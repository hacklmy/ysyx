module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input         io_from_lsu_rready,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [31:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  input         io_from_lsu_bready,
  output        io_to_lsu_arready,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_awready,
  output        io_to_lsu_wready,
  output        io_to_lsu_bvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output        io_to_axi_awvalid,
  output [31:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input         io_from_axi_arready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid,
  input         io_from_axi_awready,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [63:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [63:0] _RAND_260;
  reg [31:0] _RAND_261;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = ~reset; // @[d_cache.scala 15:11]
  reg [63:0] ram_0_0; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_1; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_2; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_3; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_4; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_5; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_6; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_7; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_8; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_9; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_10; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_11; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_12; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_13; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_14; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_15; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_16; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_17; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_18; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_19; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_20; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_21; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_22; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_23; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_24; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_25; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_26; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_27; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_28; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_29; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_30; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_31; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_32; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_33; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_34; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_35; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_36; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_37; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_38; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_39; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_40; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_41; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_42; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_43; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_44; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_45; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_46; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_47; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_48; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_49; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_50; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_51; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_52; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_53; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_54; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_55; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_56; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_57; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_58; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_59; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_60; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_61; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_62; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_63; // @[d_cache.scala 18:24]
  reg [31:0] tag_0_0; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_16; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_17; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_18; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_19; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_20; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_21; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_22; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_23; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_24; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_25; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_26; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_27; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_28; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_29; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_30; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_31; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_32; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_33; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_34; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_35; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_36; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_37; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_38; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_39; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_40; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_41; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_42; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_43; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_44; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_45; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_46; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_47; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_48; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_49; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_50; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_51; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_52; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_53; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_54; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_55; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_56; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_57; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_58; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_59; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_60; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_61; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_62; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_63; // @[d_cache.scala 22:24]
  reg  valid_0_0; // @[d_cache.scala 24:26]
  reg  valid_0_1; // @[d_cache.scala 24:26]
  reg  valid_0_2; // @[d_cache.scala 24:26]
  reg  valid_0_3; // @[d_cache.scala 24:26]
  reg  valid_0_4; // @[d_cache.scala 24:26]
  reg  valid_0_5; // @[d_cache.scala 24:26]
  reg  valid_0_6; // @[d_cache.scala 24:26]
  reg  valid_0_7; // @[d_cache.scala 24:26]
  reg  valid_0_8; // @[d_cache.scala 24:26]
  reg  valid_0_9; // @[d_cache.scala 24:26]
  reg  valid_0_10; // @[d_cache.scala 24:26]
  reg  valid_0_11; // @[d_cache.scala 24:26]
  reg  valid_0_12; // @[d_cache.scala 24:26]
  reg  valid_0_13; // @[d_cache.scala 24:26]
  reg  valid_0_14; // @[d_cache.scala 24:26]
  reg  valid_0_15; // @[d_cache.scala 24:26]
  reg  valid_0_16; // @[d_cache.scala 24:26]
  reg  valid_0_17; // @[d_cache.scala 24:26]
  reg  valid_0_18; // @[d_cache.scala 24:26]
  reg  valid_0_19; // @[d_cache.scala 24:26]
  reg  valid_0_20; // @[d_cache.scala 24:26]
  reg  valid_0_21; // @[d_cache.scala 24:26]
  reg  valid_0_22; // @[d_cache.scala 24:26]
  reg  valid_0_23; // @[d_cache.scala 24:26]
  reg  valid_0_24; // @[d_cache.scala 24:26]
  reg  valid_0_25; // @[d_cache.scala 24:26]
  reg  valid_0_26; // @[d_cache.scala 24:26]
  reg  valid_0_27; // @[d_cache.scala 24:26]
  reg  valid_0_28; // @[d_cache.scala 24:26]
  reg  valid_0_29; // @[d_cache.scala 24:26]
  reg  valid_0_30; // @[d_cache.scala 24:26]
  reg  valid_0_31; // @[d_cache.scala 24:26]
  reg  valid_0_32; // @[d_cache.scala 24:26]
  reg  valid_0_33; // @[d_cache.scala 24:26]
  reg  valid_0_34; // @[d_cache.scala 24:26]
  reg  valid_0_35; // @[d_cache.scala 24:26]
  reg  valid_0_36; // @[d_cache.scala 24:26]
  reg  valid_0_37; // @[d_cache.scala 24:26]
  reg  valid_0_38; // @[d_cache.scala 24:26]
  reg  valid_0_39; // @[d_cache.scala 24:26]
  reg  valid_0_40; // @[d_cache.scala 24:26]
  reg  valid_0_41; // @[d_cache.scala 24:26]
  reg  valid_0_42; // @[d_cache.scala 24:26]
  reg  valid_0_43; // @[d_cache.scala 24:26]
  reg  valid_0_44; // @[d_cache.scala 24:26]
  reg  valid_0_45; // @[d_cache.scala 24:26]
  reg  valid_0_46; // @[d_cache.scala 24:26]
  reg  valid_0_47; // @[d_cache.scala 24:26]
  reg  valid_0_48; // @[d_cache.scala 24:26]
  reg  valid_0_49; // @[d_cache.scala 24:26]
  reg  valid_0_50; // @[d_cache.scala 24:26]
  reg  valid_0_51; // @[d_cache.scala 24:26]
  reg  valid_0_52; // @[d_cache.scala 24:26]
  reg  valid_0_53; // @[d_cache.scala 24:26]
  reg  valid_0_54; // @[d_cache.scala 24:26]
  reg  valid_0_55; // @[d_cache.scala 24:26]
  reg  valid_0_56; // @[d_cache.scala 24:26]
  reg  valid_0_57; // @[d_cache.scala 24:26]
  reg  valid_0_58; // @[d_cache.scala 24:26]
  reg  valid_0_59; // @[d_cache.scala 24:26]
  reg  valid_0_60; // @[d_cache.scala 24:26]
  reg  valid_0_61; // @[d_cache.scala 24:26]
  reg  valid_0_62; // @[d_cache.scala 24:26]
  reg  valid_0_63; // @[d_cache.scala 24:26]
  reg  dirty_0_0; // @[d_cache.scala 26:26]
  reg  dirty_0_1; // @[d_cache.scala 26:26]
  reg  dirty_0_2; // @[d_cache.scala 26:26]
  reg  dirty_0_3; // @[d_cache.scala 26:26]
  reg  dirty_0_4; // @[d_cache.scala 26:26]
  reg  dirty_0_5; // @[d_cache.scala 26:26]
  reg  dirty_0_6; // @[d_cache.scala 26:26]
  reg  dirty_0_7; // @[d_cache.scala 26:26]
  reg  dirty_0_8; // @[d_cache.scala 26:26]
  reg  dirty_0_9; // @[d_cache.scala 26:26]
  reg  dirty_0_10; // @[d_cache.scala 26:26]
  reg  dirty_0_11; // @[d_cache.scala 26:26]
  reg  dirty_0_12; // @[d_cache.scala 26:26]
  reg  dirty_0_13; // @[d_cache.scala 26:26]
  reg  dirty_0_14; // @[d_cache.scala 26:26]
  reg  dirty_0_15; // @[d_cache.scala 26:26]
  reg  dirty_0_16; // @[d_cache.scala 26:26]
  reg  dirty_0_17; // @[d_cache.scala 26:26]
  reg  dirty_0_18; // @[d_cache.scala 26:26]
  reg  dirty_0_19; // @[d_cache.scala 26:26]
  reg  dirty_0_20; // @[d_cache.scala 26:26]
  reg  dirty_0_21; // @[d_cache.scala 26:26]
  reg  dirty_0_22; // @[d_cache.scala 26:26]
  reg  dirty_0_23; // @[d_cache.scala 26:26]
  reg  dirty_0_24; // @[d_cache.scala 26:26]
  reg  dirty_0_25; // @[d_cache.scala 26:26]
  reg  dirty_0_26; // @[d_cache.scala 26:26]
  reg  dirty_0_27; // @[d_cache.scala 26:26]
  reg  dirty_0_28; // @[d_cache.scala 26:26]
  reg  dirty_0_29; // @[d_cache.scala 26:26]
  reg  dirty_0_30; // @[d_cache.scala 26:26]
  reg  dirty_0_31; // @[d_cache.scala 26:26]
  reg  dirty_0_32; // @[d_cache.scala 26:26]
  reg  dirty_0_33; // @[d_cache.scala 26:26]
  reg  dirty_0_34; // @[d_cache.scala 26:26]
  reg  dirty_0_35; // @[d_cache.scala 26:26]
  reg  dirty_0_36; // @[d_cache.scala 26:26]
  reg  dirty_0_37; // @[d_cache.scala 26:26]
  reg  dirty_0_38; // @[d_cache.scala 26:26]
  reg  dirty_0_39; // @[d_cache.scala 26:26]
  reg  dirty_0_40; // @[d_cache.scala 26:26]
  reg  dirty_0_41; // @[d_cache.scala 26:26]
  reg  dirty_0_42; // @[d_cache.scala 26:26]
  reg  dirty_0_43; // @[d_cache.scala 26:26]
  reg  dirty_0_44; // @[d_cache.scala 26:26]
  reg  dirty_0_45; // @[d_cache.scala 26:26]
  reg  dirty_0_46; // @[d_cache.scala 26:26]
  reg  dirty_0_47; // @[d_cache.scala 26:26]
  reg  dirty_0_48; // @[d_cache.scala 26:26]
  reg  dirty_0_49; // @[d_cache.scala 26:26]
  reg  dirty_0_50; // @[d_cache.scala 26:26]
  reg  dirty_0_51; // @[d_cache.scala 26:26]
  reg  dirty_0_52; // @[d_cache.scala 26:26]
  reg  dirty_0_53; // @[d_cache.scala 26:26]
  reg  dirty_0_54; // @[d_cache.scala 26:26]
  reg  dirty_0_55; // @[d_cache.scala 26:26]
  reg  dirty_0_56; // @[d_cache.scala 26:26]
  reg  dirty_0_57; // @[d_cache.scala 26:26]
  reg  dirty_0_58; // @[d_cache.scala 26:26]
  reg  dirty_0_59; // @[d_cache.scala 26:26]
  reg  dirty_0_60; // @[d_cache.scala 26:26]
  reg  dirty_0_61; // @[d_cache.scala 26:26]
  reg  dirty_0_62; // @[d_cache.scala 26:26]
  reg  dirty_0_63; // @[d_cache.scala 26:26]
  reg  way0_hit; // @[d_cache.scala 28:27]
  reg [63:0] write_back_data; // @[d_cache.scala 31:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 32:34]
  reg [1:0] unuse_way; // @[d_cache.scala 35:28]
  reg [63:0] receive_data; // @[d_cache.scala 36:31]
  wire [2:0] offset = io_from_lsu_araddr[2:0]; // @[d_cache.scala 39:36]
  wire [5:0] index = io_from_lsu_araddr[8:3]; // @[d_cache.scala 40:35]
  wire [22:0] tag = io_from_lsu_araddr[31:9]; // @[d_cache.scala 41:33]
  wire [5:0] _shift_bit_T_8 = offset == 3'h7 ? 6'h38 : 6'h0; // @[d_cache.scala 50:24]
  wire [5:0] _shift_bit_T_9 = offset == 3'h6 ? 6'h30 : _shift_bit_T_8; // @[d_cache.scala 49:24]
  wire [5:0] _shift_bit_T_10 = offset == 3'h5 ? 6'h28 : _shift_bit_T_9; // @[d_cache.scala 48:24]
  wire [5:0] _shift_bit_T_11 = offset == 3'h4 ? 6'h20 : _shift_bit_T_10; // @[d_cache.scala 47:24]
  wire [5:0] _shift_bit_T_12 = offset == 3'h3 ? 6'h18 : _shift_bit_T_11; // @[d_cache.scala 46:24]
  wire [5:0] _shift_bit_T_13 = offset == 3'h2 ? 6'h10 : _shift_bit_T_12; // @[d_cache.scala 45:24]
  wire [5:0] _shift_bit_T_14 = offset == 3'h1 ? 6'h8 : _shift_bit_T_13; // @[d_cache.scala 44:24]
  wire [5:0] shift_bit = offset == 3'h0 ? 6'h0 : _shift_bit_T_14; // @[d_cache.scala 43:24]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 55:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 54:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 53:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 52:20]
  wire [31:0] _GEN_1 = 6'h1 == index ? tag_0_1 : tag_0_0; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_2 = 6'h2 == index ? tag_0_2 : _GEN_1; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_3 = 6'h3 == index ? tag_0_3 : _GEN_2; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_4 = 6'h4 == index ? tag_0_4 : _GEN_3; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_5 = 6'h5 == index ? tag_0_5 : _GEN_4; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_6 = 6'h6 == index ? tag_0_6 : _GEN_5; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_7 = 6'h7 == index ? tag_0_7 : _GEN_6; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_8 = 6'h8 == index ? tag_0_8 : _GEN_7; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_9 = 6'h9 == index ? tag_0_9 : _GEN_8; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_10 = 6'ha == index ? tag_0_10 : _GEN_9; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_11 = 6'hb == index ? tag_0_11 : _GEN_10; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_12 = 6'hc == index ? tag_0_12 : _GEN_11; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_13 = 6'hd == index ? tag_0_13 : _GEN_12; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_14 = 6'he == index ? tag_0_14 : _GEN_13; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_15 = 6'hf == index ? tag_0_15 : _GEN_14; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_16 = 6'h10 == index ? tag_0_16 : _GEN_15; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_17 = 6'h11 == index ? tag_0_17 : _GEN_16; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_18 = 6'h12 == index ? tag_0_18 : _GEN_17; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_19 = 6'h13 == index ? tag_0_19 : _GEN_18; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_20 = 6'h14 == index ? tag_0_20 : _GEN_19; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_21 = 6'h15 == index ? tag_0_21 : _GEN_20; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_22 = 6'h16 == index ? tag_0_22 : _GEN_21; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_23 = 6'h17 == index ? tag_0_23 : _GEN_22; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_24 = 6'h18 == index ? tag_0_24 : _GEN_23; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_25 = 6'h19 == index ? tag_0_25 : _GEN_24; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_26 = 6'h1a == index ? tag_0_26 : _GEN_25; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_27 = 6'h1b == index ? tag_0_27 : _GEN_26; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_28 = 6'h1c == index ? tag_0_28 : _GEN_27; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_29 = 6'h1d == index ? tag_0_29 : _GEN_28; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_30 = 6'h1e == index ? tag_0_30 : _GEN_29; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_31 = 6'h1f == index ? tag_0_31 : _GEN_30; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_32 = 6'h20 == index ? tag_0_32 : _GEN_31; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_33 = 6'h21 == index ? tag_0_33 : _GEN_32; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_34 = 6'h22 == index ? tag_0_34 : _GEN_33; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_35 = 6'h23 == index ? tag_0_35 : _GEN_34; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_36 = 6'h24 == index ? tag_0_36 : _GEN_35; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_37 = 6'h25 == index ? tag_0_37 : _GEN_36; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_38 = 6'h26 == index ? tag_0_38 : _GEN_37; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_39 = 6'h27 == index ? tag_0_39 : _GEN_38; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_40 = 6'h28 == index ? tag_0_40 : _GEN_39; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_41 = 6'h29 == index ? tag_0_41 : _GEN_40; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_42 = 6'h2a == index ? tag_0_42 : _GEN_41; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_43 = 6'h2b == index ? tag_0_43 : _GEN_42; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_44 = 6'h2c == index ? tag_0_44 : _GEN_43; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_45 = 6'h2d == index ? tag_0_45 : _GEN_44; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_46 = 6'h2e == index ? tag_0_46 : _GEN_45; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_47 = 6'h2f == index ? tag_0_47 : _GEN_46; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_48 = 6'h30 == index ? tag_0_48 : _GEN_47; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_49 = 6'h31 == index ? tag_0_49 : _GEN_48; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_50 = 6'h32 == index ? tag_0_50 : _GEN_49; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_51 = 6'h33 == index ? tag_0_51 : _GEN_50; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_52 = 6'h34 == index ? tag_0_52 : _GEN_51; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_53 = 6'h35 == index ? tag_0_53 : _GEN_52; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_54 = 6'h36 == index ? tag_0_54 : _GEN_53; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_55 = 6'h37 == index ? tag_0_55 : _GEN_54; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_56 = 6'h38 == index ? tag_0_56 : _GEN_55; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_57 = 6'h39 == index ? tag_0_57 : _GEN_56; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_58 = 6'h3a == index ? tag_0_58 : _GEN_57; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_59 = 6'h3b == index ? tag_0_59 : _GEN_58; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_60 = 6'h3c == index ? tag_0_60 : _GEN_59; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_61 = 6'h3d == index ? tag_0_61 : _GEN_60; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_62 = 6'h3e == index ? tag_0_62 : _GEN_61; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_63 = 6'h3f == index ? tag_0_63 : _GEN_62; // @[d_cache.scala 57:{24,24}]
  wire [31:0] _GEN_3460 = {{9'd0}, tag}; // @[d_cache.scala 57:24]
  wire  _GEN_65 = 6'h1 == index ? valid_0_1 : valid_0_0; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_66 = 6'h2 == index ? valid_0_2 : _GEN_65; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_67 = 6'h3 == index ? valid_0_3 : _GEN_66; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_68 = 6'h4 == index ? valid_0_4 : _GEN_67; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_69 = 6'h5 == index ? valid_0_5 : _GEN_68; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_70 = 6'h6 == index ? valid_0_6 : _GEN_69; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_71 = 6'h7 == index ? valid_0_7 : _GEN_70; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_72 = 6'h8 == index ? valid_0_8 : _GEN_71; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_73 = 6'h9 == index ? valid_0_9 : _GEN_72; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_74 = 6'ha == index ? valid_0_10 : _GEN_73; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_75 = 6'hb == index ? valid_0_11 : _GEN_74; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_76 = 6'hc == index ? valid_0_12 : _GEN_75; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_77 = 6'hd == index ? valid_0_13 : _GEN_76; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_78 = 6'he == index ? valid_0_14 : _GEN_77; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_79 = 6'hf == index ? valid_0_15 : _GEN_78; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_80 = 6'h10 == index ? valid_0_16 : _GEN_79; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_81 = 6'h11 == index ? valid_0_17 : _GEN_80; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_82 = 6'h12 == index ? valid_0_18 : _GEN_81; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_83 = 6'h13 == index ? valid_0_19 : _GEN_82; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_84 = 6'h14 == index ? valid_0_20 : _GEN_83; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_85 = 6'h15 == index ? valid_0_21 : _GEN_84; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_86 = 6'h16 == index ? valid_0_22 : _GEN_85; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_87 = 6'h17 == index ? valid_0_23 : _GEN_86; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_88 = 6'h18 == index ? valid_0_24 : _GEN_87; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_89 = 6'h19 == index ? valid_0_25 : _GEN_88; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_90 = 6'h1a == index ? valid_0_26 : _GEN_89; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_91 = 6'h1b == index ? valid_0_27 : _GEN_90; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_92 = 6'h1c == index ? valid_0_28 : _GEN_91; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_93 = 6'h1d == index ? valid_0_29 : _GEN_92; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_94 = 6'h1e == index ? valid_0_30 : _GEN_93; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_95 = 6'h1f == index ? valid_0_31 : _GEN_94; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_96 = 6'h20 == index ? valid_0_32 : _GEN_95; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_97 = 6'h21 == index ? valid_0_33 : _GEN_96; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_98 = 6'h22 == index ? valid_0_34 : _GEN_97; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_99 = 6'h23 == index ? valid_0_35 : _GEN_98; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_100 = 6'h24 == index ? valid_0_36 : _GEN_99; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_101 = 6'h25 == index ? valid_0_37 : _GEN_100; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_102 = 6'h26 == index ? valid_0_38 : _GEN_101; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_103 = 6'h27 == index ? valid_0_39 : _GEN_102; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_104 = 6'h28 == index ? valid_0_40 : _GEN_103; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_105 = 6'h29 == index ? valid_0_41 : _GEN_104; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_106 = 6'h2a == index ? valid_0_42 : _GEN_105; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_107 = 6'h2b == index ? valid_0_43 : _GEN_106; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_108 = 6'h2c == index ? valid_0_44 : _GEN_107; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_109 = 6'h2d == index ? valid_0_45 : _GEN_108; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_110 = 6'h2e == index ? valid_0_46 : _GEN_109; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_111 = 6'h2f == index ? valid_0_47 : _GEN_110; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_112 = 6'h30 == index ? valid_0_48 : _GEN_111; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_113 = 6'h31 == index ? valid_0_49 : _GEN_112; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_114 = 6'h32 == index ? valid_0_50 : _GEN_113; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_115 = 6'h33 == index ? valid_0_51 : _GEN_114; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_116 = 6'h34 == index ? valid_0_52 : _GEN_115; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_117 = 6'h35 == index ? valid_0_53 : _GEN_116; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_118 = 6'h36 == index ? valid_0_54 : _GEN_117; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_119 = 6'h37 == index ? valid_0_55 : _GEN_118; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_120 = 6'h38 == index ? valid_0_56 : _GEN_119; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_121 = 6'h39 == index ? valid_0_57 : _GEN_120; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_122 = 6'h3a == index ? valid_0_58 : _GEN_121; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_123 = 6'h3b == index ? valid_0_59 : _GEN_122; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_124 = 6'h3c == index ? valid_0_60 : _GEN_123; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_125 = 6'h3d == index ? valid_0_61 : _GEN_124; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_126 = 6'h3e == index ? valid_0_62 : _GEN_125; // @[d_cache.scala 57:{50,50}]
  wire  _GEN_127 = 6'h3f == index ? valid_0_63 : _GEN_126; // @[d_cache.scala 57:{50,50}]
  wire  _T_4 = _GEN_63 == _GEN_3460 & _GEN_127; // @[d_cache.scala 57:33]
  wire  _T_5 = ~_GEN_127; // @[d_cache.scala 68:25]
  reg [2:0] state; // @[d_cache.scala 76:24]
  wire  _T_10 = 3'h0 == state; // @[d_cache.scala 81:18]
  wire  _T_11 = 3'h1 == state; // @[d_cache.scala 81:18]
  wire  _GEN_133 = 6'h1 == index ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_134 = 6'h2 == index ? dirty_0_2 : _GEN_133; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_135 = 6'h3 == index ? dirty_0_3 : _GEN_134; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_136 = 6'h4 == index ? dirty_0_4 : _GEN_135; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_137 = 6'h5 == index ? dirty_0_5 : _GEN_136; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_138 = 6'h6 == index ? dirty_0_6 : _GEN_137; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_139 = 6'h7 == index ? dirty_0_7 : _GEN_138; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_140 = 6'h8 == index ? dirty_0_8 : _GEN_139; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_141 = 6'h9 == index ? dirty_0_9 : _GEN_140; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_142 = 6'ha == index ? dirty_0_10 : _GEN_141; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_143 = 6'hb == index ? dirty_0_11 : _GEN_142; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_144 = 6'hc == index ? dirty_0_12 : _GEN_143; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_145 = 6'hd == index ? dirty_0_13 : _GEN_144; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_146 = 6'he == index ? dirty_0_14 : _GEN_145; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_147 = 6'hf == index ? dirty_0_15 : _GEN_146; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_148 = 6'h10 == index ? dirty_0_16 : _GEN_147; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_149 = 6'h11 == index ? dirty_0_17 : _GEN_148; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_150 = 6'h12 == index ? dirty_0_18 : _GEN_149; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_151 = 6'h13 == index ? dirty_0_19 : _GEN_150; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_152 = 6'h14 == index ? dirty_0_20 : _GEN_151; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_153 = 6'h15 == index ? dirty_0_21 : _GEN_152; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_154 = 6'h16 == index ? dirty_0_22 : _GEN_153; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_155 = 6'h17 == index ? dirty_0_23 : _GEN_154; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_156 = 6'h18 == index ? dirty_0_24 : _GEN_155; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_157 = 6'h19 == index ? dirty_0_25 : _GEN_156; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_158 = 6'h1a == index ? dirty_0_26 : _GEN_157; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_159 = 6'h1b == index ? dirty_0_27 : _GEN_158; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_160 = 6'h1c == index ? dirty_0_28 : _GEN_159; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_161 = 6'h1d == index ? dirty_0_29 : _GEN_160; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_162 = 6'h1e == index ? dirty_0_30 : _GEN_161; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_163 = 6'h1f == index ? dirty_0_31 : _GEN_162; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_164 = 6'h20 == index ? dirty_0_32 : _GEN_163; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_165 = 6'h21 == index ? dirty_0_33 : _GEN_164; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_166 = 6'h22 == index ? dirty_0_34 : _GEN_165; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_167 = 6'h23 == index ? dirty_0_35 : _GEN_166; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_168 = 6'h24 == index ? dirty_0_36 : _GEN_167; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_169 = 6'h25 == index ? dirty_0_37 : _GEN_168; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_170 = 6'h26 == index ? dirty_0_38 : _GEN_169; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_171 = 6'h27 == index ? dirty_0_39 : _GEN_170; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_172 = 6'h28 == index ? dirty_0_40 : _GEN_171; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_173 = 6'h29 == index ? dirty_0_41 : _GEN_172; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_174 = 6'h2a == index ? dirty_0_42 : _GEN_173; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_175 = 6'h2b == index ? dirty_0_43 : _GEN_174; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_176 = 6'h2c == index ? dirty_0_44 : _GEN_175; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_177 = 6'h2d == index ? dirty_0_45 : _GEN_176; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_178 = 6'h2e == index ? dirty_0_46 : _GEN_177; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_179 = 6'h2f == index ? dirty_0_47 : _GEN_178; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_180 = 6'h30 == index ? dirty_0_48 : _GEN_179; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_181 = 6'h31 == index ? dirty_0_49 : _GEN_180; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_182 = 6'h32 == index ? dirty_0_50 : _GEN_181; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_183 = 6'h33 == index ? dirty_0_51 : _GEN_182; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_184 = 6'h34 == index ? dirty_0_52 : _GEN_183; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_185 = 6'h35 == index ? dirty_0_53 : _GEN_184; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_186 = 6'h36 == index ? dirty_0_54 : _GEN_185; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_187 = 6'h37 == index ? dirty_0_55 : _GEN_186; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_188 = 6'h38 == index ? dirty_0_56 : _GEN_187; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_189 = 6'h39 == index ? dirty_0_57 : _GEN_188; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_190 = 6'h3a == index ? dirty_0_58 : _GEN_189; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_191 = 6'h3b == index ? dirty_0_59 : _GEN_190; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_192 = 6'h3c == index ? dirty_0_60 : _GEN_191; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_193 = 6'h3d == index ? dirty_0_61 : _GEN_192; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_194 = 6'h3e == index ? dirty_0_62 : _GEN_193; // @[d_cache.scala 93:{27,27}]
  wire  _GEN_195 = 6'h3f == index ? dirty_0_63 : _GEN_194; // @[d_cache.scala 93:{27,27}]
  wire [2:0] _GEN_196 = io_from_lsu_rready ? 3'h0 : state; // @[d_cache.scala 76:24 92:41 94:27]
  wire [63:0] _GEN_3461 = {{32'd0}, io_from_lsu_wdata}; // @[d_cache.scala 109:53]
  wire [63:0] _ram_0_T = _GEN_3461 & wmask; // @[d_cache.scala 109:53]
  wire [126:0] _GEN_3789 = {{63'd0}, _ram_0_T}; // @[d_cache.scala 109:62]
  wire [126:0] _ram_0_T_1 = _GEN_3789 << shift_bit; // @[d_cache.scala 109:62]
  wire [126:0] _GEN_3790 = {{63'd0}, wmask}; // @[d_cache.scala 109:102]
  wire [126:0] _ram_0_T_2 = _GEN_3790 << shift_bit; // @[d_cache.scala 109:102]
  wire [126:0] _ram_0_T_3 = ~_ram_0_T_2; // @[d_cache.scala 109:94]
  wire [63:0] _GEN_199 = 6'h1 == index ? ram_0_1 : ram_0_0; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_200 = 6'h2 == index ? ram_0_2 : _GEN_199; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_201 = 6'h3 == index ? ram_0_3 : _GEN_200; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_202 = 6'h4 == index ? ram_0_4 : _GEN_201; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_203 = 6'h5 == index ? ram_0_5 : _GEN_202; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_204 = 6'h6 == index ? ram_0_6 : _GEN_203; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_205 = 6'h7 == index ? ram_0_7 : _GEN_204; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_206 = 6'h8 == index ? ram_0_8 : _GEN_205; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_207 = 6'h9 == index ? ram_0_9 : _GEN_206; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_208 = 6'ha == index ? ram_0_10 : _GEN_207; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_209 = 6'hb == index ? ram_0_11 : _GEN_208; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_210 = 6'hc == index ? ram_0_12 : _GEN_209; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_211 = 6'hd == index ? ram_0_13 : _GEN_210; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_212 = 6'he == index ? ram_0_14 : _GEN_211; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_213 = 6'hf == index ? ram_0_15 : _GEN_212; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_214 = 6'h10 == index ? ram_0_16 : _GEN_213; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_215 = 6'h11 == index ? ram_0_17 : _GEN_214; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_216 = 6'h12 == index ? ram_0_18 : _GEN_215; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_217 = 6'h13 == index ? ram_0_19 : _GEN_216; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_218 = 6'h14 == index ? ram_0_20 : _GEN_217; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_219 = 6'h15 == index ? ram_0_21 : _GEN_218; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_220 = 6'h16 == index ? ram_0_22 : _GEN_219; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_221 = 6'h17 == index ? ram_0_23 : _GEN_220; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_222 = 6'h18 == index ? ram_0_24 : _GEN_221; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_223 = 6'h19 == index ? ram_0_25 : _GEN_222; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_224 = 6'h1a == index ? ram_0_26 : _GEN_223; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_225 = 6'h1b == index ? ram_0_27 : _GEN_224; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_226 = 6'h1c == index ? ram_0_28 : _GEN_225; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_227 = 6'h1d == index ? ram_0_29 : _GEN_226; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_228 = 6'h1e == index ? ram_0_30 : _GEN_227; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_229 = 6'h1f == index ? ram_0_31 : _GEN_228; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_230 = 6'h20 == index ? ram_0_32 : _GEN_229; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_231 = 6'h21 == index ? ram_0_33 : _GEN_230; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_232 = 6'h22 == index ? ram_0_34 : _GEN_231; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_233 = 6'h23 == index ? ram_0_35 : _GEN_232; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_234 = 6'h24 == index ? ram_0_36 : _GEN_233; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_235 = 6'h25 == index ? ram_0_37 : _GEN_234; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_236 = 6'h26 == index ? ram_0_38 : _GEN_235; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_237 = 6'h27 == index ? ram_0_39 : _GEN_236; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_238 = 6'h28 == index ? ram_0_40 : _GEN_237; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_239 = 6'h29 == index ? ram_0_41 : _GEN_238; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_240 = 6'h2a == index ? ram_0_42 : _GEN_239; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_241 = 6'h2b == index ? ram_0_43 : _GEN_240; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_242 = 6'h2c == index ? ram_0_44 : _GEN_241; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_243 = 6'h2d == index ? ram_0_45 : _GEN_242; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_244 = 6'h2e == index ? ram_0_46 : _GEN_243; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_245 = 6'h2f == index ? ram_0_47 : _GEN_244; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_246 = 6'h30 == index ? ram_0_48 : _GEN_245; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_247 = 6'h31 == index ? ram_0_49 : _GEN_246; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_248 = 6'h32 == index ? ram_0_50 : _GEN_247; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_249 = 6'h33 == index ? ram_0_51 : _GEN_248; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_250 = 6'h34 == index ? ram_0_52 : _GEN_249; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_251 = 6'h35 == index ? ram_0_53 : _GEN_250; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_252 = 6'h36 == index ? ram_0_54 : _GEN_251; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_253 = 6'h37 == index ? ram_0_55 : _GEN_252; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_254 = 6'h38 == index ? ram_0_56 : _GEN_253; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_255 = 6'h39 == index ? ram_0_57 : _GEN_254; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_256 = 6'h3a == index ? ram_0_58 : _GEN_255; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_257 = 6'h3b == index ? ram_0_59 : _GEN_256; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_258 = 6'h3c == index ? ram_0_60 : _GEN_257; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_259 = 6'h3d == index ? ram_0_61 : _GEN_258; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_260 = 6'h3e == index ? ram_0_62 : _GEN_259; // @[d_cache.scala 109:{92,92}]
  wire [63:0] _GEN_261 = 6'h3f == index ? ram_0_63 : _GEN_260; // @[d_cache.scala 109:{92,92}]
  wire [126:0] _GEN_3462 = {{63'd0}, _GEN_261}; // @[d_cache.scala 109:92]
  wire [126:0] _ram_0_T_4 = _GEN_3462 & _ram_0_T_3; // @[d_cache.scala 109:92]
  wire [126:0] _ram_0_T_5 = _ram_0_T_1 | _ram_0_T_4; // @[d_cache.scala 109:76]
  wire [63:0] _GEN_262 = 6'h0 == index ? _ram_0_T_5[63:0] : ram_0_0; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_263 = 6'h1 == index ? _ram_0_T_5[63:0] : ram_0_1; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_264 = 6'h2 == index ? _ram_0_T_5[63:0] : ram_0_2; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_265 = 6'h3 == index ? _ram_0_T_5[63:0] : ram_0_3; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_266 = 6'h4 == index ? _ram_0_T_5[63:0] : ram_0_4; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_267 = 6'h5 == index ? _ram_0_T_5[63:0] : ram_0_5; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_268 = 6'h6 == index ? _ram_0_T_5[63:0] : ram_0_6; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_269 = 6'h7 == index ? _ram_0_T_5[63:0] : ram_0_7; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_270 = 6'h8 == index ? _ram_0_T_5[63:0] : ram_0_8; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_271 = 6'h9 == index ? _ram_0_T_5[63:0] : ram_0_9; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_272 = 6'ha == index ? _ram_0_T_5[63:0] : ram_0_10; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_273 = 6'hb == index ? _ram_0_T_5[63:0] : ram_0_11; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_274 = 6'hc == index ? _ram_0_T_5[63:0] : ram_0_12; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_275 = 6'hd == index ? _ram_0_T_5[63:0] : ram_0_13; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_276 = 6'he == index ? _ram_0_T_5[63:0] : ram_0_14; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_277 = 6'hf == index ? _ram_0_T_5[63:0] : ram_0_15; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_278 = 6'h10 == index ? _ram_0_T_5[63:0] : ram_0_16; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_279 = 6'h11 == index ? _ram_0_T_5[63:0] : ram_0_17; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_280 = 6'h12 == index ? _ram_0_T_5[63:0] : ram_0_18; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_281 = 6'h13 == index ? _ram_0_T_5[63:0] : ram_0_19; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_282 = 6'h14 == index ? _ram_0_T_5[63:0] : ram_0_20; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_283 = 6'h15 == index ? _ram_0_T_5[63:0] : ram_0_21; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_284 = 6'h16 == index ? _ram_0_T_5[63:0] : ram_0_22; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_285 = 6'h17 == index ? _ram_0_T_5[63:0] : ram_0_23; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_286 = 6'h18 == index ? _ram_0_T_5[63:0] : ram_0_24; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_287 = 6'h19 == index ? _ram_0_T_5[63:0] : ram_0_25; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_288 = 6'h1a == index ? _ram_0_T_5[63:0] : ram_0_26; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_289 = 6'h1b == index ? _ram_0_T_5[63:0] : ram_0_27; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_290 = 6'h1c == index ? _ram_0_T_5[63:0] : ram_0_28; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_291 = 6'h1d == index ? _ram_0_T_5[63:0] : ram_0_29; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_292 = 6'h1e == index ? _ram_0_T_5[63:0] : ram_0_30; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_293 = 6'h1f == index ? _ram_0_T_5[63:0] : ram_0_31; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_294 = 6'h20 == index ? _ram_0_T_5[63:0] : ram_0_32; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_295 = 6'h21 == index ? _ram_0_T_5[63:0] : ram_0_33; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_296 = 6'h22 == index ? _ram_0_T_5[63:0] : ram_0_34; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_297 = 6'h23 == index ? _ram_0_T_5[63:0] : ram_0_35; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_298 = 6'h24 == index ? _ram_0_T_5[63:0] : ram_0_36; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_299 = 6'h25 == index ? _ram_0_T_5[63:0] : ram_0_37; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_300 = 6'h26 == index ? _ram_0_T_5[63:0] : ram_0_38; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_301 = 6'h27 == index ? _ram_0_T_5[63:0] : ram_0_39; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_302 = 6'h28 == index ? _ram_0_T_5[63:0] : ram_0_40; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_303 = 6'h29 == index ? _ram_0_T_5[63:0] : ram_0_41; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_304 = 6'h2a == index ? _ram_0_T_5[63:0] : ram_0_42; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_305 = 6'h2b == index ? _ram_0_T_5[63:0] : ram_0_43; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_306 = 6'h2c == index ? _ram_0_T_5[63:0] : ram_0_44; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_307 = 6'h2d == index ? _ram_0_T_5[63:0] : ram_0_45; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_308 = 6'h2e == index ? _ram_0_T_5[63:0] : ram_0_46; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_309 = 6'h2f == index ? _ram_0_T_5[63:0] : ram_0_47; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_310 = 6'h30 == index ? _ram_0_T_5[63:0] : ram_0_48; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_311 = 6'h31 == index ? _ram_0_T_5[63:0] : ram_0_49; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_312 = 6'h32 == index ? _ram_0_T_5[63:0] : ram_0_50; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_313 = 6'h33 == index ? _ram_0_T_5[63:0] : ram_0_51; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_314 = 6'h34 == index ? _ram_0_T_5[63:0] : ram_0_52; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_315 = 6'h35 == index ? _ram_0_T_5[63:0] : ram_0_53; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_316 = 6'h36 == index ? _ram_0_T_5[63:0] : ram_0_54; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_317 = 6'h37 == index ? _ram_0_T_5[63:0] : ram_0_55; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_318 = 6'h38 == index ? _ram_0_T_5[63:0] : ram_0_56; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_319 = 6'h39 == index ? _ram_0_T_5[63:0] : ram_0_57; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_320 = 6'h3a == index ? _ram_0_T_5[63:0] : ram_0_58; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_321 = 6'h3b == index ? _ram_0_T_5[63:0] : ram_0_59; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_322 = 6'h3c == index ? _ram_0_T_5[63:0] : ram_0_60; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_323 = 6'h3d == index ? _ram_0_T_5[63:0] : ram_0_61; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_324 = 6'h3e == index ? _ram_0_T_5[63:0] : ram_0_62; // @[d_cache.scala 109:{30,30} 18:24]
  wire [63:0] _GEN_325 = 6'h3f == index ? _ram_0_T_5[63:0] : ram_0_63; // @[d_cache.scala 109:{30,30} 18:24]
  wire  _GEN_3463 = 6'h0 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_326 = 6'h0 == index | valid_0_0; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3464 = 6'h1 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_327 = 6'h1 == index | valid_0_1; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3465 = 6'h2 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_328 = 6'h2 == index | valid_0_2; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3466 = 6'h3 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_329 = 6'h3 == index | valid_0_3; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3467 = 6'h4 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_330 = 6'h4 == index | valid_0_4; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3468 = 6'h5 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_331 = 6'h5 == index | valid_0_5; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3469 = 6'h6 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_332 = 6'h6 == index | valid_0_6; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3470 = 6'h7 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_333 = 6'h7 == index | valid_0_7; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3471 = 6'h8 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_334 = 6'h8 == index | valid_0_8; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3472 = 6'h9 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_335 = 6'h9 == index | valid_0_9; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3473 = 6'ha == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_336 = 6'ha == index | valid_0_10; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3474 = 6'hb == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_337 = 6'hb == index | valid_0_11; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3475 = 6'hc == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_338 = 6'hc == index | valid_0_12; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3476 = 6'hd == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_339 = 6'hd == index | valid_0_13; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3477 = 6'he == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_340 = 6'he == index | valid_0_14; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3478 = 6'hf == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_341 = 6'hf == index | valid_0_15; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3479 = 6'h10 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_342 = 6'h10 == index | valid_0_16; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3480 = 6'h11 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_343 = 6'h11 == index | valid_0_17; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3481 = 6'h12 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_344 = 6'h12 == index | valid_0_18; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3482 = 6'h13 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_345 = 6'h13 == index | valid_0_19; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3483 = 6'h14 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_346 = 6'h14 == index | valid_0_20; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3484 = 6'h15 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_347 = 6'h15 == index | valid_0_21; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3485 = 6'h16 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_348 = 6'h16 == index | valid_0_22; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3486 = 6'h17 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_349 = 6'h17 == index | valid_0_23; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3487 = 6'h18 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_350 = 6'h18 == index | valid_0_24; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3488 = 6'h19 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_351 = 6'h19 == index | valid_0_25; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3489 = 6'h1a == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_352 = 6'h1a == index | valid_0_26; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3490 = 6'h1b == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_353 = 6'h1b == index | valid_0_27; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3491 = 6'h1c == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_354 = 6'h1c == index | valid_0_28; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3492 = 6'h1d == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_355 = 6'h1d == index | valid_0_29; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3493 = 6'h1e == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_356 = 6'h1e == index | valid_0_30; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3494 = 6'h1f == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_357 = 6'h1f == index | valid_0_31; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3495 = 6'h20 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_358 = 6'h20 == index | valid_0_32; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3496 = 6'h21 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_359 = 6'h21 == index | valid_0_33; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3497 = 6'h22 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_360 = 6'h22 == index | valid_0_34; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3498 = 6'h23 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_361 = 6'h23 == index | valid_0_35; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3499 = 6'h24 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_362 = 6'h24 == index | valid_0_36; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3500 = 6'h25 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_363 = 6'h25 == index | valid_0_37; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3501 = 6'h26 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_364 = 6'h26 == index | valid_0_38; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3502 = 6'h27 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_365 = 6'h27 == index | valid_0_39; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3503 = 6'h28 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_366 = 6'h28 == index | valid_0_40; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3504 = 6'h29 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_367 = 6'h29 == index | valid_0_41; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3505 = 6'h2a == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_368 = 6'h2a == index | valid_0_42; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3506 = 6'h2b == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_369 = 6'h2b == index | valid_0_43; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3507 = 6'h2c == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_370 = 6'h2c == index | valid_0_44; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3508 = 6'h2d == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_371 = 6'h2d == index | valid_0_45; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3509 = 6'h2e == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_372 = 6'h2e == index | valid_0_46; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3510 = 6'h2f == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_373 = 6'h2f == index | valid_0_47; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3511 = 6'h30 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_374 = 6'h30 == index | valid_0_48; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3512 = 6'h31 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_375 = 6'h31 == index | valid_0_49; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3513 = 6'h32 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_376 = 6'h32 == index | valid_0_50; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3514 = 6'h33 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_377 = 6'h33 == index | valid_0_51; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3515 = 6'h34 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_378 = 6'h34 == index | valid_0_52; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3516 = 6'h35 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_379 = 6'h35 == index | valid_0_53; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3517 = 6'h36 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_380 = 6'h36 == index | valid_0_54; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3518 = 6'h37 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_381 = 6'h37 == index | valid_0_55; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3519 = 6'h38 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_382 = 6'h38 == index | valid_0_56; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3520 = 6'h39 == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_383 = 6'h39 == index | valid_0_57; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3521 = 6'h3a == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_384 = 6'h3a == index | valid_0_58; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3522 = 6'h3b == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_385 = 6'h3b == index | valid_0_59; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3523 = 6'h3c == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_386 = 6'h3c == index | valid_0_60; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3524 = 6'h3d == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_387 = 6'h3d == index | valid_0_61; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3525 = 6'h3e == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_388 = 6'h3e == index | valid_0_62; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_3526 = 6'h3f == index; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_389 = 6'h3f == index | valid_0_63; // @[d_cache.scala 112:{32,32} 24:26]
  wire  _GEN_390 = _GEN_3463 | dirty_0_0; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_391 = _GEN_3464 | dirty_0_1; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_392 = _GEN_3465 | dirty_0_2; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_393 = _GEN_3466 | dirty_0_3; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_394 = _GEN_3467 | dirty_0_4; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_395 = _GEN_3468 | dirty_0_5; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_396 = _GEN_3469 | dirty_0_6; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_397 = _GEN_3470 | dirty_0_7; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_398 = _GEN_3471 | dirty_0_8; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_399 = _GEN_3472 | dirty_0_9; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_400 = _GEN_3473 | dirty_0_10; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_401 = _GEN_3474 | dirty_0_11; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_402 = _GEN_3475 | dirty_0_12; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_403 = _GEN_3476 | dirty_0_13; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_404 = _GEN_3477 | dirty_0_14; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_405 = _GEN_3478 | dirty_0_15; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_406 = _GEN_3479 | dirty_0_16; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_407 = _GEN_3480 | dirty_0_17; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_408 = _GEN_3481 | dirty_0_18; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_409 = _GEN_3482 | dirty_0_19; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_410 = _GEN_3483 | dirty_0_20; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_411 = _GEN_3484 | dirty_0_21; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_412 = _GEN_3485 | dirty_0_22; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_413 = _GEN_3486 | dirty_0_23; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_414 = _GEN_3487 | dirty_0_24; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_415 = _GEN_3488 | dirty_0_25; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_416 = _GEN_3489 | dirty_0_26; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_417 = _GEN_3490 | dirty_0_27; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_418 = _GEN_3491 | dirty_0_28; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_419 = _GEN_3492 | dirty_0_29; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_420 = _GEN_3493 | dirty_0_30; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_421 = _GEN_3494 | dirty_0_31; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_422 = _GEN_3495 | dirty_0_32; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_423 = _GEN_3496 | dirty_0_33; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_424 = _GEN_3497 | dirty_0_34; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_425 = _GEN_3498 | dirty_0_35; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_426 = _GEN_3499 | dirty_0_36; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_427 = _GEN_3500 | dirty_0_37; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_428 = _GEN_3501 | dirty_0_38; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_429 = _GEN_3502 | dirty_0_39; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_430 = _GEN_3503 | dirty_0_40; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_431 = _GEN_3504 | dirty_0_41; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_432 = _GEN_3505 | dirty_0_42; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_433 = _GEN_3506 | dirty_0_43; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_434 = _GEN_3507 | dirty_0_44; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_435 = _GEN_3508 | dirty_0_45; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_436 = _GEN_3509 | dirty_0_46; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_437 = _GEN_3510 | dirty_0_47; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_438 = _GEN_3511 | dirty_0_48; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_439 = _GEN_3512 | dirty_0_49; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_440 = _GEN_3513 | dirty_0_50; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_441 = _GEN_3514 | dirty_0_51; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_442 = _GEN_3515 | dirty_0_52; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_443 = _GEN_3516 | dirty_0_53; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_444 = _GEN_3517 | dirty_0_54; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_445 = _GEN_3518 | dirty_0_55; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_446 = _GEN_3519 | dirty_0_56; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_447 = _GEN_3520 | dirty_0_57; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_448 = _GEN_3521 | dirty_0_58; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_449 = _GEN_3522 | dirty_0_59; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_450 = _GEN_3523 | dirty_0_60; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_451 = _GEN_3524 | dirty_0_61; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_452 = _GEN_3525 | dirty_0_62; // @[d_cache.scala 113:{32,32} 26:26]
  wire  _GEN_453 = _GEN_3526 | dirty_0_63; // @[d_cache.scala 113:{32,32} 26:26]
  wire [2:0] _GEN_454 = way0_hit ? 3'h0 : 3'h4; // @[d_cache.scala 107:27 108:23 124:23]
  wire [63:0] _GEN_455 = way0_hit ? _GEN_262 : ram_0_0; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_456 = way0_hit ? _GEN_263 : ram_0_1; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_457 = way0_hit ? _GEN_264 : ram_0_2; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_458 = way0_hit ? _GEN_265 : ram_0_3; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_459 = way0_hit ? _GEN_266 : ram_0_4; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_460 = way0_hit ? _GEN_267 : ram_0_5; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_461 = way0_hit ? _GEN_268 : ram_0_6; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_462 = way0_hit ? _GEN_269 : ram_0_7; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_463 = way0_hit ? _GEN_270 : ram_0_8; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_464 = way0_hit ? _GEN_271 : ram_0_9; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_465 = way0_hit ? _GEN_272 : ram_0_10; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_466 = way0_hit ? _GEN_273 : ram_0_11; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_467 = way0_hit ? _GEN_274 : ram_0_12; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_468 = way0_hit ? _GEN_275 : ram_0_13; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_469 = way0_hit ? _GEN_276 : ram_0_14; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_470 = way0_hit ? _GEN_277 : ram_0_15; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_471 = way0_hit ? _GEN_278 : ram_0_16; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_472 = way0_hit ? _GEN_279 : ram_0_17; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_473 = way0_hit ? _GEN_280 : ram_0_18; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_474 = way0_hit ? _GEN_281 : ram_0_19; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_475 = way0_hit ? _GEN_282 : ram_0_20; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_476 = way0_hit ? _GEN_283 : ram_0_21; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_477 = way0_hit ? _GEN_284 : ram_0_22; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_478 = way0_hit ? _GEN_285 : ram_0_23; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_479 = way0_hit ? _GEN_286 : ram_0_24; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_480 = way0_hit ? _GEN_287 : ram_0_25; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_481 = way0_hit ? _GEN_288 : ram_0_26; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_482 = way0_hit ? _GEN_289 : ram_0_27; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_483 = way0_hit ? _GEN_290 : ram_0_28; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_484 = way0_hit ? _GEN_291 : ram_0_29; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_485 = way0_hit ? _GEN_292 : ram_0_30; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_486 = way0_hit ? _GEN_293 : ram_0_31; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_487 = way0_hit ? _GEN_294 : ram_0_32; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_488 = way0_hit ? _GEN_295 : ram_0_33; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_489 = way0_hit ? _GEN_296 : ram_0_34; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_490 = way0_hit ? _GEN_297 : ram_0_35; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_491 = way0_hit ? _GEN_298 : ram_0_36; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_492 = way0_hit ? _GEN_299 : ram_0_37; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_493 = way0_hit ? _GEN_300 : ram_0_38; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_494 = way0_hit ? _GEN_301 : ram_0_39; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_495 = way0_hit ? _GEN_302 : ram_0_40; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_496 = way0_hit ? _GEN_303 : ram_0_41; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_497 = way0_hit ? _GEN_304 : ram_0_42; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_498 = way0_hit ? _GEN_305 : ram_0_43; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_499 = way0_hit ? _GEN_306 : ram_0_44; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_500 = way0_hit ? _GEN_307 : ram_0_45; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_501 = way0_hit ? _GEN_308 : ram_0_46; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_502 = way0_hit ? _GEN_309 : ram_0_47; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_503 = way0_hit ? _GEN_310 : ram_0_48; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_504 = way0_hit ? _GEN_311 : ram_0_49; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_505 = way0_hit ? _GEN_312 : ram_0_50; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_506 = way0_hit ? _GEN_313 : ram_0_51; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_507 = way0_hit ? _GEN_314 : ram_0_52; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_508 = way0_hit ? _GEN_315 : ram_0_53; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_509 = way0_hit ? _GEN_316 : ram_0_54; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_510 = way0_hit ? _GEN_317 : ram_0_55; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_511 = way0_hit ? _GEN_318 : ram_0_56; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_512 = way0_hit ? _GEN_319 : ram_0_57; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_513 = way0_hit ? _GEN_320 : ram_0_58; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_514 = way0_hit ? _GEN_321 : ram_0_59; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_515 = way0_hit ? _GEN_322 : ram_0_60; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_516 = way0_hit ? _GEN_323 : ram_0_61; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_517 = way0_hit ? _GEN_324 : ram_0_62; // @[d_cache.scala 107:27 18:24]
  wire [63:0] _GEN_518 = way0_hit ? _GEN_325 : ram_0_63; // @[d_cache.scala 107:27 18:24]
  wire  _GEN_519 = way0_hit ? _GEN_326 : valid_0_0; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_520 = way0_hit ? _GEN_327 : valid_0_1; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_521 = way0_hit ? _GEN_328 : valid_0_2; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_522 = way0_hit ? _GEN_329 : valid_0_3; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_523 = way0_hit ? _GEN_330 : valid_0_4; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_524 = way0_hit ? _GEN_331 : valid_0_5; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_525 = way0_hit ? _GEN_332 : valid_0_6; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_526 = way0_hit ? _GEN_333 : valid_0_7; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_527 = way0_hit ? _GEN_334 : valid_0_8; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_528 = way0_hit ? _GEN_335 : valid_0_9; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_529 = way0_hit ? _GEN_336 : valid_0_10; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_530 = way0_hit ? _GEN_337 : valid_0_11; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_531 = way0_hit ? _GEN_338 : valid_0_12; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_532 = way0_hit ? _GEN_339 : valid_0_13; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_533 = way0_hit ? _GEN_340 : valid_0_14; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_534 = way0_hit ? _GEN_341 : valid_0_15; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_535 = way0_hit ? _GEN_342 : valid_0_16; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_536 = way0_hit ? _GEN_343 : valid_0_17; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_537 = way0_hit ? _GEN_344 : valid_0_18; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_538 = way0_hit ? _GEN_345 : valid_0_19; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_539 = way0_hit ? _GEN_346 : valid_0_20; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_540 = way0_hit ? _GEN_347 : valid_0_21; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_541 = way0_hit ? _GEN_348 : valid_0_22; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_542 = way0_hit ? _GEN_349 : valid_0_23; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_543 = way0_hit ? _GEN_350 : valid_0_24; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_544 = way0_hit ? _GEN_351 : valid_0_25; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_545 = way0_hit ? _GEN_352 : valid_0_26; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_546 = way0_hit ? _GEN_353 : valid_0_27; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_547 = way0_hit ? _GEN_354 : valid_0_28; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_548 = way0_hit ? _GEN_355 : valid_0_29; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_549 = way0_hit ? _GEN_356 : valid_0_30; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_550 = way0_hit ? _GEN_357 : valid_0_31; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_551 = way0_hit ? _GEN_358 : valid_0_32; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_552 = way0_hit ? _GEN_359 : valid_0_33; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_553 = way0_hit ? _GEN_360 : valid_0_34; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_554 = way0_hit ? _GEN_361 : valid_0_35; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_555 = way0_hit ? _GEN_362 : valid_0_36; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_556 = way0_hit ? _GEN_363 : valid_0_37; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_557 = way0_hit ? _GEN_364 : valid_0_38; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_558 = way0_hit ? _GEN_365 : valid_0_39; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_559 = way0_hit ? _GEN_366 : valid_0_40; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_560 = way0_hit ? _GEN_367 : valid_0_41; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_561 = way0_hit ? _GEN_368 : valid_0_42; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_562 = way0_hit ? _GEN_369 : valid_0_43; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_563 = way0_hit ? _GEN_370 : valid_0_44; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_564 = way0_hit ? _GEN_371 : valid_0_45; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_565 = way0_hit ? _GEN_372 : valid_0_46; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_566 = way0_hit ? _GEN_373 : valid_0_47; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_567 = way0_hit ? _GEN_374 : valid_0_48; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_568 = way0_hit ? _GEN_375 : valid_0_49; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_569 = way0_hit ? _GEN_376 : valid_0_50; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_570 = way0_hit ? _GEN_377 : valid_0_51; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_571 = way0_hit ? _GEN_378 : valid_0_52; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_572 = way0_hit ? _GEN_379 : valid_0_53; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_573 = way0_hit ? _GEN_380 : valid_0_54; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_574 = way0_hit ? _GEN_381 : valid_0_55; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_575 = way0_hit ? _GEN_382 : valid_0_56; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_576 = way0_hit ? _GEN_383 : valid_0_57; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_577 = way0_hit ? _GEN_384 : valid_0_58; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_578 = way0_hit ? _GEN_385 : valid_0_59; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_579 = way0_hit ? _GEN_386 : valid_0_60; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_580 = way0_hit ? _GEN_387 : valid_0_61; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_581 = way0_hit ? _GEN_388 : valid_0_62; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_582 = way0_hit ? _GEN_389 : valid_0_63; // @[d_cache.scala 107:27 24:26]
  wire  _GEN_583 = way0_hit ? _GEN_390 : dirty_0_0; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_584 = way0_hit ? _GEN_391 : dirty_0_1; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_585 = way0_hit ? _GEN_392 : dirty_0_2; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_586 = way0_hit ? _GEN_393 : dirty_0_3; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_587 = way0_hit ? _GEN_394 : dirty_0_4; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_588 = way0_hit ? _GEN_395 : dirty_0_5; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_589 = way0_hit ? _GEN_396 : dirty_0_6; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_590 = way0_hit ? _GEN_397 : dirty_0_7; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_591 = way0_hit ? _GEN_398 : dirty_0_8; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_592 = way0_hit ? _GEN_399 : dirty_0_9; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_593 = way0_hit ? _GEN_400 : dirty_0_10; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_594 = way0_hit ? _GEN_401 : dirty_0_11; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_595 = way0_hit ? _GEN_402 : dirty_0_12; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_596 = way0_hit ? _GEN_403 : dirty_0_13; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_597 = way0_hit ? _GEN_404 : dirty_0_14; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_598 = way0_hit ? _GEN_405 : dirty_0_15; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_599 = way0_hit ? _GEN_406 : dirty_0_16; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_600 = way0_hit ? _GEN_407 : dirty_0_17; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_601 = way0_hit ? _GEN_408 : dirty_0_18; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_602 = way0_hit ? _GEN_409 : dirty_0_19; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_603 = way0_hit ? _GEN_410 : dirty_0_20; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_604 = way0_hit ? _GEN_411 : dirty_0_21; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_605 = way0_hit ? _GEN_412 : dirty_0_22; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_606 = way0_hit ? _GEN_413 : dirty_0_23; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_607 = way0_hit ? _GEN_414 : dirty_0_24; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_608 = way0_hit ? _GEN_415 : dirty_0_25; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_609 = way0_hit ? _GEN_416 : dirty_0_26; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_610 = way0_hit ? _GEN_417 : dirty_0_27; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_611 = way0_hit ? _GEN_418 : dirty_0_28; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_612 = way0_hit ? _GEN_419 : dirty_0_29; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_613 = way0_hit ? _GEN_420 : dirty_0_30; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_614 = way0_hit ? _GEN_421 : dirty_0_31; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_615 = way0_hit ? _GEN_422 : dirty_0_32; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_616 = way0_hit ? _GEN_423 : dirty_0_33; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_617 = way0_hit ? _GEN_424 : dirty_0_34; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_618 = way0_hit ? _GEN_425 : dirty_0_35; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_619 = way0_hit ? _GEN_426 : dirty_0_36; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_620 = way0_hit ? _GEN_427 : dirty_0_37; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_621 = way0_hit ? _GEN_428 : dirty_0_38; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_622 = way0_hit ? _GEN_429 : dirty_0_39; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_623 = way0_hit ? _GEN_430 : dirty_0_40; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_624 = way0_hit ? _GEN_431 : dirty_0_41; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_625 = way0_hit ? _GEN_432 : dirty_0_42; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_626 = way0_hit ? _GEN_433 : dirty_0_43; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_627 = way0_hit ? _GEN_434 : dirty_0_44; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_628 = way0_hit ? _GEN_435 : dirty_0_45; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_629 = way0_hit ? _GEN_436 : dirty_0_46; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_630 = way0_hit ? _GEN_437 : dirty_0_47; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_631 = way0_hit ? _GEN_438 : dirty_0_48; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_632 = way0_hit ? _GEN_439 : dirty_0_49; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_633 = way0_hit ? _GEN_440 : dirty_0_50; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_634 = way0_hit ? _GEN_441 : dirty_0_51; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_635 = way0_hit ? _GEN_442 : dirty_0_52; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_636 = way0_hit ? _GEN_443 : dirty_0_53; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_637 = way0_hit ? _GEN_444 : dirty_0_54; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_638 = way0_hit ? _GEN_445 : dirty_0_55; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_639 = way0_hit ? _GEN_446 : dirty_0_56; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_640 = way0_hit ? _GEN_447 : dirty_0_57; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_641 = way0_hit ? _GEN_448 : dirty_0_58; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_642 = way0_hit ? _GEN_449 : dirty_0_59; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_643 = way0_hit ? _GEN_450 : dirty_0_60; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_644 = way0_hit ? _GEN_451 : dirty_0_61; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_645 = way0_hit ? _GEN_452 : dirty_0_62; // @[d_cache.scala 107:27 26:26]
  wire  _GEN_646 = way0_hit ? _GEN_453 : dirty_0_63; // @[d_cache.scala 107:27 26:26]
  wire [2:0] _GEN_647 = io_from_axi_rvalid ? 3'h5 : state; // @[d_cache.scala 128:37 129:23 76:24]
  wire [63:0] _GEN_648 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[d_cache.scala 131:37 132:30 36:31]
  wire [2:0] _GEN_649 = io_from_axi_bvalid ? 3'h0 : state; // @[d_cache.scala 136:37 137:23 76:24]
  wire [63:0] _GEN_650 = 6'h0 == index ? receive_data : ram_0_0; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_651 = 6'h1 == index ? receive_data : ram_0_1; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_652 = 6'h2 == index ? receive_data : ram_0_2; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_653 = 6'h3 == index ? receive_data : ram_0_3; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_654 = 6'h4 == index ? receive_data : ram_0_4; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_655 = 6'h5 == index ? receive_data : ram_0_5; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_656 = 6'h6 == index ? receive_data : ram_0_6; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_657 = 6'h7 == index ? receive_data : ram_0_7; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_658 = 6'h8 == index ? receive_data : ram_0_8; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_659 = 6'h9 == index ? receive_data : ram_0_9; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_660 = 6'ha == index ? receive_data : ram_0_10; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_661 = 6'hb == index ? receive_data : ram_0_11; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_662 = 6'hc == index ? receive_data : ram_0_12; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_663 = 6'hd == index ? receive_data : ram_0_13; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_664 = 6'he == index ? receive_data : ram_0_14; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_665 = 6'hf == index ? receive_data : ram_0_15; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_666 = 6'h10 == index ? receive_data : ram_0_16; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_667 = 6'h11 == index ? receive_data : ram_0_17; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_668 = 6'h12 == index ? receive_data : ram_0_18; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_669 = 6'h13 == index ? receive_data : ram_0_19; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_670 = 6'h14 == index ? receive_data : ram_0_20; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_671 = 6'h15 == index ? receive_data : ram_0_21; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_672 = 6'h16 == index ? receive_data : ram_0_22; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_673 = 6'h17 == index ? receive_data : ram_0_23; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_674 = 6'h18 == index ? receive_data : ram_0_24; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_675 = 6'h19 == index ? receive_data : ram_0_25; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_676 = 6'h1a == index ? receive_data : ram_0_26; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_677 = 6'h1b == index ? receive_data : ram_0_27; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_678 = 6'h1c == index ? receive_data : ram_0_28; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_679 = 6'h1d == index ? receive_data : ram_0_29; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_680 = 6'h1e == index ? receive_data : ram_0_30; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_681 = 6'h1f == index ? receive_data : ram_0_31; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_682 = 6'h20 == index ? receive_data : ram_0_32; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_683 = 6'h21 == index ? receive_data : ram_0_33; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_684 = 6'h22 == index ? receive_data : ram_0_34; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_685 = 6'h23 == index ? receive_data : ram_0_35; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_686 = 6'h24 == index ? receive_data : ram_0_36; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_687 = 6'h25 == index ? receive_data : ram_0_37; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_688 = 6'h26 == index ? receive_data : ram_0_38; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_689 = 6'h27 == index ? receive_data : ram_0_39; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_690 = 6'h28 == index ? receive_data : ram_0_40; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_691 = 6'h29 == index ? receive_data : ram_0_41; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_692 = 6'h2a == index ? receive_data : ram_0_42; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_693 = 6'h2b == index ? receive_data : ram_0_43; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_694 = 6'h2c == index ? receive_data : ram_0_44; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_695 = 6'h2d == index ? receive_data : ram_0_45; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_696 = 6'h2e == index ? receive_data : ram_0_46; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_697 = 6'h2f == index ? receive_data : ram_0_47; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_698 = 6'h30 == index ? receive_data : ram_0_48; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_699 = 6'h31 == index ? receive_data : ram_0_49; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_700 = 6'h32 == index ? receive_data : ram_0_50; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_701 = 6'h33 == index ? receive_data : ram_0_51; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_702 = 6'h34 == index ? receive_data : ram_0_52; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_703 = 6'h35 == index ? receive_data : ram_0_53; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_704 = 6'h36 == index ? receive_data : ram_0_54; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_705 = 6'h37 == index ? receive_data : ram_0_55; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_706 = 6'h38 == index ? receive_data : ram_0_56; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_707 = 6'h39 == index ? receive_data : ram_0_57; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_708 = 6'h3a == index ? receive_data : ram_0_58; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_709 = 6'h3b == index ? receive_data : ram_0_59; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_710 = 6'h3c == index ? receive_data : ram_0_60; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_711 = 6'h3d == index ? receive_data : ram_0_61; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_712 = 6'h3e == index ? receive_data : ram_0_62; // @[d_cache.scala 143:{30,30} 18:24]
  wire [63:0] _GEN_713 = 6'h3f == index ? receive_data : ram_0_63; // @[d_cache.scala 143:{30,30} 18:24]
  wire [31:0] _GEN_714 = 6'h0 == index ? _GEN_3460 : tag_0_0; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_715 = 6'h1 == index ? _GEN_3460 : tag_0_1; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_716 = 6'h2 == index ? _GEN_3460 : tag_0_2; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_717 = 6'h3 == index ? _GEN_3460 : tag_0_3; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_718 = 6'h4 == index ? _GEN_3460 : tag_0_4; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_719 = 6'h5 == index ? _GEN_3460 : tag_0_5; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_720 = 6'h6 == index ? _GEN_3460 : tag_0_6; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_721 = 6'h7 == index ? _GEN_3460 : tag_0_7; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_722 = 6'h8 == index ? _GEN_3460 : tag_0_8; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_723 = 6'h9 == index ? _GEN_3460 : tag_0_9; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_724 = 6'ha == index ? _GEN_3460 : tag_0_10; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_725 = 6'hb == index ? _GEN_3460 : tag_0_11; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_726 = 6'hc == index ? _GEN_3460 : tag_0_12; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_727 = 6'hd == index ? _GEN_3460 : tag_0_13; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_728 = 6'he == index ? _GEN_3460 : tag_0_14; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_729 = 6'hf == index ? _GEN_3460 : tag_0_15; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_730 = 6'h10 == index ? _GEN_3460 : tag_0_16; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_731 = 6'h11 == index ? _GEN_3460 : tag_0_17; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_732 = 6'h12 == index ? _GEN_3460 : tag_0_18; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_733 = 6'h13 == index ? _GEN_3460 : tag_0_19; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_734 = 6'h14 == index ? _GEN_3460 : tag_0_20; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_735 = 6'h15 == index ? _GEN_3460 : tag_0_21; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_736 = 6'h16 == index ? _GEN_3460 : tag_0_22; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_737 = 6'h17 == index ? _GEN_3460 : tag_0_23; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_738 = 6'h18 == index ? _GEN_3460 : tag_0_24; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_739 = 6'h19 == index ? _GEN_3460 : tag_0_25; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_740 = 6'h1a == index ? _GEN_3460 : tag_0_26; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_741 = 6'h1b == index ? _GEN_3460 : tag_0_27; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_742 = 6'h1c == index ? _GEN_3460 : tag_0_28; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_743 = 6'h1d == index ? _GEN_3460 : tag_0_29; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_744 = 6'h1e == index ? _GEN_3460 : tag_0_30; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_745 = 6'h1f == index ? _GEN_3460 : tag_0_31; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_746 = 6'h20 == index ? _GEN_3460 : tag_0_32; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_747 = 6'h21 == index ? _GEN_3460 : tag_0_33; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_748 = 6'h22 == index ? _GEN_3460 : tag_0_34; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_749 = 6'h23 == index ? _GEN_3460 : tag_0_35; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_750 = 6'h24 == index ? _GEN_3460 : tag_0_36; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_751 = 6'h25 == index ? _GEN_3460 : tag_0_37; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_752 = 6'h26 == index ? _GEN_3460 : tag_0_38; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_753 = 6'h27 == index ? _GEN_3460 : tag_0_39; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_754 = 6'h28 == index ? _GEN_3460 : tag_0_40; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_755 = 6'h29 == index ? _GEN_3460 : tag_0_41; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_756 = 6'h2a == index ? _GEN_3460 : tag_0_42; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_757 = 6'h2b == index ? _GEN_3460 : tag_0_43; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_758 = 6'h2c == index ? _GEN_3460 : tag_0_44; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_759 = 6'h2d == index ? _GEN_3460 : tag_0_45; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_760 = 6'h2e == index ? _GEN_3460 : tag_0_46; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_761 = 6'h2f == index ? _GEN_3460 : tag_0_47; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_762 = 6'h30 == index ? _GEN_3460 : tag_0_48; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_763 = 6'h31 == index ? _GEN_3460 : tag_0_49; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_764 = 6'h32 == index ? _GEN_3460 : tag_0_50; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_765 = 6'h33 == index ? _GEN_3460 : tag_0_51; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_766 = 6'h34 == index ? _GEN_3460 : tag_0_52; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_767 = 6'h35 == index ? _GEN_3460 : tag_0_53; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_768 = 6'h36 == index ? _GEN_3460 : tag_0_54; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_769 = 6'h37 == index ? _GEN_3460 : tag_0_55; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_770 = 6'h38 == index ? _GEN_3460 : tag_0_56; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_771 = 6'h39 == index ? _GEN_3460 : tag_0_57; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_772 = 6'h3a == index ? _GEN_3460 : tag_0_58; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_773 = 6'h3b == index ? _GEN_3460 : tag_0_59; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_774 = 6'h3c == index ? _GEN_3460 : tag_0_60; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_775 = 6'h3d == index ? _GEN_3460 : tag_0_61; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_776 = 6'h3e == index ? _GEN_3460 : tag_0_62; // @[d_cache.scala 144:{30,30} 22:24]
  wire [31:0] _GEN_777 = 6'h3f == index ? _GEN_3460 : tag_0_63; // @[d_cache.scala 144:{30,30} 22:24]
  wire [40:0] _write_back_addr_T_1 = {_GEN_63,index,3'h0}; // @[Cat.scala 31:58]
  wire  _GEN_970 = 6'h0 == index ? 1'h0 : dirty_0_0; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_971 = 6'h1 == index ? 1'h0 : dirty_0_1; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_972 = 6'h2 == index ? 1'h0 : dirty_0_2; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_973 = 6'h3 == index ? 1'h0 : dirty_0_3; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_974 = 6'h4 == index ? 1'h0 : dirty_0_4; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_975 = 6'h5 == index ? 1'h0 : dirty_0_5; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_976 = 6'h6 == index ? 1'h0 : dirty_0_6; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_977 = 6'h7 == index ? 1'h0 : dirty_0_7; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_978 = 6'h8 == index ? 1'h0 : dirty_0_8; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_979 = 6'h9 == index ? 1'h0 : dirty_0_9; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_980 = 6'ha == index ? 1'h0 : dirty_0_10; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_981 = 6'hb == index ? 1'h0 : dirty_0_11; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_982 = 6'hc == index ? 1'h0 : dirty_0_12; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_983 = 6'hd == index ? 1'h0 : dirty_0_13; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_984 = 6'he == index ? 1'h0 : dirty_0_14; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_985 = 6'hf == index ? 1'h0 : dirty_0_15; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_986 = 6'h10 == index ? 1'h0 : dirty_0_16; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_987 = 6'h11 == index ? 1'h0 : dirty_0_17; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_988 = 6'h12 == index ? 1'h0 : dirty_0_18; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_989 = 6'h13 == index ? 1'h0 : dirty_0_19; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_990 = 6'h14 == index ? 1'h0 : dirty_0_20; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_991 = 6'h15 == index ? 1'h0 : dirty_0_21; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_992 = 6'h16 == index ? 1'h0 : dirty_0_22; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_993 = 6'h17 == index ? 1'h0 : dirty_0_23; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_994 = 6'h18 == index ? 1'h0 : dirty_0_24; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_995 = 6'h19 == index ? 1'h0 : dirty_0_25; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_996 = 6'h1a == index ? 1'h0 : dirty_0_26; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_997 = 6'h1b == index ? 1'h0 : dirty_0_27; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_998 = 6'h1c == index ? 1'h0 : dirty_0_28; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_999 = 6'h1d == index ? 1'h0 : dirty_0_29; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1000 = 6'h1e == index ? 1'h0 : dirty_0_30; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1001 = 6'h1f == index ? 1'h0 : dirty_0_31; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1002 = 6'h20 == index ? 1'h0 : dirty_0_32; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1003 = 6'h21 == index ? 1'h0 : dirty_0_33; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1004 = 6'h22 == index ? 1'h0 : dirty_0_34; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1005 = 6'h23 == index ? 1'h0 : dirty_0_35; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1006 = 6'h24 == index ? 1'h0 : dirty_0_36; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1007 = 6'h25 == index ? 1'h0 : dirty_0_37; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1008 = 6'h26 == index ? 1'h0 : dirty_0_38; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1009 = 6'h27 == index ? 1'h0 : dirty_0_39; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1010 = 6'h28 == index ? 1'h0 : dirty_0_40; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1011 = 6'h29 == index ? 1'h0 : dirty_0_41; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1012 = 6'h2a == index ? 1'h0 : dirty_0_42; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1013 = 6'h2b == index ? 1'h0 : dirty_0_43; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1014 = 6'h2c == index ? 1'h0 : dirty_0_44; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1015 = 6'h2d == index ? 1'h0 : dirty_0_45; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1016 = 6'h2e == index ? 1'h0 : dirty_0_46; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1017 = 6'h2f == index ? 1'h0 : dirty_0_47; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1018 = 6'h30 == index ? 1'h0 : dirty_0_48; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1019 = 6'h31 == index ? 1'h0 : dirty_0_49; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1020 = 6'h32 == index ? 1'h0 : dirty_0_50; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1021 = 6'h33 == index ? 1'h0 : dirty_0_51; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1022 = 6'h34 == index ? 1'h0 : dirty_0_52; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1023 = 6'h35 == index ? 1'h0 : dirty_0_53; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1024 = 6'h36 == index ? 1'h0 : dirty_0_54; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1025 = 6'h37 == index ? 1'h0 : dirty_0_55; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1026 = 6'h38 == index ? 1'h0 : dirty_0_56; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1027 = 6'h39 == index ? 1'h0 : dirty_0_57; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1028 = 6'h3a == index ? 1'h0 : dirty_0_58; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1029 = 6'h3b == index ? 1'h0 : dirty_0_59; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1030 = 6'h3c == index ? 1'h0 : dirty_0_60; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1031 = 6'h3d == index ? 1'h0 : dirty_0_61; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1032 = 6'h3e == index ? 1'h0 : dirty_0_62; // @[d_cache.scala 161:{40,40} 26:26]
  wire  _GEN_1033 = 6'h3f == index ? 1'h0 : dirty_0_63; // @[d_cache.scala 161:{40,40} 26:26]
  wire [63:0] _GEN_1290 = _GEN_195 ? _GEN_261 : write_back_data; // @[d_cache.scala 156:47 157:41 31:34]
  wire [40:0] _GEN_1291 = _GEN_195 ? _write_back_addr_T_1 : {{9'd0}, write_back_addr}; // @[d_cache.scala 156:47 158:41 32:34]
  wire [63:0] _GEN_1292 = _GEN_195 ? _GEN_650 : _GEN_650; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1293 = _GEN_195 ? _GEN_651 : _GEN_651; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1294 = _GEN_195 ? _GEN_652 : _GEN_652; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1295 = _GEN_195 ? _GEN_653 : _GEN_653; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1296 = _GEN_195 ? _GEN_654 : _GEN_654; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1297 = _GEN_195 ? _GEN_655 : _GEN_655; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1298 = _GEN_195 ? _GEN_656 : _GEN_656; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1299 = _GEN_195 ? _GEN_657 : _GEN_657; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1300 = _GEN_195 ? _GEN_658 : _GEN_658; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1301 = _GEN_195 ? _GEN_659 : _GEN_659; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1302 = _GEN_195 ? _GEN_660 : _GEN_660; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1303 = _GEN_195 ? _GEN_661 : _GEN_661; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1304 = _GEN_195 ? _GEN_662 : _GEN_662; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1305 = _GEN_195 ? _GEN_663 : _GEN_663; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1306 = _GEN_195 ? _GEN_664 : _GEN_664; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1307 = _GEN_195 ? _GEN_665 : _GEN_665; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1308 = _GEN_195 ? _GEN_666 : _GEN_666; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1309 = _GEN_195 ? _GEN_667 : _GEN_667; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1310 = _GEN_195 ? _GEN_668 : _GEN_668; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1311 = _GEN_195 ? _GEN_669 : _GEN_669; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1312 = _GEN_195 ? _GEN_670 : _GEN_670; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1313 = _GEN_195 ? _GEN_671 : _GEN_671; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1314 = _GEN_195 ? _GEN_672 : _GEN_672; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1315 = _GEN_195 ? _GEN_673 : _GEN_673; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1316 = _GEN_195 ? _GEN_674 : _GEN_674; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1317 = _GEN_195 ? _GEN_675 : _GEN_675; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1318 = _GEN_195 ? _GEN_676 : _GEN_676; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1319 = _GEN_195 ? _GEN_677 : _GEN_677; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1320 = _GEN_195 ? _GEN_678 : _GEN_678; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1321 = _GEN_195 ? _GEN_679 : _GEN_679; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1322 = _GEN_195 ? _GEN_680 : _GEN_680; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1323 = _GEN_195 ? _GEN_681 : _GEN_681; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1324 = _GEN_195 ? _GEN_682 : _GEN_682; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1325 = _GEN_195 ? _GEN_683 : _GEN_683; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1326 = _GEN_195 ? _GEN_684 : _GEN_684; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1327 = _GEN_195 ? _GEN_685 : _GEN_685; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1328 = _GEN_195 ? _GEN_686 : _GEN_686; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1329 = _GEN_195 ? _GEN_687 : _GEN_687; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1330 = _GEN_195 ? _GEN_688 : _GEN_688; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1331 = _GEN_195 ? _GEN_689 : _GEN_689; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1332 = _GEN_195 ? _GEN_690 : _GEN_690; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1333 = _GEN_195 ? _GEN_691 : _GEN_691; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1334 = _GEN_195 ? _GEN_692 : _GEN_692; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1335 = _GEN_195 ? _GEN_693 : _GEN_693; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1336 = _GEN_195 ? _GEN_694 : _GEN_694; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1337 = _GEN_195 ? _GEN_695 : _GEN_695; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1338 = _GEN_195 ? _GEN_696 : _GEN_696; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1339 = _GEN_195 ? _GEN_697 : _GEN_697; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1340 = _GEN_195 ? _GEN_698 : _GEN_698; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1341 = _GEN_195 ? _GEN_699 : _GEN_699; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1342 = _GEN_195 ? _GEN_700 : _GEN_700; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1343 = _GEN_195 ? _GEN_701 : _GEN_701; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1344 = _GEN_195 ? _GEN_702 : _GEN_702; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1345 = _GEN_195 ? _GEN_703 : _GEN_703; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1346 = _GEN_195 ? _GEN_704 : _GEN_704; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1347 = _GEN_195 ? _GEN_705 : _GEN_705; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1348 = _GEN_195 ? _GEN_706 : _GEN_706; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1349 = _GEN_195 ? _GEN_707 : _GEN_707; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1350 = _GEN_195 ? _GEN_708 : _GEN_708; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1351 = _GEN_195 ? _GEN_709 : _GEN_709; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1352 = _GEN_195 ? _GEN_710 : _GEN_710; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1353 = _GEN_195 ? _GEN_711 : _GEN_711; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1354 = _GEN_195 ? _GEN_712 : _GEN_712; // @[d_cache.scala 156:47]
  wire [63:0] _GEN_1355 = _GEN_195 ? _GEN_713 : _GEN_713; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1356 = _GEN_195 ? _GEN_714 : _GEN_714; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1357 = _GEN_195 ? _GEN_715 : _GEN_715; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1358 = _GEN_195 ? _GEN_716 : _GEN_716; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1359 = _GEN_195 ? _GEN_717 : _GEN_717; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1360 = _GEN_195 ? _GEN_718 : _GEN_718; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1361 = _GEN_195 ? _GEN_719 : _GEN_719; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1362 = _GEN_195 ? _GEN_720 : _GEN_720; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1363 = _GEN_195 ? _GEN_721 : _GEN_721; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1364 = _GEN_195 ? _GEN_722 : _GEN_722; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1365 = _GEN_195 ? _GEN_723 : _GEN_723; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1366 = _GEN_195 ? _GEN_724 : _GEN_724; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1367 = _GEN_195 ? _GEN_725 : _GEN_725; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1368 = _GEN_195 ? _GEN_726 : _GEN_726; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1369 = _GEN_195 ? _GEN_727 : _GEN_727; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1370 = _GEN_195 ? _GEN_728 : _GEN_728; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1371 = _GEN_195 ? _GEN_729 : _GEN_729; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1372 = _GEN_195 ? _GEN_730 : _GEN_730; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1373 = _GEN_195 ? _GEN_731 : _GEN_731; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1374 = _GEN_195 ? _GEN_732 : _GEN_732; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1375 = _GEN_195 ? _GEN_733 : _GEN_733; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1376 = _GEN_195 ? _GEN_734 : _GEN_734; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1377 = _GEN_195 ? _GEN_735 : _GEN_735; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1378 = _GEN_195 ? _GEN_736 : _GEN_736; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1379 = _GEN_195 ? _GEN_737 : _GEN_737; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1380 = _GEN_195 ? _GEN_738 : _GEN_738; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1381 = _GEN_195 ? _GEN_739 : _GEN_739; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1382 = _GEN_195 ? _GEN_740 : _GEN_740; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1383 = _GEN_195 ? _GEN_741 : _GEN_741; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1384 = _GEN_195 ? _GEN_742 : _GEN_742; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1385 = _GEN_195 ? _GEN_743 : _GEN_743; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1386 = _GEN_195 ? _GEN_744 : _GEN_744; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1387 = _GEN_195 ? _GEN_745 : _GEN_745; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1388 = _GEN_195 ? _GEN_746 : _GEN_746; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1389 = _GEN_195 ? _GEN_747 : _GEN_747; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1390 = _GEN_195 ? _GEN_748 : _GEN_748; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1391 = _GEN_195 ? _GEN_749 : _GEN_749; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1392 = _GEN_195 ? _GEN_750 : _GEN_750; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1393 = _GEN_195 ? _GEN_751 : _GEN_751; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1394 = _GEN_195 ? _GEN_752 : _GEN_752; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1395 = _GEN_195 ? _GEN_753 : _GEN_753; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1396 = _GEN_195 ? _GEN_754 : _GEN_754; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1397 = _GEN_195 ? _GEN_755 : _GEN_755; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1398 = _GEN_195 ? _GEN_756 : _GEN_756; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1399 = _GEN_195 ? _GEN_757 : _GEN_757; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1400 = _GEN_195 ? _GEN_758 : _GEN_758; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1401 = _GEN_195 ? _GEN_759 : _GEN_759; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1402 = _GEN_195 ? _GEN_760 : _GEN_760; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1403 = _GEN_195 ? _GEN_761 : _GEN_761; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1404 = _GEN_195 ? _GEN_762 : _GEN_762; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1405 = _GEN_195 ? _GEN_763 : _GEN_763; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1406 = _GEN_195 ? _GEN_764 : _GEN_764; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1407 = _GEN_195 ? _GEN_765 : _GEN_765; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1408 = _GEN_195 ? _GEN_766 : _GEN_766; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1409 = _GEN_195 ? _GEN_767 : _GEN_767; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1410 = _GEN_195 ? _GEN_768 : _GEN_768; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1411 = _GEN_195 ? _GEN_769 : _GEN_769; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1412 = _GEN_195 ? _GEN_770 : _GEN_770; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1413 = _GEN_195 ? _GEN_771 : _GEN_771; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1414 = _GEN_195 ? _GEN_772 : _GEN_772; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1415 = _GEN_195 ? _GEN_773 : _GEN_773; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1416 = _GEN_195 ? _GEN_774 : _GEN_774; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1417 = _GEN_195 ? _GEN_775 : _GEN_775; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1418 = _GEN_195 ? _GEN_776 : _GEN_776; // @[d_cache.scala 156:47]
  wire [31:0] _GEN_1419 = _GEN_195 ? _GEN_777 : _GEN_777; // @[d_cache.scala 156:47]
  wire  _GEN_1420 = _GEN_195 ? _GEN_970 : dirty_0_0; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1421 = _GEN_195 ? _GEN_971 : dirty_0_1; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1422 = _GEN_195 ? _GEN_972 : dirty_0_2; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1423 = _GEN_195 ? _GEN_973 : dirty_0_3; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1424 = _GEN_195 ? _GEN_974 : dirty_0_4; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1425 = _GEN_195 ? _GEN_975 : dirty_0_5; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1426 = _GEN_195 ? _GEN_976 : dirty_0_6; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1427 = _GEN_195 ? _GEN_977 : dirty_0_7; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1428 = _GEN_195 ? _GEN_978 : dirty_0_8; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1429 = _GEN_195 ? _GEN_979 : dirty_0_9; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1430 = _GEN_195 ? _GEN_980 : dirty_0_10; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1431 = _GEN_195 ? _GEN_981 : dirty_0_11; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1432 = _GEN_195 ? _GEN_982 : dirty_0_12; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1433 = _GEN_195 ? _GEN_983 : dirty_0_13; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1434 = _GEN_195 ? _GEN_984 : dirty_0_14; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1435 = _GEN_195 ? _GEN_985 : dirty_0_15; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1436 = _GEN_195 ? _GEN_986 : dirty_0_16; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1437 = _GEN_195 ? _GEN_987 : dirty_0_17; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1438 = _GEN_195 ? _GEN_988 : dirty_0_18; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1439 = _GEN_195 ? _GEN_989 : dirty_0_19; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1440 = _GEN_195 ? _GEN_990 : dirty_0_20; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1441 = _GEN_195 ? _GEN_991 : dirty_0_21; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1442 = _GEN_195 ? _GEN_992 : dirty_0_22; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1443 = _GEN_195 ? _GEN_993 : dirty_0_23; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1444 = _GEN_195 ? _GEN_994 : dirty_0_24; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1445 = _GEN_195 ? _GEN_995 : dirty_0_25; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1446 = _GEN_195 ? _GEN_996 : dirty_0_26; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1447 = _GEN_195 ? _GEN_997 : dirty_0_27; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1448 = _GEN_195 ? _GEN_998 : dirty_0_28; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1449 = _GEN_195 ? _GEN_999 : dirty_0_29; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1450 = _GEN_195 ? _GEN_1000 : dirty_0_30; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1451 = _GEN_195 ? _GEN_1001 : dirty_0_31; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1452 = _GEN_195 ? _GEN_1002 : dirty_0_32; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1453 = _GEN_195 ? _GEN_1003 : dirty_0_33; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1454 = _GEN_195 ? _GEN_1004 : dirty_0_34; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1455 = _GEN_195 ? _GEN_1005 : dirty_0_35; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1456 = _GEN_195 ? _GEN_1006 : dirty_0_36; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1457 = _GEN_195 ? _GEN_1007 : dirty_0_37; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1458 = _GEN_195 ? _GEN_1008 : dirty_0_38; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1459 = _GEN_195 ? _GEN_1009 : dirty_0_39; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1460 = _GEN_195 ? _GEN_1010 : dirty_0_40; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1461 = _GEN_195 ? _GEN_1011 : dirty_0_41; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1462 = _GEN_195 ? _GEN_1012 : dirty_0_42; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1463 = _GEN_195 ? _GEN_1013 : dirty_0_43; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1464 = _GEN_195 ? _GEN_1014 : dirty_0_44; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1465 = _GEN_195 ? _GEN_1015 : dirty_0_45; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1466 = _GEN_195 ? _GEN_1016 : dirty_0_46; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1467 = _GEN_195 ? _GEN_1017 : dirty_0_47; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1468 = _GEN_195 ? _GEN_1018 : dirty_0_48; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1469 = _GEN_195 ? _GEN_1019 : dirty_0_49; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1470 = _GEN_195 ? _GEN_1020 : dirty_0_50; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1471 = _GEN_195 ? _GEN_1021 : dirty_0_51; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1472 = _GEN_195 ? _GEN_1022 : dirty_0_52; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1473 = _GEN_195 ? _GEN_1023 : dirty_0_53; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1474 = _GEN_195 ? _GEN_1024 : dirty_0_54; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1475 = _GEN_195 ? _GEN_1025 : dirty_0_55; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1476 = _GEN_195 ? _GEN_1026 : dirty_0_56; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1477 = _GEN_195 ? _GEN_1027 : dirty_0_57; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1478 = _GEN_195 ? _GEN_1028 : dirty_0_58; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1479 = _GEN_195 ? _GEN_1029 : dirty_0_59; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1480 = _GEN_195 ? _GEN_1030 : dirty_0_60; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1481 = _GEN_195 ? _GEN_1031 : dirty_0_61; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1482 = _GEN_195 ? _GEN_1032 : dirty_0_62; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1483 = _GEN_195 ? _GEN_1033 : dirty_0_63; // @[d_cache.scala 156:47 26:26]
  wire  _GEN_1484 = _GEN_195 ? _GEN_326 : _GEN_326; // @[d_cache.scala 156:47]
  wire  _GEN_1485 = _GEN_195 ? _GEN_327 : _GEN_327; // @[d_cache.scala 156:47]
  wire  _GEN_1486 = _GEN_195 ? _GEN_328 : _GEN_328; // @[d_cache.scala 156:47]
  wire  _GEN_1487 = _GEN_195 ? _GEN_329 : _GEN_329; // @[d_cache.scala 156:47]
  wire  _GEN_1488 = _GEN_195 ? _GEN_330 : _GEN_330; // @[d_cache.scala 156:47]
  wire  _GEN_1489 = _GEN_195 ? _GEN_331 : _GEN_331; // @[d_cache.scala 156:47]
  wire  _GEN_1490 = _GEN_195 ? _GEN_332 : _GEN_332; // @[d_cache.scala 156:47]
  wire  _GEN_1491 = _GEN_195 ? _GEN_333 : _GEN_333; // @[d_cache.scala 156:47]
  wire  _GEN_1492 = _GEN_195 ? _GEN_334 : _GEN_334; // @[d_cache.scala 156:47]
  wire  _GEN_1493 = _GEN_195 ? _GEN_335 : _GEN_335; // @[d_cache.scala 156:47]
  wire  _GEN_1494 = _GEN_195 ? _GEN_336 : _GEN_336; // @[d_cache.scala 156:47]
  wire  _GEN_1495 = _GEN_195 ? _GEN_337 : _GEN_337; // @[d_cache.scala 156:47]
  wire  _GEN_1496 = _GEN_195 ? _GEN_338 : _GEN_338; // @[d_cache.scala 156:47]
  wire  _GEN_1497 = _GEN_195 ? _GEN_339 : _GEN_339; // @[d_cache.scala 156:47]
  wire  _GEN_1498 = _GEN_195 ? _GEN_340 : _GEN_340; // @[d_cache.scala 156:47]
  wire  _GEN_1499 = _GEN_195 ? _GEN_341 : _GEN_341; // @[d_cache.scala 156:47]
  wire  _GEN_1500 = _GEN_195 ? _GEN_342 : _GEN_342; // @[d_cache.scala 156:47]
  wire  _GEN_1501 = _GEN_195 ? _GEN_343 : _GEN_343; // @[d_cache.scala 156:47]
  wire  _GEN_1502 = _GEN_195 ? _GEN_344 : _GEN_344; // @[d_cache.scala 156:47]
  wire  _GEN_1503 = _GEN_195 ? _GEN_345 : _GEN_345; // @[d_cache.scala 156:47]
  wire  _GEN_1504 = _GEN_195 ? _GEN_346 : _GEN_346; // @[d_cache.scala 156:47]
  wire  _GEN_1505 = _GEN_195 ? _GEN_347 : _GEN_347; // @[d_cache.scala 156:47]
  wire  _GEN_1506 = _GEN_195 ? _GEN_348 : _GEN_348; // @[d_cache.scala 156:47]
  wire  _GEN_1507 = _GEN_195 ? _GEN_349 : _GEN_349; // @[d_cache.scala 156:47]
  wire  _GEN_1508 = _GEN_195 ? _GEN_350 : _GEN_350; // @[d_cache.scala 156:47]
  wire  _GEN_1509 = _GEN_195 ? _GEN_351 : _GEN_351; // @[d_cache.scala 156:47]
  wire  _GEN_1510 = _GEN_195 ? _GEN_352 : _GEN_352; // @[d_cache.scala 156:47]
  wire  _GEN_1511 = _GEN_195 ? _GEN_353 : _GEN_353; // @[d_cache.scala 156:47]
  wire  _GEN_1512 = _GEN_195 ? _GEN_354 : _GEN_354; // @[d_cache.scala 156:47]
  wire  _GEN_1513 = _GEN_195 ? _GEN_355 : _GEN_355; // @[d_cache.scala 156:47]
  wire  _GEN_1514 = _GEN_195 ? _GEN_356 : _GEN_356; // @[d_cache.scala 156:47]
  wire  _GEN_1515 = _GEN_195 ? _GEN_357 : _GEN_357; // @[d_cache.scala 156:47]
  wire  _GEN_1516 = _GEN_195 ? _GEN_358 : _GEN_358; // @[d_cache.scala 156:47]
  wire  _GEN_1517 = _GEN_195 ? _GEN_359 : _GEN_359; // @[d_cache.scala 156:47]
  wire  _GEN_1518 = _GEN_195 ? _GEN_360 : _GEN_360; // @[d_cache.scala 156:47]
  wire  _GEN_1519 = _GEN_195 ? _GEN_361 : _GEN_361; // @[d_cache.scala 156:47]
  wire  _GEN_1520 = _GEN_195 ? _GEN_362 : _GEN_362; // @[d_cache.scala 156:47]
  wire  _GEN_1521 = _GEN_195 ? _GEN_363 : _GEN_363; // @[d_cache.scala 156:47]
  wire  _GEN_1522 = _GEN_195 ? _GEN_364 : _GEN_364; // @[d_cache.scala 156:47]
  wire  _GEN_1523 = _GEN_195 ? _GEN_365 : _GEN_365; // @[d_cache.scala 156:47]
  wire  _GEN_1524 = _GEN_195 ? _GEN_366 : _GEN_366; // @[d_cache.scala 156:47]
  wire  _GEN_1525 = _GEN_195 ? _GEN_367 : _GEN_367; // @[d_cache.scala 156:47]
  wire  _GEN_1526 = _GEN_195 ? _GEN_368 : _GEN_368; // @[d_cache.scala 156:47]
  wire  _GEN_1527 = _GEN_195 ? _GEN_369 : _GEN_369; // @[d_cache.scala 156:47]
  wire  _GEN_1528 = _GEN_195 ? _GEN_370 : _GEN_370; // @[d_cache.scala 156:47]
  wire  _GEN_1529 = _GEN_195 ? _GEN_371 : _GEN_371; // @[d_cache.scala 156:47]
  wire  _GEN_1530 = _GEN_195 ? _GEN_372 : _GEN_372; // @[d_cache.scala 156:47]
  wire  _GEN_1531 = _GEN_195 ? _GEN_373 : _GEN_373; // @[d_cache.scala 156:47]
  wire  _GEN_1532 = _GEN_195 ? _GEN_374 : _GEN_374; // @[d_cache.scala 156:47]
  wire  _GEN_1533 = _GEN_195 ? _GEN_375 : _GEN_375; // @[d_cache.scala 156:47]
  wire  _GEN_1534 = _GEN_195 ? _GEN_376 : _GEN_376; // @[d_cache.scala 156:47]
  wire  _GEN_1535 = _GEN_195 ? _GEN_377 : _GEN_377; // @[d_cache.scala 156:47]
  wire  _GEN_1536 = _GEN_195 ? _GEN_378 : _GEN_378; // @[d_cache.scala 156:47]
  wire  _GEN_1537 = _GEN_195 ? _GEN_379 : _GEN_379; // @[d_cache.scala 156:47]
  wire  _GEN_1538 = _GEN_195 ? _GEN_380 : _GEN_380; // @[d_cache.scala 156:47]
  wire  _GEN_1539 = _GEN_195 ? _GEN_381 : _GEN_381; // @[d_cache.scala 156:47]
  wire  _GEN_1540 = _GEN_195 ? _GEN_382 : _GEN_382; // @[d_cache.scala 156:47]
  wire  _GEN_1541 = _GEN_195 ? _GEN_383 : _GEN_383; // @[d_cache.scala 156:47]
  wire  _GEN_1542 = _GEN_195 ? _GEN_384 : _GEN_384; // @[d_cache.scala 156:47]
  wire  _GEN_1543 = _GEN_195 ? _GEN_385 : _GEN_385; // @[d_cache.scala 156:47]
  wire  _GEN_1544 = _GEN_195 ? _GEN_386 : _GEN_386; // @[d_cache.scala 156:47]
  wire  _GEN_1545 = _GEN_195 ? _GEN_387 : _GEN_387; // @[d_cache.scala 156:47]
  wire  _GEN_1546 = _GEN_195 ? _GEN_388 : _GEN_388; // @[d_cache.scala 156:47]
  wire  _GEN_1547 = _GEN_195 ? _GEN_389 : _GEN_389; // @[d_cache.scala 156:47]
  wire [2:0] _GEN_1548 = _GEN_195 ? 3'h6 : 3'h7; // @[d_cache.scala 156:47 163:31 166:31]
  wire [2:0] _GEN_1549 = unuse_way == 2'h1 ? 3'h7 : _GEN_1548; // @[d_cache.scala 141:34 142:23]
  wire [63:0] _GEN_1550 = unuse_way == 2'h1 ? _GEN_650 : _GEN_1292; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1551 = unuse_way == 2'h1 ? _GEN_651 : _GEN_1293; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1552 = unuse_way == 2'h1 ? _GEN_652 : _GEN_1294; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1553 = unuse_way == 2'h1 ? _GEN_653 : _GEN_1295; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1554 = unuse_way == 2'h1 ? _GEN_654 : _GEN_1296; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1555 = unuse_way == 2'h1 ? _GEN_655 : _GEN_1297; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1556 = unuse_way == 2'h1 ? _GEN_656 : _GEN_1298; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1557 = unuse_way == 2'h1 ? _GEN_657 : _GEN_1299; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1558 = unuse_way == 2'h1 ? _GEN_658 : _GEN_1300; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1559 = unuse_way == 2'h1 ? _GEN_659 : _GEN_1301; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1560 = unuse_way == 2'h1 ? _GEN_660 : _GEN_1302; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1561 = unuse_way == 2'h1 ? _GEN_661 : _GEN_1303; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1562 = unuse_way == 2'h1 ? _GEN_662 : _GEN_1304; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1563 = unuse_way == 2'h1 ? _GEN_663 : _GEN_1305; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1564 = unuse_way == 2'h1 ? _GEN_664 : _GEN_1306; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1565 = unuse_way == 2'h1 ? _GEN_665 : _GEN_1307; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1566 = unuse_way == 2'h1 ? _GEN_666 : _GEN_1308; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1567 = unuse_way == 2'h1 ? _GEN_667 : _GEN_1309; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1568 = unuse_way == 2'h1 ? _GEN_668 : _GEN_1310; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1569 = unuse_way == 2'h1 ? _GEN_669 : _GEN_1311; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1570 = unuse_way == 2'h1 ? _GEN_670 : _GEN_1312; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1571 = unuse_way == 2'h1 ? _GEN_671 : _GEN_1313; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1572 = unuse_way == 2'h1 ? _GEN_672 : _GEN_1314; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1573 = unuse_way == 2'h1 ? _GEN_673 : _GEN_1315; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1574 = unuse_way == 2'h1 ? _GEN_674 : _GEN_1316; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1575 = unuse_way == 2'h1 ? _GEN_675 : _GEN_1317; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1576 = unuse_way == 2'h1 ? _GEN_676 : _GEN_1318; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1577 = unuse_way == 2'h1 ? _GEN_677 : _GEN_1319; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1578 = unuse_way == 2'h1 ? _GEN_678 : _GEN_1320; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1579 = unuse_way == 2'h1 ? _GEN_679 : _GEN_1321; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1580 = unuse_way == 2'h1 ? _GEN_680 : _GEN_1322; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1581 = unuse_way == 2'h1 ? _GEN_681 : _GEN_1323; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1582 = unuse_way == 2'h1 ? _GEN_682 : _GEN_1324; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1583 = unuse_way == 2'h1 ? _GEN_683 : _GEN_1325; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1584 = unuse_way == 2'h1 ? _GEN_684 : _GEN_1326; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1585 = unuse_way == 2'h1 ? _GEN_685 : _GEN_1327; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1586 = unuse_way == 2'h1 ? _GEN_686 : _GEN_1328; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1587 = unuse_way == 2'h1 ? _GEN_687 : _GEN_1329; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1588 = unuse_way == 2'h1 ? _GEN_688 : _GEN_1330; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1589 = unuse_way == 2'h1 ? _GEN_689 : _GEN_1331; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1590 = unuse_way == 2'h1 ? _GEN_690 : _GEN_1332; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1591 = unuse_way == 2'h1 ? _GEN_691 : _GEN_1333; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1592 = unuse_way == 2'h1 ? _GEN_692 : _GEN_1334; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1593 = unuse_way == 2'h1 ? _GEN_693 : _GEN_1335; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1594 = unuse_way == 2'h1 ? _GEN_694 : _GEN_1336; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1595 = unuse_way == 2'h1 ? _GEN_695 : _GEN_1337; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1596 = unuse_way == 2'h1 ? _GEN_696 : _GEN_1338; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1597 = unuse_way == 2'h1 ? _GEN_697 : _GEN_1339; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1598 = unuse_way == 2'h1 ? _GEN_698 : _GEN_1340; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1599 = unuse_way == 2'h1 ? _GEN_699 : _GEN_1341; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1600 = unuse_way == 2'h1 ? _GEN_700 : _GEN_1342; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1601 = unuse_way == 2'h1 ? _GEN_701 : _GEN_1343; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1602 = unuse_way == 2'h1 ? _GEN_702 : _GEN_1344; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1603 = unuse_way == 2'h1 ? _GEN_703 : _GEN_1345; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1604 = unuse_way == 2'h1 ? _GEN_704 : _GEN_1346; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1605 = unuse_way == 2'h1 ? _GEN_705 : _GEN_1347; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1606 = unuse_way == 2'h1 ? _GEN_706 : _GEN_1348; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1607 = unuse_way == 2'h1 ? _GEN_707 : _GEN_1349; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1608 = unuse_way == 2'h1 ? _GEN_708 : _GEN_1350; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1609 = unuse_way == 2'h1 ? _GEN_709 : _GEN_1351; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1610 = unuse_way == 2'h1 ? _GEN_710 : _GEN_1352; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1611 = unuse_way == 2'h1 ? _GEN_711 : _GEN_1353; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1612 = unuse_way == 2'h1 ? _GEN_712 : _GEN_1354; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1613 = unuse_way == 2'h1 ? _GEN_713 : _GEN_1355; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1614 = unuse_way == 2'h1 ? _GEN_714 : _GEN_1356; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1615 = unuse_way == 2'h1 ? _GEN_715 : _GEN_1357; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1616 = unuse_way == 2'h1 ? _GEN_716 : _GEN_1358; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1617 = unuse_way == 2'h1 ? _GEN_717 : _GEN_1359; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1618 = unuse_way == 2'h1 ? _GEN_718 : _GEN_1360; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1619 = unuse_way == 2'h1 ? _GEN_719 : _GEN_1361; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1620 = unuse_way == 2'h1 ? _GEN_720 : _GEN_1362; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1621 = unuse_way == 2'h1 ? _GEN_721 : _GEN_1363; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1622 = unuse_way == 2'h1 ? _GEN_722 : _GEN_1364; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1623 = unuse_way == 2'h1 ? _GEN_723 : _GEN_1365; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1624 = unuse_way == 2'h1 ? _GEN_724 : _GEN_1366; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1625 = unuse_way == 2'h1 ? _GEN_725 : _GEN_1367; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1626 = unuse_way == 2'h1 ? _GEN_726 : _GEN_1368; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1627 = unuse_way == 2'h1 ? _GEN_727 : _GEN_1369; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1628 = unuse_way == 2'h1 ? _GEN_728 : _GEN_1370; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1629 = unuse_way == 2'h1 ? _GEN_729 : _GEN_1371; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1630 = unuse_way == 2'h1 ? _GEN_730 : _GEN_1372; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1631 = unuse_way == 2'h1 ? _GEN_731 : _GEN_1373; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1632 = unuse_way == 2'h1 ? _GEN_732 : _GEN_1374; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1633 = unuse_way == 2'h1 ? _GEN_733 : _GEN_1375; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1634 = unuse_way == 2'h1 ? _GEN_734 : _GEN_1376; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1635 = unuse_way == 2'h1 ? _GEN_735 : _GEN_1377; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1636 = unuse_way == 2'h1 ? _GEN_736 : _GEN_1378; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1637 = unuse_way == 2'h1 ? _GEN_737 : _GEN_1379; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1638 = unuse_way == 2'h1 ? _GEN_738 : _GEN_1380; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1639 = unuse_way == 2'h1 ? _GEN_739 : _GEN_1381; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1640 = unuse_way == 2'h1 ? _GEN_740 : _GEN_1382; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1641 = unuse_way == 2'h1 ? _GEN_741 : _GEN_1383; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1642 = unuse_way == 2'h1 ? _GEN_742 : _GEN_1384; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1643 = unuse_way == 2'h1 ? _GEN_743 : _GEN_1385; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1644 = unuse_way == 2'h1 ? _GEN_744 : _GEN_1386; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1645 = unuse_way == 2'h1 ? _GEN_745 : _GEN_1387; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1646 = unuse_way == 2'h1 ? _GEN_746 : _GEN_1388; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1647 = unuse_way == 2'h1 ? _GEN_747 : _GEN_1389; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1648 = unuse_way == 2'h1 ? _GEN_748 : _GEN_1390; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1649 = unuse_way == 2'h1 ? _GEN_749 : _GEN_1391; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1650 = unuse_way == 2'h1 ? _GEN_750 : _GEN_1392; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1651 = unuse_way == 2'h1 ? _GEN_751 : _GEN_1393; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1652 = unuse_way == 2'h1 ? _GEN_752 : _GEN_1394; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1653 = unuse_way == 2'h1 ? _GEN_753 : _GEN_1395; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1654 = unuse_way == 2'h1 ? _GEN_754 : _GEN_1396; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1655 = unuse_way == 2'h1 ? _GEN_755 : _GEN_1397; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1656 = unuse_way == 2'h1 ? _GEN_756 : _GEN_1398; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1657 = unuse_way == 2'h1 ? _GEN_757 : _GEN_1399; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1658 = unuse_way == 2'h1 ? _GEN_758 : _GEN_1400; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1659 = unuse_way == 2'h1 ? _GEN_759 : _GEN_1401; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1660 = unuse_way == 2'h1 ? _GEN_760 : _GEN_1402; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1661 = unuse_way == 2'h1 ? _GEN_761 : _GEN_1403; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1662 = unuse_way == 2'h1 ? _GEN_762 : _GEN_1404; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1663 = unuse_way == 2'h1 ? _GEN_763 : _GEN_1405; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1664 = unuse_way == 2'h1 ? _GEN_764 : _GEN_1406; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1665 = unuse_way == 2'h1 ? _GEN_765 : _GEN_1407; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1666 = unuse_way == 2'h1 ? _GEN_766 : _GEN_1408; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1667 = unuse_way == 2'h1 ? _GEN_767 : _GEN_1409; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1668 = unuse_way == 2'h1 ? _GEN_768 : _GEN_1410; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1669 = unuse_way == 2'h1 ? _GEN_769 : _GEN_1411; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1670 = unuse_way == 2'h1 ? _GEN_770 : _GEN_1412; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1671 = unuse_way == 2'h1 ? _GEN_771 : _GEN_1413; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1672 = unuse_way == 2'h1 ? _GEN_772 : _GEN_1414; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1673 = unuse_way == 2'h1 ? _GEN_773 : _GEN_1415; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1674 = unuse_way == 2'h1 ? _GEN_774 : _GEN_1416; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1675 = unuse_way == 2'h1 ? _GEN_775 : _GEN_1417; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1676 = unuse_way == 2'h1 ? _GEN_776 : _GEN_1418; // @[d_cache.scala 141:34]
  wire [31:0] _GEN_1677 = unuse_way == 2'h1 ? _GEN_777 : _GEN_1419; // @[d_cache.scala 141:34]
  wire  _GEN_1678 = unuse_way == 2'h1 ? _GEN_326 : _GEN_1484; // @[d_cache.scala 141:34]
  wire  _GEN_1679 = unuse_way == 2'h1 ? _GEN_327 : _GEN_1485; // @[d_cache.scala 141:34]
  wire  _GEN_1680 = unuse_way == 2'h1 ? _GEN_328 : _GEN_1486; // @[d_cache.scala 141:34]
  wire  _GEN_1681 = unuse_way == 2'h1 ? _GEN_329 : _GEN_1487; // @[d_cache.scala 141:34]
  wire  _GEN_1682 = unuse_way == 2'h1 ? _GEN_330 : _GEN_1488; // @[d_cache.scala 141:34]
  wire  _GEN_1683 = unuse_way == 2'h1 ? _GEN_331 : _GEN_1489; // @[d_cache.scala 141:34]
  wire  _GEN_1684 = unuse_way == 2'h1 ? _GEN_332 : _GEN_1490; // @[d_cache.scala 141:34]
  wire  _GEN_1685 = unuse_way == 2'h1 ? _GEN_333 : _GEN_1491; // @[d_cache.scala 141:34]
  wire  _GEN_1686 = unuse_way == 2'h1 ? _GEN_334 : _GEN_1492; // @[d_cache.scala 141:34]
  wire  _GEN_1687 = unuse_way == 2'h1 ? _GEN_335 : _GEN_1493; // @[d_cache.scala 141:34]
  wire  _GEN_1688 = unuse_way == 2'h1 ? _GEN_336 : _GEN_1494; // @[d_cache.scala 141:34]
  wire  _GEN_1689 = unuse_way == 2'h1 ? _GEN_337 : _GEN_1495; // @[d_cache.scala 141:34]
  wire  _GEN_1690 = unuse_way == 2'h1 ? _GEN_338 : _GEN_1496; // @[d_cache.scala 141:34]
  wire  _GEN_1691 = unuse_way == 2'h1 ? _GEN_339 : _GEN_1497; // @[d_cache.scala 141:34]
  wire  _GEN_1692 = unuse_way == 2'h1 ? _GEN_340 : _GEN_1498; // @[d_cache.scala 141:34]
  wire  _GEN_1693 = unuse_way == 2'h1 ? _GEN_341 : _GEN_1499; // @[d_cache.scala 141:34]
  wire  _GEN_1694 = unuse_way == 2'h1 ? _GEN_342 : _GEN_1500; // @[d_cache.scala 141:34]
  wire  _GEN_1695 = unuse_way == 2'h1 ? _GEN_343 : _GEN_1501; // @[d_cache.scala 141:34]
  wire  _GEN_1696 = unuse_way == 2'h1 ? _GEN_344 : _GEN_1502; // @[d_cache.scala 141:34]
  wire  _GEN_1697 = unuse_way == 2'h1 ? _GEN_345 : _GEN_1503; // @[d_cache.scala 141:34]
  wire  _GEN_1698 = unuse_way == 2'h1 ? _GEN_346 : _GEN_1504; // @[d_cache.scala 141:34]
  wire  _GEN_1699 = unuse_way == 2'h1 ? _GEN_347 : _GEN_1505; // @[d_cache.scala 141:34]
  wire  _GEN_1700 = unuse_way == 2'h1 ? _GEN_348 : _GEN_1506; // @[d_cache.scala 141:34]
  wire  _GEN_1701 = unuse_way == 2'h1 ? _GEN_349 : _GEN_1507; // @[d_cache.scala 141:34]
  wire  _GEN_1702 = unuse_way == 2'h1 ? _GEN_350 : _GEN_1508; // @[d_cache.scala 141:34]
  wire  _GEN_1703 = unuse_way == 2'h1 ? _GEN_351 : _GEN_1509; // @[d_cache.scala 141:34]
  wire  _GEN_1704 = unuse_way == 2'h1 ? _GEN_352 : _GEN_1510; // @[d_cache.scala 141:34]
  wire  _GEN_1705 = unuse_way == 2'h1 ? _GEN_353 : _GEN_1511; // @[d_cache.scala 141:34]
  wire  _GEN_1706 = unuse_way == 2'h1 ? _GEN_354 : _GEN_1512; // @[d_cache.scala 141:34]
  wire  _GEN_1707 = unuse_way == 2'h1 ? _GEN_355 : _GEN_1513; // @[d_cache.scala 141:34]
  wire  _GEN_1708 = unuse_way == 2'h1 ? _GEN_356 : _GEN_1514; // @[d_cache.scala 141:34]
  wire  _GEN_1709 = unuse_way == 2'h1 ? _GEN_357 : _GEN_1515; // @[d_cache.scala 141:34]
  wire  _GEN_1710 = unuse_way == 2'h1 ? _GEN_358 : _GEN_1516; // @[d_cache.scala 141:34]
  wire  _GEN_1711 = unuse_way == 2'h1 ? _GEN_359 : _GEN_1517; // @[d_cache.scala 141:34]
  wire  _GEN_1712 = unuse_way == 2'h1 ? _GEN_360 : _GEN_1518; // @[d_cache.scala 141:34]
  wire  _GEN_1713 = unuse_way == 2'h1 ? _GEN_361 : _GEN_1519; // @[d_cache.scala 141:34]
  wire  _GEN_1714 = unuse_way == 2'h1 ? _GEN_362 : _GEN_1520; // @[d_cache.scala 141:34]
  wire  _GEN_1715 = unuse_way == 2'h1 ? _GEN_363 : _GEN_1521; // @[d_cache.scala 141:34]
  wire  _GEN_1716 = unuse_way == 2'h1 ? _GEN_364 : _GEN_1522; // @[d_cache.scala 141:34]
  wire  _GEN_1717 = unuse_way == 2'h1 ? _GEN_365 : _GEN_1523; // @[d_cache.scala 141:34]
  wire  _GEN_1718 = unuse_way == 2'h1 ? _GEN_366 : _GEN_1524; // @[d_cache.scala 141:34]
  wire  _GEN_1719 = unuse_way == 2'h1 ? _GEN_367 : _GEN_1525; // @[d_cache.scala 141:34]
  wire  _GEN_1720 = unuse_way == 2'h1 ? _GEN_368 : _GEN_1526; // @[d_cache.scala 141:34]
  wire  _GEN_1721 = unuse_way == 2'h1 ? _GEN_369 : _GEN_1527; // @[d_cache.scala 141:34]
  wire  _GEN_1722 = unuse_way == 2'h1 ? _GEN_370 : _GEN_1528; // @[d_cache.scala 141:34]
  wire  _GEN_1723 = unuse_way == 2'h1 ? _GEN_371 : _GEN_1529; // @[d_cache.scala 141:34]
  wire  _GEN_1724 = unuse_way == 2'h1 ? _GEN_372 : _GEN_1530; // @[d_cache.scala 141:34]
  wire  _GEN_1725 = unuse_way == 2'h1 ? _GEN_373 : _GEN_1531; // @[d_cache.scala 141:34]
  wire  _GEN_1726 = unuse_way == 2'h1 ? _GEN_374 : _GEN_1532; // @[d_cache.scala 141:34]
  wire  _GEN_1727 = unuse_way == 2'h1 ? _GEN_375 : _GEN_1533; // @[d_cache.scala 141:34]
  wire  _GEN_1728 = unuse_way == 2'h1 ? _GEN_376 : _GEN_1534; // @[d_cache.scala 141:34]
  wire  _GEN_1729 = unuse_way == 2'h1 ? _GEN_377 : _GEN_1535; // @[d_cache.scala 141:34]
  wire  _GEN_1730 = unuse_way == 2'h1 ? _GEN_378 : _GEN_1536; // @[d_cache.scala 141:34]
  wire  _GEN_1731 = unuse_way == 2'h1 ? _GEN_379 : _GEN_1537; // @[d_cache.scala 141:34]
  wire  _GEN_1732 = unuse_way == 2'h1 ? _GEN_380 : _GEN_1538; // @[d_cache.scala 141:34]
  wire  _GEN_1733 = unuse_way == 2'h1 ? _GEN_381 : _GEN_1539; // @[d_cache.scala 141:34]
  wire  _GEN_1734 = unuse_way == 2'h1 ? _GEN_382 : _GEN_1540; // @[d_cache.scala 141:34]
  wire  _GEN_1735 = unuse_way == 2'h1 ? _GEN_383 : _GEN_1541; // @[d_cache.scala 141:34]
  wire  _GEN_1736 = unuse_way == 2'h1 ? _GEN_384 : _GEN_1542; // @[d_cache.scala 141:34]
  wire  _GEN_1737 = unuse_way == 2'h1 ? _GEN_385 : _GEN_1543; // @[d_cache.scala 141:34]
  wire  _GEN_1738 = unuse_way == 2'h1 ? _GEN_386 : _GEN_1544; // @[d_cache.scala 141:34]
  wire  _GEN_1739 = unuse_way == 2'h1 ? _GEN_387 : _GEN_1545; // @[d_cache.scala 141:34]
  wire  _GEN_1740 = unuse_way == 2'h1 ? _GEN_388 : _GEN_1546; // @[d_cache.scala 141:34]
  wire  _GEN_1741 = unuse_way == 2'h1 ? _GEN_389 : _GEN_1547; // @[d_cache.scala 141:34]
  wire [63:0] _GEN_1742 = unuse_way == 2'h1 ? write_back_data : _GEN_1290; // @[d_cache.scala 141:34 31:34]
  wire [40:0] _GEN_1743 = unuse_way == 2'h1 ? {{9'd0}, write_back_addr} : _GEN_1291; // @[d_cache.scala 141:34 32:34]
  wire  _GEN_1744 = unuse_way == 2'h1 ? dirty_0_0 : _GEN_1420; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1745 = unuse_way == 2'h1 ? dirty_0_1 : _GEN_1421; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1746 = unuse_way == 2'h1 ? dirty_0_2 : _GEN_1422; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1747 = unuse_way == 2'h1 ? dirty_0_3 : _GEN_1423; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1748 = unuse_way == 2'h1 ? dirty_0_4 : _GEN_1424; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1749 = unuse_way == 2'h1 ? dirty_0_5 : _GEN_1425; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1750 = unuse_way == 2'h1 ? dirty_0_6 : _GEN_1426; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1751 = unuse_way == 2'h1 ? dirty_0_7 : _GEN_1427; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1752 = unuse_way == 2'h1 ? dirty_0_8 : _GEN_1428; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1753 = unuse_way == 2'h1 ? dirty_0_9 : _GEN_1429; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1754 = unuse_way == 2'h1 ? dirty_0_10 : _GEN_1430; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1755 = unuse_way == 2'h1 ? dirty_0_11 : _GEN_1431; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1756 = unuse_way == 2'h1 ? dirty_0_12 : _GEN_1432; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1757 = unuse_way == 2'h1 ? dirty_0_13 : _GEN_1433; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1758 = unuse_way == 2'h1 ? dirty_0_14 : _GEN_1434; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1759 = unuse_way == 2'h1 ? dirty_0_15 : _GEN_1435; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1760 = unuse_way == 2'h1 ? dirty_0_16 : _GEN_1436; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1761 = unuse_way == 2'h1 ? dirty_0_17 : _GEN_1437; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1762 = unuse_way == 2'h1 ? dirty_0_18 : _GEN_1438; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1763 = unuse_way == 2'h1 ? dirty_0_19 : _GEN_1439; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1764 = unuse_way == 2'h1 ? dirty_0_20 : _GEN_1440; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1765 = unuse_way == 2'h1 ? dirty_0_21 : _GEN_1441; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1766 = unuse_way == 2'h1 ? dirty_0_22 : _GEN_1442; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1767 = unuse_way == 2'h1 ? dirty_0_23 : _GEN_1443; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1768 = unuse_way == 2'h1 ? dirty_0_24 : _GEN_1444; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1769 = unuse_way == 2'h1 ? dirty_0_25 : _GEN_1445; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1770 = unuse_way == 2'h1 ? dirty_0_26 : _GEN_1446; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1771 = unuse_way == 2'h1 ? dirty_0_27 : _GEN_1447; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1772 = unuse_way == 2'h1 ? dirty_0_28 : _GEN_1448; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1773 = unuse_way == 2'h1 ? dirty_0_29 : _GEN_1449; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1774 = unuse_way == 2'h1 ? dirty_0_30 : _GEN_1450; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1775 = unuse_way == 2'h1 ? dirty_0_31 : _GEN_1451; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1776 = unuse_way == 2'h1 ? dirty_0_32 : _GEN_1452; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1777 = unuse_way == 2'h1 ? dirty_0_33 : _GEN_1453; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1778 = unuse_way == 2'h1 ? dirty_0_34 : _GEN_1454; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1779 = unuse_way == 2'h1 ? dirty_0_35 : _GEN_1455; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1780 = unuse_way == 2'h1 ? dirty_0_36 : _GEN_1456; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1781 = unuse_way == 2'h1 ? dirty_0_37 : _GEN_1457; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1782 = unuse_way == 2'h1 ? dirty_0_38 : _GEN_1458; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1783 = unuse_way == 2'h1 ? dirty_0_39 : _GEN_1459; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1784 = unuse_way == 2'h1 ? dirty_0_40 : _GEN_1460; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1785 = unuse_way == 2'h1 ? dirty_0_41 : _GEN_1461; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1786 = unuse_way == 2'h1 ? dirty_0_42 : _GEN_1462; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1787 = unuse_way == 2'h1 ? dirty_0_43 : _GEN_1463; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1788 = unuse_way == 2'h1 ? dirty_0_44 : _GEN_1464; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1789 = unuse_way == 2'h1 ? dirty_0_45 : _GEN_1465; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1790 = unuse_way == 2'h1 ? dirty_0_46 : _GEN_1466; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1791 = unuse_way == 2'h1 ? dirty_0_47 : _GEN_1467; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1792 = unuse_way == 2'h1 ? dirty_0_48 : _GEN_1468; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1793 = unuse_way == 2'h1 ? dirty_0_49 : _GEN_1469; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1794 = unuse_way == 2'h1 ? dirty_0_50 : _GEN_1470; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1795 = unuse_way == 2'h1 ? dirty_0_51 : _GEN_1471; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1796 = unuse_way == 2'h1 ? dirty_0_52 : _GEN_1472; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1797 = unuse_way == 2'h1 ? dirty_0_53 : _GEN_1473; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1798 = unuse_way == 2'h1 ? dirty_0_54 : _GEN_1474; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1799 = unuse_way == 2'h1 ? dirty_0_55 : _GEN_1475; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1800 = unuse_way == 2'h1 ? dirty_0_56 : _GEN_1476; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1801 = unuse_way == 2'h1 ? dirty_0_57 : _GEN_1477; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1802 = unuse_way == 2'h1 ? dirty_0_58 : _GEN_1478; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1803 = unuse_way == 2'h1 ? dirty_0_59 : _GEN_1479; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1804 = unuse_way == 2'h1 ? dirty_0_60 : _GEN_1480; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1805 = unuse_way == 2'h1 ? dirty_0_61 : _GEN_1481; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1806 = unuse_way == 2'h1 ? dirty_0_62 : _GEN_1482; // @[d_cache.scala 141:34 26:26]
  wire  _GEN_1807 = unuse_way == 2'h1 ? dirty_0_63 : _GEN_1483; // @[d_cache.scala 141:34 26:26]
  wire [2:0] _GEN_1808 = io_from_axi_bvalid ? 3'h7 : state; // @[d_cache.scala 193:37 194:23 76:24]
  wire [2:0] _GEN_1809 = 3'h7 == state ? 3'h1 : state; // @[d_cache.scala 81:18 198:19 76:24]
  wire [2:0] _GEN_1810 = 3'h6 == state ? _GEN_1808 : _GEN_1809; // @[d_cache.scala 81:18]
  wire [2:0] _GEN_1811 = 3'h5 == state ? _GEN_1549 : _GEN_1810; // @[d_cache.scala 81:18]
  wire [63:0] _GEN_1812 = 3'h5 == state ? _GEN_1550 : ram_0_0; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1813 = 3'h5 == state ? _GEN_1551 : ram_0_1; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1814 = 3'h5 == state ? _GEN_1552 : ram_0_2; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1815 = 3'h5 == state ? _GEN_1553 : ram_0_3; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1816 = 3'h5 == state ? _GEN_1554 : ram_0_4; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1817 = 3'h5 == state ? _GEN_1555 : ram_0_5; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1818 = 3'h5 == state ? _GEN_1556 : ram_0_6; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1819 = 3'h5 == state ? _GEN_1557 : ram_0_7; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1820 = 3'h5 == state ? _GEN_1558 : ram_0_8; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1821 = 3'h5 == state ? _GEN_1559 : ram_0_9; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1822 = 3'h5 == state ? _GEN_1560 : ram_0_10; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1823 = 3'h5 == state ? _GEN_1561 : ram_0_11; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1824 = 3'h5 == state ? _GEN_1562 : ram_0_12; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1825 = 3'h5 == state ? _GEN_1563 : ram_0_13; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1826 = 3'h5 == state ? _GEN_1564 : ram_0_14; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1827 = 3'h5 == state ? _GEN_1565 : ram_0_15; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1828 = 3'h5 == state ? _GEN_1566 : ram_0_16; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1829 = 3'h5 == state ? _GEN_1567 : ram_0_17; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1830 = 3'h5 == state ? _GEN_1568 : ram_0_18; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1831 = 3'h5 == state ? _GEN_1569 : ram_0_19; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1832 = 3'h5 == state ? _GEN_1570 : ram_0_20; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1833 = 3'h5 == state ? _GEN_1571 : ram_0_21; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1834 = 3'h5 == state ? _GEN_1572 : ram_0_22; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1835 = 3'h5 == state ? _GEN_1573 : ram_0_23; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1836 = 3'h5 == state ? _GEN_1574 : ram_0_24; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1837 = 3'h5 == state ? _GEN_1575 : ram_0_25; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1838 = 3'h5 == state ? _GEN_1576 : ram_0_26; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1839 = 3'h5 == state ? _GEN_1577 : ram_0_27; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1840 = 3'h5 == state ? _GEN_1578 : ram_0_28; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1841 = 3'h5 == state ? _GEN_1579 : ram_0_29; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1842 = 3'h5 == state ? _GEN_1580 : ram_0_30; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1843 = 3'h5 == state ? _GEN_1581 : ram_0_31; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1844 = 3'h5 == state ? _GEN_1582 : ram_0_32; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1845 = 3'h5 == state ? _GEN_1583 : ram_0_33; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1846 = 3'h5 == state ? _GEN_1584 : ram_0_34; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1847 = 3'h5 == state ? _GEN_1585 : ram_0_35; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1848 = 3'h5 == state ? _GEN_1586 : ram_0_36; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1849 = 3'h5 == state ? _GEN_1587 : ram_0_37; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1850 = 3'h5 == state ? _GEN_1588 : ram_0_38; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1851 = 3'h5 == state ? _GEN_1589 : ram_0_39; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1852 = 3'h5 == state ? _GEN_1590 : ram_0_40; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1853 = 3'h5 == state ? _GEN_1591 : ram_0_41; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1854 = 3'h5 == state ? _GEN_1592 : ram_0_42; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1855 = 3'h5 == state ? _GEN_1593 : ram_0_43; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1856 = 3'h5 == state ? _GEN_1594 : ram_0_44; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1857 = 3'h5 == state ? _GEN_1595 : ram_0_45; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1858 = 3'h5 == state ? _GEN_1596 : ram_0_46; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1859 = 3'h5 == state ? _GEN_1597 : ram_0_47; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1860 = 3'h5 == state ? _GEN_1598 : ram_0_48; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1861 = 3'h5 == state ? _GEN_1599 : ram_0_49; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1862 = 3'h5 == state ? _GEN_1600 : ram_0_50; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1863 = 3'h5 == state ? _GEN_1601 : ram_0_51; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1864 = 3'h5 == state ? _GEN_1602 : ram_0_52; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1865 = 3'h5 == state ? _GEN_1603 : ram_0_53; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1866 = 3'h5 == state ? _GEN_1604 : ram_0_54; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1867 = 3'h5 == state ? _GEN_1605 : ram_0_55; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1868 = 3'h5 == state ? _GEN_1606 : ram_0_56; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1869 = 3'h5 == state ? _GEN_1607 : ram_0_57; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1870 = 3'h5 == state ? _GEN_1608 : ram_0_58; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1871 = 3'h5 == state ? _GEN_1609 : ram_0_59; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1872 = 3'h5 == state ? _GEN_1610 : ram_0_60; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1873 = 3'h5 == state ? _GEN_1611 : ram_0_61; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1874 = 3'h5 == state ? _GEN_1612 : ram_0_62; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_1875 = 3'h5 == state ? _GEN_1613 : ram_0_63; // @[d_cache.scala 81:18 18:24]
  wire [31:0] _GEN_1876 = 3'h5 == state ? _GEN_1614 : tag_0_0; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1877 = 3'h5 == state ? _GEN_1615 : tag_0_1; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1878 = 3'h5 == state ? _GEN_1616 : tag_0_2; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1879 = 3'h5 == state ? _GEN_1617 : tag_0_3; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1880 = 3'h5 == state ? _GEN_1618 : tag_0_4; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1881 = 3'h5 == state ? _GEN_1619 : tag_0_5; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1882 = 3'h5 == state ? _GEN_1620 : tag_0_6; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1883 = 3'h5 == state ? _GEN_1621 : tag_0_7; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1884 = 3'h5 == state ? _GEN_1622 : tag_0_8; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1885 = 3'h5 == state ? _GEN_1623 : tag_0_9; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1886 = 3'h5 == state ? _GEN_1624 : tag_0_10; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1887 = 3'h5 == state ? _GEN_1625 : tag_0_11; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1888 = 3'h5 == state ? _GEN_1626 : tag_0_12; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1889 = 3'h5 == state ? _GEN_1627 : tag_0_13; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1890 = 3'h5 == state ? _GEN_1628 : tag_0_14; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1891 = 3'h5 == state ? _GEN_1629 : tag_0_15; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1892 = 3'h5 == state ? _GEN_1630 : tag_0_16; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1893 = 3'h5 == state ? _GEN_1631 : tag_0_17; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1894 = 3'h5 == state ? _GEN_1632 : tag_0_18; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1895 = 3'h5 == state ? _GEN_1633 : tag_0_19; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1896 = 3'h5 == state ? _GEN_1634 : tag_0_20; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1897 = 3'h5 == state ? _GEN_1635 : tag_0_21; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1898 = 3'h5 == state ? _GEN_1636 : tag_0_22; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1899 = 3'h5 == state ? _GEN_1637 : tag_0_23; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1900 = 3'h5 == state ? _GEN_1638 : tag_0_24; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1901 = 3'h5 == state ? _GEN_1639 : tag_0_25; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1902 = 3'h5 == state ? _GEN_1640 : tag_0_26; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1903 = 3'h5 == state ? _GEN_1641 : tag_0_27; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1904 = 3'h5 == state ? _GEN_1642 : tag_0_28; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1905 = 3'h5 == state ? _GEN_1643 : tag_0_29; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1906 = 3'h5 == state ? _GEN_1644 : tag_0_30; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1907 = 3'h5 == state ? _GEN_1645 : tag_0_31; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1908 = 3'h5 == state ? _GEN_1646 : tag_0_32; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1909 = 3'h5 == state ? _GEN_1647 : tag_0_33; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1910 = 3'h5 == state ? _GEN_1648 : tag_0_34; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1911 = 3'h5 == state ? _GEN_1649 : tag_0_35; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1912 = 3'h5 == state ? _GEN_1650 : tag_0_36; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1913 = 3'h5 == state ? _GEN_1651 : tag_0_37; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1914 = 3'h5 == state ? _GEN_1652 : tag_0_38; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1915 = 3'h5 == state ? _GEN_1653 : tag_0_39; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1916 = 3'h5 == state ? _GEN_1654 : tag_0_40; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1917 = 3'h5 == state ? _GEN_1655 : tag_0_41; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1918 = 3'h5 == state ? _GEN_1656 : tag_0_42; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1919 = 3'h5 == state ? _GEN_1657 : tag_0_43; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1920 = 3'h5 == state ? _GEN_1658 : tag_0_44; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1921 = 3'h5 == state ? _GEN_1659 : tag_0_45; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1922 = 3'h5 == state ? _GEN_1660 : tag_0_46; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1923 = 3'h5 == state ? _GEN_1661 : tag_0_47; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1924 = 3'h5 == state ? _GEN_1662 : tag_0_48; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1925 = 3'h5 == state ? _GEN_1663 : tag_0_49; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1926 = 3'h5 == state ? _GEN_1664 : tag_0_50; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1927 = 3'h5 == state ? _GEN_1665 : tag_0_51; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1928 = 3'h5 == state ? _GEN_1666 : tag_0_52; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1929 = 3'h5 == state ? _GEN_1667 : tag_0_53; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1930 = 3'h5 == state ? _GEN_1668 : tag_0_54; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1931 = 3'h5 == state ? _GEN_1669 : tag_0_55; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1932 = 3'h5 == state ? _GEN_1670 : tag_0_56; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1933 = 3'h5 == state ? _GEN_1671 : tag_0_57; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1934 = 3'h5 == state ? _GEN_1672 : tag_0_58; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1935 = 3'h5 == state ? _GEN_1673 : tag_0_59; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1936 = 3'h5 == state ? _GEN_1674 : tag_0_60; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1937 = 3'h5 == state ? _GEN_1675 : tag_0_61; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1938 = 3'h5 == state ? _GEN_1676 : tag_0_62; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_1939 = 3'h5 == state ? _GEN_1677 : tag_0_63; // @[d_cache.scala 81:18 22:24]
  wire  _GEN_1940 = 3'h5 == state ? _GEN_1678 : valid_0_0; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1941 = 3'h5 == state ? _GEN_1679 : valid_0_1; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1942 = 3'h5 == state ? _GEN_1680 : valid_0_2; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1943 = 3'h5 == state ? _GEN_1681 : valid_0_3; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1944 = 3'h5 == state ? _GEN_1682 : valid_0_4; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1945 = 3'h5 == state ? _GEN_1683 : valid_0_5; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1946 = 3'h5 == state ? _GEN_1684 : valid_0_6; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1947 = 3'h5 == state ? _GEN_1685 : valid_0_7; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1948 = 3'h5 == state ? _GEN_1686 : valid_0_8; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1949 = 3'h5 == state ? _GEN_1687 : valid_0_9; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1950 = 3'h5 == state ? _GEN_1688 : valid_0_10; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1951 = 3'h5 == state ? _GEN_1689 : valid_0_11; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1952 = 3'h5 == state ? _GEN_1690 : valid_0_12; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1953 = 3'h5 == state ? _GEN_1691 : valid_0_13; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1954 = 3'h5 == state ? _GEN_1692 : valid_0_14; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1955 = 3'h5 == state ? _GEN_1693 : valid_0_15; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1956 = 3'h5 == state ? _GEN_1694 : valid_0_16; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1957 = 3'h5 == state ? _GEN_1695 : valid_0_17; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1958 = 3'h5 == state ? _GEN_1696 : valid_0_18; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1959 = 3'h5 == state ? _GEN_1697 : valid_0_19; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1960 = 3'h5 == state ? _GEN_1698 : valid_0_20; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1961 = 3'h5 == state ? _GEN_1699 : valid_0_21; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1962 = 3'h5 == state ? _GEN_1700 : valid_0_22; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1963 = 3'h5 == state ? _GEN_1701 : valid_0_23; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1964 = 3'h5 == state ? _GEN_1702 : valid_0_24; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1965 = 3'h5 == state ? _GEN_1703 : valid_0_25; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1966 = 3'h5 == state ? _GEN_1704 : valid_0_26; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1967 = 3'h5 == state ? _GEN_1705 : valid_0_27; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1968 = 3'h5 == state ? _GEN_1706 : valid_0_28; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1969 = 3'h5 == state ? _GEN_1707 : valid_0_29; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1970 = 3'h5 == state ? _GEN_1708 : valid_0_30; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1971 = 3'h5 == state ? _GEN_1709 : valid_0_31; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1972 = 3'h5 == state ? _GEN_1710 : valid_0_32; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1973 = 3'h5 == state ? _GEN_1711 : valid_0_33; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1974 = 3'h5 == state ? _GEN_1712 : valid_0_34; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1975 = 3'h5 == state ? _GEN_1713 : valid_0_35; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1976 = 3'h5 == state ? _GEN_1714 : valid_0_36; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1977 = 3'h5 == state ? _GEN_1715 : valid_0_37; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1978 = 3'h5 == state ? _GEN_1716 : valid_0_38; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1979 = 3'h5 == state ? _GEN_1717 : valid_0_39; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1980 = 3'h5 == state ? _GEN_1718 : valid_0_40; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1981 = 3'h5 == state ? _GEN_1719 : valid_0_41; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1982 = 3'h5 == state ? _GEN_1720 : valid_0_42; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1983 = 3'h5 == state ? _GEN_1721 : valid_0_43; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1984 = 3'h5 == state ? _GEN_1722 : valid_0_44; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1985 = 3'h5 == state ? _GEN_1723 : valid_0_45; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1986 = 3'h5 == state ? _GEN_1724 : valid_0_46; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1987 = 3'h5 == state ? _GEN_1725 : valid_0_47; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1988 = 3'h5 == state ? _GEN_1726 : valid_0_48; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1989 = 3'h5 == state ? _GEN_1727 : valid_0_49; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1990 = 3'h5 == state ? _GEN_1728 : valid_0_50; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1991 = 3'h5 == state ? _GEN_1729 : valid_0_51; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1992 = 3'h5 == state ? _GEN_1730 : valid_0_52; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1993 = 3'h5 == state ? _GEN_1731 : valid_0_53; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1994 = 3'h5 == state ? _GEN_1732 : valid_0_54; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1995 = 3'h5 == state ? _GEN_1733 : valid_0_55; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1996 = 3'h5 == state ? _GEN_1734 : valid_0_56; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1997 = 3'h5 == state ? _GEN_1735 : valid_0_57; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1998 = 3'h5 == state ? _GEN_1736 : valid_0_58; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_1999 = 3'h5 == state ? _GEN_1737 : valid_0_59; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2000 = 3'h5 == state ? _GEN_1738 : valid_0_60; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2001 = 3'h5 == state ? _GEN_1739 : valid_0_61; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2002 = 3'h5 == state ? _GEN_1740 : valid_0_62; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2003 = 3'h5 == state ? _GEN_1741 : valid_0_63; // @[d_cache.scala 81:18 24:26]
  wire [63:0] _GEN_2004 = 3'h5 == state ? _GEN_1742 : write_back_data; // @[d_cache.scala 81:18 31:34]
  wire [40:0] _GEN_2005 = 3'h5 == state ? _GEN_1743 : {{9'd0}, write_back_addr}; // @[d_cache.scala 81:18 32:34]
  wire  _GEN_2006 = 3'h5 == state ? _GEN_1744 : dirty_0_0; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2007 = 3'h5 == state ? _GEN_1745 : dirty_0_1; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2008 = 3'h5 == state ? _GEN_1746 : dirty_0_2; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2009 = 3'h5 == state ? _GEN_1747 : dirty_0_3; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2010 = 3'h5 == state ? _GEN_1748 : dirty_0_4; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2011 = 3'h5 == state ? _GEN_1749 : dirty_0_5; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2012 = 3'h5 == state ? _GEN_1750 : dirty_0_6; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2013 = 3'h5 == state ? _GEN_1751 : dirty_0_7; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2014 = 3'h5 == state ? _GEN_1752 : dirty_0_8; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2015 = 3'h5 == state ? _GEN_1753 : dirty_0_9; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2016 = 3'h5 == state ? _GEN_1754 : dirty_0_10; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2017 = 3'h5 == state ? _GEN_1755 : dirty_0_11; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2018 = 3'h5 == state ? _GEN_1756 : dirty_0_12; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2019 = 3'h5 == state ? _GEN_1757 : dirty_0_13; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2020 = 3'h5 == state ? _GEN_1758 : dirty_0_14; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2021 = 3'h5 == state ? _GEN_1759 : dirty_0_15; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2022 = 3'h5 == state ? _GEN_1760 : dirty_0_16; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2023 = 3'h5 == state ? _GEN_1761 : dirty_0_17; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2024 = 3'h5 == state ? _GEN_1762 : dirty_0_18; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2025 = 3'h5 == state ? _GEN_1763 : dirty_0_19; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2026 = 3'h5 == state ? _GEN_1764 : dirty_0_20; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2027 = 3'h5 == state ? _GEN_1765 : dirty_0_21; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2028 = 3'h5 == state ? _GEN_1766 : dirty_0_22; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2029 = 3'h5 == state ? _GEN_1767 : dirty_0_23; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2030 = 3'h5 == state ? _GEN_1768 : dirty_0_24; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2031 = 3'h5 == state ? _GEN_1769 : dirty_0_25; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2032 = 3'h5 == state ? _GEN_1770 : dirty_0_26; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2033 = 3'h5 == state ? _GEN_1771 : dirty_0_27; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2034 = 3'h5 == state ? _GEN_1772 : dirty_0_28; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2035 = 3'h5 == state ? _GEN_1773 : dirty_0_29; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2036 = 3'h5 == state ? _GEN_1774 : dirty_0_30; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2037 = 3'h5 == state ? _GEN_1775 : dirty_0_31; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2038 = 3'h5 == state ? _GEN_1776 : dirty_0_32; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2039 = 3'h5 == state ? _GEN_1777 : dirty_0_33; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2040 = 3'h5 == state ? _GEN_1778 : dirty_0_34; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2041 = 3'h5 == state ? _GEN_1779 : dirty_0_35; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2042 = 3'h5 == state ? _GEN_1780 : dirty_0_36; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2043 = 3'h5 == state ? _GEN_1781 : dirty_0_37; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2044 = 3'h5 == state ? _GEN_1782 : dirty_0_38; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2045 = 3'h5 == state ? _GEN_1783 : dirty_0_39; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2046 = 3'h5 == state ? _GEN_1784 : dirty_0_40; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2047 = 3'h5 == state ? _GEN_1785 : dirty_0_41; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2048 = 3'h5 == state ? _GEN_1786 : dirty_0_42; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2049 = 3'h5 == state ? _GEN_1787 : dirty_0_43; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2050 = 3'h5 == state ? _GEN_1788 : dirty_0_44; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2051 = 3'h5 == state ? _GEN_1789 : dirty_0_45; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2052 = 3'h5 == state ? _GEN_1790 : dirty_0_46; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2053 = 3'h5 == state ? _GEN_1791 : dirty_0_47; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2054 = 3'h5 == state ? _GEN_1792 : dirty_0_48; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2055 = 3'h5 == state ? _GEN_1793 : dirty_0_49; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2056 = 3'h5 == state ? _GEN_1794 : dirty_0_50; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2057 = 3'h5 == state ? _GEN_1795 : dirty_0_51; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2058 = 3'h5 == state ? _GEN_1796 : dirty_0_52; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2059 = 3'h5 == state ? _GEN_1797 : dirty_0_53; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2060 = 3'h5 == state ? _GEN_1798 : dirty_0_54; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2061 = 3'h5 == state ? _GEN_1799 : dirty_0_55; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2062 = 3'h5 == state ? _GEN_1800 : dirty_0_56; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2063 = 3'h5 == state ? _GEN_1801 : dirty_0_57; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2064 = 3'h5 == state ? _GEN_1802 : dirty_0_58; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2065 = 3'h5 == state ? _GEN_1803 : dirty_0_59; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2066 = 3'h5 == state ? _GEN_1804 : dirty_0_60; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2067 = 3'h5 == state ? _GEN_1805 : dirty_0_61; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2068 = 3'h5 == state ? _GEN_1806 : dirty_0_62; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2069 = 3'h5 == state ? _GEN_1807 : dirty_0_63; // @[d_cache.scala 81:18 26:26]
  wire [2:0] _GEN_2070 = 3'h4 == state ? _GEN_649 : _GEN_1811; // @[d_cache.scala 81:18]
  wire [63:0] _GEN_2071 = 3'h4 == state ? ram_0_0 : _GEN_1812; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2072 = 3'h4 == state ? ram_0_1 : _GEN_1813; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2073 = 3'h4 == state ? ram_0_2 : _GEN_1814; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2074 = 3'h4 == state ? ram_0_3 : _GEN_1815; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2075 = 3'h4 == state ? ram_0_4 : _GEN_1816; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2076 = 3'h4 == state ? ram_0_5 : _GEN_1817; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2077 = 3'h4 == state ? ram_0_6 : _GEN_1818; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2078 = 3'h4 == state ? ram_0_7 : _GEN_1819; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2079 = 3'h4 == state ? ram_0_8 : _GEN_1820; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2080 = 3'h4 == state ? ram_0_9 : _GEN_1821; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2081 = 3'h4 == state ? ram_0_10 : _GEN_1822; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2082 = 3'h4 == state ? ram_0_11 : _GEN_1823; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2083 = 3'h4 == state ? ram_0_12 : _GEN_1824; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2084 = 3'h4 == state ? ram_0_13 : _GEN_1825; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2085 = 3'h4 == state ? ram_0_14 : _GEN_1826; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2086 = 3'h4 == state ? ram_0_15 : _GEN_1827; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2087 = 3'h4 == state ? ram_0_16 : _GEN_1828; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2088 = 3'h4 == state ? ram_0_17 : _GEN_1829; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2089 = 3'h4 == state ? ram_0_18 : _GEN_1830; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2090 = 3'h4 == state ? ram_0_19 : _GEN_1831; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2091 = 3'h4 == state ? ram_0_20 : _GEN_1832; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2092 = 3'h4 == state ? ram_0_21 : _GEN_1833; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2093 = 3'h4 == state ? ram_0_22 : _GEN_1834; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2094 = 3'h4 == state ? ram_0_23 : _GEN_1835; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2095 = 3'h4 == state ? ram_0_24 : _GEN_1836; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2096 = 3'h4 == state ? ram_0_25 : _GEN_1837; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2097 = 3'h4 == state ? ram_0_26 : _GEN_1838; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2098 = 3'h4 == state ? ram_0_27 : _GEN_1839; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2099 = 3'h4 == state ? ram_0_28 : _GEN_1840; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2100 = 3'h4 == state ? ram_0_29 : _GEN_1841; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2101 = 3'h4 == state ? ram_0_30 : _GEN_1842; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2102 = 3'h4 == state ? ram_0_31 : _GEN_1843; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2103 = 3'h4 == state ? ram_0_32 : _GEN_1844; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2104 = 3'h4 == state ? ram_0_33 : _GEN_1845; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2105 = 3'h4 == state ? ram_0_34 : _GEN_1846; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2106 = 3'h4 == state ? ram_0_35 : _GEN_1847; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2107 = 3'h4 == state ? ram_0_36 : _GEN_1848; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2108 = 3'h4 == state ? ram_0_37 : _GEN_1849; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2109 = 3'h4 == state ? ram_0_38 : _GEN_1850; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2110 = 3'h4 == state ? ram_0_39 : _GEN_1851; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2111 = 3'h4 == state ? ram_0_40 : _GEN_1852; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2112 = 3'h4 == state ? ram_0_41 : _GEN_1853; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2113 = 3'h4 == state ? ram_0_42 : _GEN_1854; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2114 = 3'h4 == state ? ram_0_43 : _GEN_1855; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2115 = 3'h4 == state ? ram_0_44 : _GEN_1856; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2116 = 3'h4 == state ? ram_0_45 : _GEN_1857; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2117 = 3'h4 == state ? ram_0_46 : _GEN_1858; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2118 = 3'h4 == state ? ram_0_47 : _GEN_1859; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2119 = 3'h4 == state ? ram_0_48 : _GEN_1860; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2120 = 3'h4 == state ? ram_0_49 : _GEN_1861; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2121 = 3'h4 == state ? ram_0_50 : _GEN_1862; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2122 = 3'h4 == state ? ram_0_51 : _GEN_1863; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2123 = 3'h4 == state ? ram_0_52 : _GEN_1864; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2124 = 3'h4 == state ? ram_0_53 : _GEN_1865; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2125 = 3'h4 == state ? ram_0_54 : _GEN_1866; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2126 = 3'h4 == state ? ram_0_55 : _GEN_1867; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2127 = 3'h4 == state ? ram_0_56 : _GEN_1868; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2128 = 3'h4 == state ? ram_0_57 : _GEN_1869; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2129 = 3'h4 == state ? ram_0_58 : _GEN_1870; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2130 = 3'h4 == state ? ram_0_59 : _GEN_1871; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2131 = 3'h4 == state ? ram_0_60 : _GEN_1872; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2132 = 3'h4 == state ? ram_0_61 : _GEN_1873; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2133 = 3'h4 == state ? ram_0_62 : _GEN_1874; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2134 = 3'h4 == state ? ram_0_63 : _GEN_1875; // @[d_cache.scala 81:18 18:24]
  wire [31:0] _GEN_2135 = 3'h4 == state ? tag_0_0 : _GEN_1876; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2136 = 3'h4 == state ? tag_0_1 : _GEN_1877; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2137 = 3'h4 == state ? tag_0_2 : _GEN_1878; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2138 = 3'h4 == state ? tag_0_3 : _GEN_1879; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2139 = 3'h4 == state ? tag_0_4 : _GEN_1880; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2140 = 3'h4 == state ? tag_0_5 : _GEN_1881; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2141 = 3'h4 == state ? tag_0_6 : _GEN_1882; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2142 = 3'h4 == state ? tag_0_7 : _GEN_1883; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2143 = 3'h4 == state ? tag_0_8 : _GEN_1884; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2144 = 3'h4 == state ? tag_0_9 : _GEN_1885; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2145 = 3'h4 == state ? tag_0_10 : _GEN_1886; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2146 = 3'h4 == state ? tag_0_11 : _GEN_1887; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2147 = 3'h4 == state ? tag_0_12 : _GEN_1888; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2148 = 3'h4 == state ? tag_0_13 : _GEN_1889; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2149 = 3'h4 == state ? tag_0_14 : _GEN_1890; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2150 = 3'h4 == state ? tag_0_15 : _GEN_1891; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2151 = 3'h4 == state ? tag_0_16 : _GEN_1892; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2152 = 3'h4 == state ? tag_0_17 : _GEN_1893; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2153 = 3'h4 == state ? tag_0_18 : _GEN_1894; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2154 = 3'h4 == state ? tag_0_19 : _GEN_1895; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2155 = 3'h4 == state ? tag_0_20 : _GEN_1896; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2156 = 3'h4 == state ? tag_0_21 : _GEN_1897; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2157 = 3'h4 == state ? tag_0_22 : _GEN_1898; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2158 = 3'h4 == state ? tag_0_23 : _GEN_1899; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2159 = 3'h4 == state ? tag_0_24 : _GEN_1900; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2160 = 3'h4 == state ? tag_0_25 : _GEN_1901; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2161 = 3'h4 == state ? tag_0_26 : _GEN_1902; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2162 = 3'h4 == state ? tag_0_27 : _GEN_1903; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2163 = 3'h4 == state ? tag_0_28 : _GEN_1904; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2164 = 3'h4 == state ? tag_0_29 : _GEN_1905; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2165 = 3'h4 == state ? tag_0_30 : _GEN_1906; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2166 = 3'h4 == state ? tag_0_31 : _GEN_1907; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2167 = 3'h4 == state ? tag_0_32 : _GEN_1908; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2168 = 3'h4 == state ? tag_0_33 : _GEN_1909; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2169 = 3'h4 == state ? tag_0_34 : _GEN_1910; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2170 = 3'h4 == state ? tag_0_35 : _GEN_1911; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2171 = 3'h4 == state ? tag_0_36 : _GEN_1912; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2172 = 3'h4 == state ? tag_0_37 : _GEN_1913; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2173 = 3'h4 == state ? tag_0_38 : _GEN_1914; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2174 = 3'h4 == state ? tag_0_39 : _GEN_1915; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2175 = 3'h4 == state ? tag_0_40 : _GEN_1916; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2176 = 3'h4 == state ? tag_0_41 : _GEN_1917; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2177 = 3'h4 == state ? tag_0_42 : _GEN_1918; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2178 = 3'h4 == state ? tag_0_43 : _GEN_1919; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2179 = 3'h4 == state ? tag_0_44 : _GEN_1920; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2180 = 3'h4 == state ? tag_0_45 : _GEN_1921; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2181 = 3'h4 == state ? tag_0_46 : _GEN_1922; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2182 = 3'h4 == state ? tag_0_47 : _GEN_1923; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2183 = 3'h4 == state ? tag_0_48 : _GEN_1924; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2184 = 3'h4 == state ? tag_0_49 : _GEN_1925; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2185 = 3'h4 == state ? tag_0_50 : _GEN_1926; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2186 = 3'h4 == state ? tag_0_51 : _GEN_1927; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2187 = 3'h4 == state ? tag_0_52 : _GEN_1928; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2188 = 3'h4 == state ? tag_0_53 : _GEN_1929; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2189 = 3'h4 == state ? tag_0_54 : _GEN_1930; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2190 = 3'h4 == state ? tag_0_55 : _GEN_1931; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2191 = 3'h4 == state ? tag_0_56 : _GEN_1932; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2192 = 3'h4 == state ? tag_0_57 : _GEN_1933; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2193 = 3'h4 == state ? tag_0_58 : _GEN_1934; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2194 = 3'h4 == state ? tag_0_59 : _GEN_1935; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2195 = 3'h4 == state ? tag_0_60 : _GEN_1936; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2196 = 3'h4 == state ? tag_0_61 : _GEN_1937; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2197 = 3'h4 == state ? tag_0_62 : _GEN_1938; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2198 = 3'h4 == state ? tag_0_63 : _GEN_1939; // @[d_cache.scala 81:18 22:24]
  wire  _GEN_2199 = 3'h4 == state ? valid_0_0 : _GEN_1940; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2200 = 3'h4 == state ? valid_0_1 : _GEN_1941; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2201 = 3'h4 == state ? valid_0_2 : _GEN_1942; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2202 = 3'h4 == state ? valid_0_3 : _GEN_1943; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2203 = 3'h4 == state ? valid_0_4 : _GEN_1944; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2204 = 3'h4 == state ? valid_0_5 : _GEN_1945; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2205 = 3'h4 == state ? valid_0_6 : _GEN_1946; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2206 = 3'h4 == state ? valid_0_7 : _GEN_1947; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2207 = 3'h4 == state ? valid_0_8 : _GEN_1948; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2208 = 3'h4 == state ? valid_0_9 : _GEN_1949; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2209 = 3'h4 == state ? valid_0_10 : _GEN_1950; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2210 = 3'h4 == state ? valid_0_11 : _GEN_1951; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2211 = 3'h4 == state ? valid_0_12 : _GEN_1952; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2212 = 3'h4 == state ? valid_0_13 : _GEN_1953; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2213 = 3'h4 == state ? valid_0_14 : _GEN_1954; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2214 = 3'h4 == state ? valid_0_15 : _GEN_1955; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2215 = 3'h4 == state ? valid_0_16 : _GEN_1956; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2216 = 3'h4 == state ? valid_0_17 : _GEN_1957; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2217 = 3'h4 == state ? valid_0_18 : _GEN_1958; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2218 = 3'h4 == state ? valid_0_19 : _GEN_1959; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2219 = 3'h4 == state ? valid_0_20 : _GEN_1960; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2220 = 3'h4 == state ? valid_0_21 : _GEN_1961; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2221 = 3'h4 == state ? valid_0_22 : _GEN_1962; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2222 = 3'h4 == state ? valid_0_23 : _GEN_1963; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2223 = 3'h4 == state ? valid_0_24 : _GEN_1964; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2224 = 3'h4 == state ? valid_0_25 : _GEN_1965; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2225 = 3'h4 == state ? valid_0_26 : _GEN_1966; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2226 = 3'h4 == state ? valid_0_27 : _GEN_1967; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2227 = 3'h4 == state ? valid_0_28 : _GEN_1968; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2228 = 3'h4 == state ? valid_0_29 : _GEN_1969; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2229 = 3'h4 == state ? valid_0_30 : _GEN_1970; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2230 = 3'h4 == state ? valid_0_31 : _GEN_1971; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2231 = 3'h4 == state ? valid_0_32 : _GEN_1972; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2232 = 3'h4 == state ? valid_0_33 : _GEN_1973; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2233 = 3'h4 == state ? valid_0_34 : _GEN_1974; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2234 = 3'h4 == state ? valid_0_35 : _GEN_1975; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2235 = 3'h4 == state ? valid_0_36 : _GEN_1976; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2236 = 3'h4 == state ? valid_0_37 : _GEN_1977; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2237 = 3'h4 == state ? valid_0_38 : _GEN_1978; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2238 = 3'h4 == state ? valid_0_39 : _GEN_1979; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2239 = 3'h4 == state ? valid_0_40 : _GEN_1980; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2240 = 3'h4 == state ? valid_0_41 : _GEN_1981; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2241 = 3'h4 == state ? valid_0_42 : _GEN_1982; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2242 = 3'h4 == state ? valid_0_43 : _GEN_1983; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2243 = 3'h4 == state ? valid_0_44 : _GEN_1984; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2244 = 3'h4 == state ? valid_0_45 : _GEN_1985; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2245 = 3'h4 == state ? valid_0_46 : _GEN_1986; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2246 = 3'h4 == state ? valid_0_47 : _GEN_1987; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2247 = 3'h4 == state ? valid_0_48 : _GEN_1988; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2248 = 3'h4 == state ? valid_0_49 : _GEN_1989; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2249 = 3'h4 == state ? valid_0_50 : _GEN_1990; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2250 = 3'h4 == state ? valid_0_51 : _GEN_1991; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2251 = 3'h4 == state ? valid_0_52 : _GEN_1992; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2252 = 3'h4 == state ? valid_0_53 : _GEN_1993; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2253 = 3'h4 == state ? valid_0_54 : _GEN_1994; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2254 = 3'h4 == state ? valid_0_55 : _GEN_1995; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2255 = 3'h4 == state ? valid_0_56 : _GEN_1996; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2256 = 3'h4 == state ? valid_0_57 : _GEN_1997; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2257 = 3'h4 == state ? valid_0_58 : _GEN_1998; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2258 = 3'h4 == state ? valid_0_59 : _GEN_1999; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2259 = 3'h4 == state ? valid_0_60 : _GEN_2000; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2260 = 3'h4 == state ? valid_0_61 : _GEN_2001; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2261 = 3'h4 == state ? valid_0_62 : _GEN_2002; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2262 = 3'h4 == state ? valid_0_63 : _GEN_2003; // @[d_cache.scala 81:18 24:26]
  wire [63:0] _GEN_2263 = 3'h4 == state ? write_back_data : _GEN_2004; // @[d_cache.scala 81:18 31:34]
  wire [40:0] _GEN_2264 = 3'h4 == state ? {{9'd0}, write_back_addr} : _GEN_2005; // @[d_cache.scala 81:18 32:34]
  wire  _GEN_2265 = 3'h4 == state ? dirty_0_0 : _GEN_2006; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2266 = 3'h4 == state ? dirty_0_1 : _GEN_2007; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2267 = 3'h4 == state ? dirty_0_2 : _GEN_2008; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2268 = 3'h4 == state ? dirty_0_3 : _GEN_2009; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2269 = 3'h4 == state ? dirty_0_4 : _GEN_2010; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2270 = 3'h4 == state ? dirty_0_5 : _GEN_2011; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2271 = 3'h4 == state ? dirty_0_6 : _GEN_2012; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2272 = 3'h4 == state ? dirty_0_7 : _GEN_2013; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2273 = 3'h4 == state ? dirty_0_8 : _GEN_2014; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2274 = 3'h4 == state ? dirty_0_9 : _GEN_2015; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2275 = 3'h4 == state ? dirty_0_10 : _GEN_2016; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2276 = 3'h4 == state ? dirty_0_11 : _GEN_2017; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2277 = 3'h4 == state ? dirty_0_12 : _GEN_2018; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2278 = 3'h4 == state ? dirty_0_13 : _GEN_2019; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2279 = 3'h4 == state ? dirty_0_14 : _GEN_2020; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2280 = 3'h4 == state ? dirty_0_15 : _GEN_2021; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2281 = 3'h4 == state ? dirty_0_16 : _GEN_2022; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2282 = 3'h4 == state ? dirty_0_17 : _GEN_2023; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2283 = 3'h4 == state ? dirty_0_18 : _GEN_2024; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2284 = 3'h4 == state ? dirty_0_19 : _GEN_2025; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2285 = 3'h4 == state ? dirty_0_20 : _GEN_2026; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2286 = 3'h4 == state ? dirty_0_21 : _GEN_2027; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2287 = 3'h4 == state ? dirty_0_22 : _GEN_2028; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2288 = 3'h4 == state ? dirty_0_23 : _GEN_2029; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2289 = 3'h4 == state ? dirty_0_24 : _GEN_2030; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2290 = 3'h4 == state ? dirty_0_25 : _GEN_2031; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2291 = 3'h4 == state ? dirty_0_26 : _GEN_2032; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2292 = 3'h4 == state ? dirty_0_27 : _GEN_2033; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2293 = 3'h4 == state ? dirty_0_28 : _GEN_2034; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2294 = 3'h4 == state ? dirty_0_29 : _GEN_2035; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2295 = 3'h4 == state ? dirty_0_30 : _GEN_2036; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2296 = 3'h4 == state ? dirty_0_31 : _GEN_2037; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2297 = 3'h4 == state ? dirty_0_32 : _GEN_2038; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2298 = 3'h4 == state ? dirty_0_33 : _GEN_2039; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2299 = 3'h4 == state ? dirty_0_34 : _GEN_2040; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2300 = 3'h4 == state ? dirty_0_35 : _GEN_2041; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2301 = 3'h4 == state ? dirty_0_36 : _GEN_2042; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2302 = 3'h4 == state ? dirty_0_37 : _GEN_2043; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2303 = 3'h4 == state ? dirty_0_38 : _GEN_2044; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2304 = 3'h4 == state ? dirty_0_39 : _GEN_2045; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2305 = 3'h4 == state ? dirty_0_40 : _GEN_2046; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2306 = 3'h4 == state ? dirty_0_41 : _GEN_2047; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2307 = 3'h4 == state ? dirty_0_42 : _GEN_2048; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2308 = 3'h4 == state ? dirty_0_43 : _GEN_2049; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2309 = 3'h4 == state ? dirty_0_44 : _GEN_2050; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2310 = 3'h4 == state ? dirty_0_45 : _GEN_2051; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2311 = 3'h4 == state ? dirty_0_46 : _GEN_2052; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2312 = 3'h4 == state ? dirty_0_47 : _GEN_2053; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2313 = 3'h4 == state ? dirty_0_48 : _GEN_2054; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2314 = 3'h4 == state ? dirty_0_49 : _GEN_2055; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2315 = 3'h4 == state ? dirty_0_50 : _GEN_2056; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2316 = 3'h4 == state ? dirty_0_51 : _GEN_2057; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2317 = 3'h4 == state ? dirty_0_52 : _GEN_2058; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2318 = 3'h4 == state ? dirty_0_53 : _GEN_2059; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2319 = 3'h4 == state ? dirty_0_54 : _GEN_2060; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2320 = 3'h4 == state ? dirty_0_55 : _GEN_2061; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2321 = 3'h4 == state ? dirty_0_56 : _GEN_2062; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2322 = 3'h4 == state ? dirty_0_57 : _GEN_2063; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2323 = 3'h4 == state ? dirty_0_58 : _GEN_2064; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2324 = 3'h4 == state ? dirty_0_59 : _GEN_2065; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2325 = 3'h4 == state ? dirty_0_60 : _GEN_2066; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2326 = 3'h4 == state ? dirty_0_61 : _GEN_2067; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2327 = 3'h4 == state ? dirty_0_62 : _GEN_2068; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2328 = 3'h4 == state ? dirty_0_63 : _GEN_2069; // @[d_cache.scala 81:18 26:26]
  wire [2:0] _GEN_2329 = 3'h3 == state ? _GEN_647 : _GEN_2070; // @[d_cache.scala 81:18]
  wire [63:0] _GEN_2330 = 3'h3 == state ? _GEN_648 : receive_data; // @[d_cache.scala 81:18 36:31]
  wire [63:0] _GEN_2331 = 3'h3 == state ? ram_0_0 : _GEN_2071; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2332 = 3'h3 == state ? ram_0_1 : _GEN_2072; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2333 = 3'h3 == state ? ram_0_2 : _GEN_2073; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2334 = 3'h3 == state ? ram_0_3 : _GEN_2074; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2335 = 3'h3 == state ? ram_0_4 : _GEN_2075; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2336 = 3'h3 == state ? ram_0_5 : _GEN_2076; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2337 = 3'h3 == state ? ram_0_6 : _GEN_2077; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2338 = 3'h3 == state ? ram_0_7 : _GEN_2078; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2339 = 3'h3 == state ? ram_0_8 : _GEN_2079; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2340 = 3'h3 == state ? ram_0_9 : _GEN_2080; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2341 = 3'h3 == state ? ram_0_10 : _GEN_2081; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2342 = 3'h3 == state ? ram_0_11 : _GEN_2082; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2343 = 3'h3 == state ? ram_0_12 : _GEN_2083; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2344 = 3'h3 == state ? ram_0_13 : _GEN_2084; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2345 = 3'h3 == state ? ram_0_14 : _GEN_2085; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2346 = 3'h3 == state ? ram_0_15 : _GEN_2086; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2347 = 3'h3 == state ? ram_0_16 : _GEN_2087; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2348 = 3'h3 == state ? ram_0_17 : _GEN_2088; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2349 = 3'h3 == state ? ram_0_18 : _GEN_2089; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2350 = 3'h3 == state ? ram_0_19 : _GEN_2090; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2351 = 3'h3 == state ? ram_0_20 : _GEN_2091; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2352 = 3'h3 == state ? ram_0_21 : _GEN_2092; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2353 = 3'h3 == state ? ram_0_22 : _GEN_2093; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2354 = 3'h3 == state ? ram_0_23 : _GEN_2094; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2355 = 3'h3 == state ? ram_0_24 : _GEN_2095; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2356 = 3'h3 == state ? ram_0_25 : _GEN_2096; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2357 = 3'h3 == state ? ram_0_26 : _GEN_2097; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2358 = 3'h3 == state ? ram_0_27 : _GEN_2098; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2359 = 3'h3 == state ? ram_0_28 : _GEN_2099; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2360 = 3'h3 == state ? ram_0_29 : _GEN_2100; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2361 = 3'h3 == state ? ram_0_30 : _GEN_2101; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2362 = 3'h3 == state ? ram_0_31 : _GEN_2102; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2363 = 3'h3 == state ? ram_0_32 : _GEN_2103; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2364 = 3'h3 == state ? ram_0_33 : _GEN_2104; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2365 = 3'h3 == state ? ram_0_34 : _GEN_2105; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2366 = 3'h3 == state ? ram_0_35 : _GEN_2106; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2367 = 3'h3 == state ? ram_0_36 : _GEN_2107; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2368 = 3'h3 == state ? ram_0_37 : _GEN_2108; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2369 = 3'h3 == state ? ram_0_38 : _GEN_2109; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2370 = 3'h3 == state ? ram_0_39 : _GEN_2110; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2371 = 3'h3 == state ? ram_0_40 : _GEN_2111; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2372 = 3'h3 == state ? ram_0_41 : _GEN_2112; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2373 = 3'h3 == state ? ram_0_42 : _GEN_2113; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2374 = 3'h3 == state ? ram_0_43 : _GEN_2114; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2375 = 3'h3 == state ? ram_0_44 : _GEN_2115; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2376 = 3'h3 == state ? ram_0_45 : _GEN_2116; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2377 = 3'h3 == state ? ram_0_46 : _GEN_2117; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2378 = 3'h3 == state ? ram_0_47 : _GEN_2118; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2379 = 3'h3 == state ? ram_0_48 : _GEN_2119; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2380 = 3'h3 == state ? ram_0_49 : _GEN_2120; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2381 = 3'h3 == state ? ram_0_50 : _GEN_2121; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2382 = 3'h3 == state ? ram_0_51 : _GEN_2122; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2383 = 3'h3 == state ? ram_0_52 : _GEN_2123; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2384 = 3'h3 == state ? ram_0_53 : _GEN_2124; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2385 = 3'h3 == state ? ram_0_54 : _GEN_2125; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2386 = 3'h3 == state ? ram_0_55 : _GEN_2126; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2387 = 3'h3 == state ? ram_0_56 : _GEN_2127; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2388 = 3'h3 == state ? ram_0_57 : _GEN_2128; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2389 = 3'h3 == state ? ram_0_58 : _GEN_2129; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2390 = 3'h3 == state ? ram_0_59 : _GEN_2130; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2391 = 3'h3 == state ? ram_0_60 : _GEN_2131; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2392 = 3'h3 == state ? ram_0_61 : _GEN_2132; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2393 = 3'h3 == state ? ram_0_62 : _GEN_2133; // @[d_cache.scala 81:18 18:24]
  wire [63:0] _GEN_2394 = 3'h3 == state ? ram_0_63 : _GEN_2134; // @[d_cache.scala 81:18 18:24]
  wire [31:0] _GEN_2395 = 3'h3 == state ? tag_0_0 : _GEN_2135; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2396 = 3'h3 == state ? tag_0_1 : _GEN_2136; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2397 = 3'h3 == state ? tag_0_2 : _GEN_2137; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2398 = 3'h3 == state ? tag_0_3 : _GEN_2138; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2399 = 3'h3 == state ? tag_0_4 : _GEN_2139; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2400 = 3'h3 == state ? tag_0_5 : _GEN_2140; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2401 = 3'h3 == state ? tag_0_6 : _GEN_2141; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2402 = 3'h3 == state ? tag_0_7 : _GEN_2142; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2403 = 3'h3 == state ? tag_0_8 : _GEN_2143; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2404 = 3'h3 == state ? tag_0_9 : _GEN_2144; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2405 = 3'h3 == state ? tag_0_10 : _GEN_2145; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2406 = 3'h3 == state ? tag_0_11 : _GEN_2146; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2407 = 3'h3 == state ? tag_0_12 : _GEN_2147; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2408 = 3'h3 == state ? tag_0_13 : _GEN_2148; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2409 = 3'h3 == state ? tag_0_14 : _GEN_2149; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2410 = 3'h3 == state ? tag_0_15 : _GEN_2150; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2411 = 3'h3 == state ? tag_0_16 : _GEN_2151; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2412 = 3'h3 == state ? tag_0_17 : _GEN_2152; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2413 = 3'h3 == state ? tag_0_18 : _GEN_2153; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2414 = 3'h3 == state ? tag_0_19 : _GEN_2154; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2415 = 3'h3 == state ? tag_0_20 : _GEN_2155; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2416 = 3'h3 == state ? tag_0_21 : _GEN_2156; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2417 = 3'h3 == state ? tag_0_22 : _GEN_2157; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2418 = 3'h3 == state ? tag_0_23 : _GEN_2158; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2419 = 3'h3 == state ? tag_0_24 : _GEN_2159; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2420 = 3'h3 == state ? tag_0_25 : _GEN_2160; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2421 = 3'h3 == state ? tag_0_26 : _GEN_2161; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2422 = 3'h3 == state ? tag_0_27 : _GEN_2162; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2423 = 3'h3 == state ? tag_0_28 : _GEN_2163; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2424 = 3'h3 == state ? tag_0_29 : _GEN_2164; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2425 = 3'h3 == state ? tag_0_30 : _GEN_2165; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2426 = 3'h3 == state ? tag_0_31 : _GEN_2166; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2427 = 3'h3 == state ? tag_0_32 : _GEN_2167; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2428 = 3'h3 == state ? tag_0_33 : _GEN_2168; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2429 = 3'h3 == state ? tag_0_34 : _GEN_2169; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2430 = 3'h3 == state ? tag_0_35 : _GEN_2170; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2431 = 3'h3 == state ? tag_0_36 : _GEN_2171; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2432 = 3'h3 == state ? tag_0_37 : _GEN_2172; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2433 = 3'h3 == state ? tag_0_38 : _GEN_2173; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2434 = 3'h3 == state ? tag_0_39 : _GEN_2174; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2435 = 3'h3 == state ? tag_0_40 : _GEN_2175; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2436 = 3'h3 == state ? tag_0_41 : _GEN_2176; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2437 = 3'h3 == state ? tag_0_42 : _GEN_2177; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2438 = 3'h3 == state ? tag_0_43 : _GEN_2178; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2439 = 3'h3 == state ? tag_0_44 : _GEN_2179; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2440 = 3'h3 == state ? tag_0_45 : _GEN_2180; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2441 = 3'h3 == state ? tag_0_46 : _GEN_2181; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2442 = 3'h3 == state ? tag_0_47 : _GEN_2182; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2443 = 3'h3 == state ? tag_0_48 : _GEN_2183; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2444 = 3'h3 == state ? tag_0_49 : _GEN_2184; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2445 = 3'h3 == state ? tag_0_50 : _GEN_2185; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2446 = 3'h3 == state ? tag_0_51 : _GEN_2186; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2447 = 3'h3 == state ? tag_0_52 : _GEN_2187; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2448 = 3'h3 == state ? tag_0_53 : _GEN_2188; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2449 = 3'h3 == state ? tag_0_54 : _GEN_2189; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2450 = 3'h3 == state ? tag_0_55 : _GEN_2190; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2451 = 3'h3 == state ? tag_0_56 : _GEN_2191; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2452 = 3'h3 == state ? tag_0_57 : _GEN_2192; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2453 = 3'h3 == state ? tag_0_58 : _GEN_2193; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2454 = 3'h3 == state ? tag_0_59 : _GEN_2194; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2455 = 3'h3 == state ? tag_0_60 : _GEN_2195; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2456 = 3'h3 == state ? tag_0_61 : _GEN_2196; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2457 = 3'h3 == state ? tag_0_62 : _GEN_2197; // @[d_cache.scala 81:18 22:24]
  wire [31:0] _GEN_2458 = 3'h3 == state ? tag_0_63 : _GEN_2198; // @[d_cache.scala 81:18 22:24]
  wire  _GEN_2459 = 3'h3 == state ? valid_0_0 : _GEN_2199; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2460 = 3'h3 == state ? valid_0_1 : _GEN_2200; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2461 = 3'h3 == state ? valid_0_2 : _GEN_2201; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2462 = 3'h3 == state ? valid_0_3 : _GEN_2202; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2463 = 3'h3 == state ? valid_0_4 : _GEN_2203; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2464 = 3'h3 == state ? valid_0_5 : _GEN_2204; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2465 = 3'h3 == state ? valid_0_6 : _GEN_2205; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2466 = 3'h3 == state ? valid_0_7 : _GEN_2206; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2467 = 3'h3 == state ? valid_0_8 : _GEN_2207; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2468 = 3'h3 == state ? valid_0_9 : _GEN_2208; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2469 = 3'h3 == state ? valid_0_10 : _GEN_2209; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2470 = 3'h3 == state ? valid_0_11 : _GEN_2210; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2471 = 3'h3 == state ? valid_0_12 : _GEN_2211; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2472 = 3'h3 == state ? valid_0_13 : _GEN_2212; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2473 = 3'h3 == state ? valid_0_14 : _GEN_2213; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2474 = 3'h3 == state ? valid_0_15 : _GEN_2214; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2475 = 3'h3 == state ? valid_0_16 : _GEN_2215; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2476 = 3'h3 == state ? valid_0_17 : _GEN_2216; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2477 = 3'h3 == state ? valid_0_18 : _GEN_2217; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2478 = 3'h3 == state ? valid_0_19 : _GEN_2218; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2479 = 3'h3 == state ? valid_0_20 : _GEN_2219; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2480 = 3'h3 == state ? valid_0_21 : _GEN_2220; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2481 = 3'h3 == state ? valid_0_22 : _GEN_2221; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2482 = 3'h3 == state ? valid_0_23 : _GEN_2222; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2483 = 3'h3 == state ? valid_0_24 : _GEN_2223; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2484 = 3'h3 == state ? valid_0_25 : _GEN_2224; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2485 = 3'h3 == state ? valid_0_26 : _GEN_2225; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2486 = 3'h3 == state ? valid_0_27 : _GEN_2226; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2487 = 3'h3 == state ? valid_0_28 : _GEN_2227; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2488 = 3'h3 == state ? valid_0_29 : _GEN_2228; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2489 = 3'h3 == state ? valid_0_30 : _GEN_2229; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2490 = 3'h3 == state ? valid_0_31 : _GEN_2230; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2491 = 3'h3 == state ? valid_0_32 : _GEN_2231; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2492 = 3'h3 == state ? valid_0_33 : _GEN_2232; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2493 = 3'h3 == state ? valid_0_34 : _GEN_2233; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2494 = 3'h3 == state ? valid_0_35 : _GEN_2234; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2495 = 3'h3 == state ? valid_0_36 : _GEN_2235; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2496 = 3'h3 == state ? valid_0_37 : _GEN_2236; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2497 = 3'h3 == state ? valid_0_38 : _GEN_2237; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2498 = 3'h3 == state ? valid_0_39 : _GEN_2238; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2499 = 3'h3 == state ? valid_0_40 : _GEN_2239; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2500 = 3'h3 == state ? valid_0_41 : _GEN_2240; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2501 = 3'h3 == state ? valid_0_42 : _GEN_2241; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2502 = 3'h3 == state ? valid_0_43 : _GEN_2242; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2503 = 3'h3 == state ? valid_0_44 : _GEN_2243; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2504 = 3'h3 == state ? valid_0_45 : _GEN_2244; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2505 = 3'h3 == state ? valid_0_46 : _GEN_2245; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2506 = 3'h3 == state ? valid_0_47 : _GEN_2246; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2507 = 3'h3 == state ? valid_0_48 : _GEN_2247; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2508 = 3'h3 == state ? valid_0_49 : _GEN_2248; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2509 = 3'h3 == state ? valid_0_50 : _GEN_2249; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2510 = 3'h3 == state ? valid_0_51 : _GEN_2250; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2511 = 3'h3 == state ? valid_0_52 : _GEN_2251; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2512 = 3'h3 == state ? valid_0_53 : _GEN_2252; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2513 = 3'h3 == state ? valid_0_54 : _GEN_2253; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2514 = 3'h3 == state ? valid_0_55 : _GEN_2254; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2515 = 3'h3 == state ? valid_0_56 : _GEN_2255; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2516 = 3'h3 == state ? valid_0_57 : _GEN_2256; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2517 = 3'h3 == state ? valid_0_58 : _GEN_2257; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2518 = 3'h3 == state ? valid_0_59 : _GEN_2258; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2519 = 3'h3 == state ? valid_0_60 : _GEN_2259; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2520 = 3'h3 == state ? valid_0_61 : _GEN_2260; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2521 = 3'h3 == state ? valid_0_62 : _GEN_2261; // @[d_cache.scala 81:18 24:26]
  wire  _GEN_2522 = 3'h3 == state ? valid_0_63 : _GEN_2262; // @[d_cache.scala 81:18 24:26]
  wire [63:0] _GEN_2523 = 3'h3 == state ? write_back_data : _GEN_2263; // @[d_cache.scala 81:18 31:34]
  wire [40:0] _GEN_2524 = 3'h3 == state ? {{9'd0}, write_back_addr} : _GEN_2264; // @[d_cache.scala 81:18 32:34]
  wire  _GEN_2525 = 3'h3 == state ? dirty_0_0 : _GEN_2265; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2526 = 3'h3 == state ? dirty_0_1 : _GEN_2266; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2527 = 3'h3 == state ? dirty_0_2 : _GEN_2267; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2528 = 3'h3 == state ? dirty_0_3 : _GEN_2268; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2529 = 3'h3 == state ? dirty_0_4 : _GEN_2269; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2530 = 3'h3 == state ? dirty_0_5 : _GEN_2270; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2531 = 3'h3 == state ? dirty_0_6 : _GEN_2271; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2532 = 3'h3 == state ? dirty_0_7 : _GEN_2272; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2533 = 3'h3 == state ? dirty_0_8 : _GEN_2273; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2534 = 3'h3 == state ? dirty_0_9 : _GEN_2274; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2535 = 3'h3 == state ? dirty_0_10 : _GEN_2275; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2536 = 3'h3 == state ? dirty_0_11 : _GEN_2276; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2537 = 3'h3 == state ? dirty_0_12 : _GEN_2277; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2538 = 3'h3 == state ? dirty_0_13 : _GEN_2278; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2539 = 3'h3 == state ? dirty_0_14 : _GEN_2279; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2540 = 3'h3 == state ? dirty_0_15 : _GEN_2280; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2541 = 3'h3 == state ? dirty_0_16 : _GEN_2281; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2542 = 3'h3 == state ? dirty_0_17 : _GEN_2282; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2543 = 3'h3 == state ? dirty_0_18 : _GEN_2283; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2544 = 3'h3 == state ? dirty_0_19 : _GEN_2284; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2545 = 3'h3 == state ? dirty_0_20 : _GEN_2285; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2546 = 3'h3 == state ? dirty_0_21 : _GEN_2286; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2547 = 3'h3 == state ? dirty_0_22 : _GEN_2287; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2548 = 3'h3 == state ? dirty_0_23 : _GEN_2288; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2549 = 3'h3 == state ? dirty_0_24 : _GEN_2289; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2550 = 3'h3 == state ? dirty_0_25 : _GEN_2290; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2551 = 3'h3 == state ? dirty_0_26 : _GEN_2291; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2552 = 3'h3 == state ? dirty_0_27 : _GEN_2292; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2553 = 3'h3 == state ? dirty_0_28 : _GEN_2293; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2554 = 3'h3 == state ? dirty_0_29 : _GEN_2294; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2555 = 3'h3 == state ? dirty_0_30 : _GEN_2295; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2556 = 3'h3 == state ? dirty_0_31 : _GEN_2296; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2557 = 3'h3 == state ? dirty_0_32 : _GEN_2297; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2558 = 3'h3 == state ? dirty_0_33 : _GEN_2298; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2559 = 3'h3 == state ? dirty_0_34 : _GEN_2299; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2560 = 3'h3 == state ? dirty_0_35 : _GEN_2300; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2561 = 3'h3 == state ? dirty_0_36 : _GEN_2301; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2562 = 3'h3 == state ? dirty_0_37 : _GEN_2302; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2563 = 3'h3 == state ? dirty_0_38 : _GEN_2303; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2564 = 3'h3 == state ? dirty_0_39 : _GEN_2304; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2565 = 3'h3 == state ? dirty_0_40 : _GEN_2305; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2566 = 3'h3 == state ? dirty_0_41 : _GEN_2306; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2567 = 3'h3 == state ? dirty_0_42 : _GEN_2307; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2568 = 3'h3 == state ? dirty_0_43 : _GEN_2308; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2569 = 3'h3 == state ? dirty_0_44 : _GEN_2309; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2570 = 3'h3 == state ? dirty_0_45 : _GEN_2310; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2571 = 3'h3 == state ? dirty_0_46 : _GEN_2311; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2572 = 3'h3 == state ? dirty_0_47 : _GEN_2312; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2573 = 3'h3 == state ? dirty_0_48 : _GEN_2313; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2574 = 3'h3 == state ? dirty_0_49 : _GEN_2314; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2575 = 3'h3 == state ? dirty_0_50 : _GEN_2315; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2576 = 3'h3 == state ? dirty_0_51 : _GEN_2316; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2577 = 3'h3 == state ? dirty_0_52 : _GEN_2317; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2578 = 3'h3 == state ? dirty_0_53 : _GEN_2318; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2579 = 3'h3 == state ? dirty_0_54 : _GEN_2319; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2580 = 3'h3 == state ? dirty_0_55 : _GEN_2320; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2581 = 3'h3 == state ? dirty_0_56 : _GEN_2321; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2582 = 3'h3 == state ? dirty_0_57 : _GEN_2322; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2583 = 3'h3 == state ? dirty_0_58 : _GEN_2323; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2584 = 3'h3 == state ? dirty_0_59 : _GEN_2324; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2585 = 3'h3 == state ? dirty_0_60 : _GEN_2325; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2586 = 3'h3 == state ? dirty_0_61 : _GEN_2326; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2587 = 3'h3 == state ? dirty_0_62 : _GEN_2327; // @[d_cache.scala 81:18 26:26]
  wire  _GEN_2588 = 3'h3 == state ? dirty_0_63 : _GEN_2328; // @[d_cache.scala 81:18 26:26]
  wire [40:0] _GEN_2848 = 3'h2 == state ? {{9'd0}, write_back_addr} : _GEN_2524; // @[d_cache.scala 81:18 32:34]
  wire [40:0] _GEN_3108 = 3'h1 == state ? {{9'd0}, write_back_addr} : _GEN_2848; // @[d_cache.scala 81:18 32:34]
  wire [40:0] _GEN_3368 = 3'h0 == state ? {{9'd0}, write_back_addr} : _GEN_3108; // @[d_cache.scala 81:18 32:34]
  wire [63:0] _io_to_lsu_rdata_T = _GEN_261 >> shift_bit; // @[d_cache.scala 228:49]
  wire [63:0] _GEN_3369 = way0_hit ? _io_to_lsu_rdata_T : 64'h0; // @[d_cache.scala 227:23 228:33 242:33]
  wire  _GEN_3373 = way0_hit ? 1'h0 : 1'h1; // @[d_cache.scala 259:23 261:35 275:35]
  wire  _T_25 = state == 3'h3; // @[d_cache.scala 281:21]
  wire [63:0] _GEN_3783 = {{32'd0}, io_from_lsu_araddr}; // @[d_cache.scala 289:48]
  wire [63:0] _io_to_axi_araddr_T = _GEN_3783 & 64'hfffffffffffffff8; // @[d_cache.scala 289:48]
  wire  _T_28 = state == 3'h6; // @[d_cache.scala 330:21]
  wire [31:0] _GEN_3376 = state == 3'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 330:35 338:26 354:26]
  wire  _GEN_3377 = state == 3'h6 ? 1'h0 : io_from_lsu_rready; // @[d_cache.scala 330:35 339:26 355:26]
  wire [31:0] _GEN_3378 = state == 3'h6 ? write_back_addr : 32'h0; // @[d_cache.scala 330:35 340:26 356:26]
  wire [63:0] _GEN_3379 = state == 3'h6 ? write_back_data : 64'h0; // @[d_cache.scala 330:35 342:25 358:25]
  wire [7:0] _GEN_3380 = state == 3'h6 ? 8'hff : 8'h0; // @[d_cache.scala 330:35 343:25 359:25]
  wire  _GEN_3382 = state == 3'h5 | _T_28; // @[d_cache.scala 314:31 316:27]
  wire [31:0] _GEN_3383 = state == 3'h5 ? io_from_lsu_araddr : _GEN_3376; // @[d_cache.scala 314:31 322:26]
  wire  _GEN_3384 = state == 3'h5 ? io_from_lsu_rready : _GEN_3377; // @[d_cache.scala 314:31 323:26]
  wire [31:0] _GEN_3385 = state == 3'h5 ? 32'h0 : _GEN_3378; // @[d_cache.scala 314:31 324:26]
  wire  _GEN_3386 = state == 3'h5 ? 1'h0 : _T_28; // @[d_cache.scala 314:31 325:27]
  wire [63:0] _GEN_3387 = state == 3'h5 ? 64'h0 : _GEN_3379; // @[d_cache.scala 314:31 326:25]
  wire [7:0] _GEN_3388 = state == 3'h5 ? 8'h0 : _GEN_3380; // @[d_cache.scala 314:31 327:25]
  wire  _GEN_3390 = state == 3'h4 | _GEN_3382; // @[d_cache.scala 297:31 299:27]
  wire  _GEN_3391 = state == 3'h4 & io_from_axi_wready; // @[d_cache.scala 297:31 301:26]
  wire  _GEN_3392 = state == 3'h4 & io_from_axi_bvalid; // @[d_cache.scala 297:31 302:26]
  wire  _GEN_3393 = state == 3'h4 & io_from_axi_awready; // @[d_cache.scala 297:31 303:27]
  wire [31:0] _GEN_3394 = state == 3'h4 ? 32'h0 : _GEN_3383; // @[d_cache.scala 297:31 305:26]
  wire  _GEN_3395 = state == 3'h4 ? io_from_lsu_rready : _GEN_3384; // @[d_cache.scala 297:31 306:26]
  wire [31:0] _GEN_3396 = state == 3'h4 ? io_from_lsu_awaddr : _GEN_3385; // @[d_cache.scala 297:31 307:26]
  wire  _GEN_3397 = state == 3'h4 ? io_from_lsu_awvalid : _GEN_3386; // @[d_cache.scala 297:31 308:27]
  wire [63:0] _GEN_3398 = state == 3'h4 ? {{32'd0}, io_from_lsu_wdata} : _GEN_3387; // @[d_cache.scala 297:31 309:25]
  wire [7:0] _GEN_3399 = state == 3'h4 ? io_from_lsu_wstrb : _GEN_3388; // @[d_cache.scala 297:31 310:25]
  wire  _GEN_3400 = state == 3'h4 ? io_from_lsu_wvalid : _GEN_3386; // @[d_cache.scala 297:31 311:26]
  wire  _GEN_3401 = state == 3'h4 ? io_from_lsu_bready : _GEN_3386; // @[d_cache.scala 297:31 312:26]
  wire  _GEN_3403 = state == 3'h3 | _GEN_3390; // @[d_cache.scala 281:31 283:27]
  wire  _GEN_3404 = state == 3'h3 ? 1'h0 : _GEN_3391; // @[d_cache.scala 281:31 285:26]
  wire  _GEN_3405 = state == 3'h3 ? 1'h0 : _GEN_3392; // @[d_cache.scala 281:31 286:26]
  wire  _GEN_3406 = state == 3'h3 ? 1'h0 : _GEN_3393; // @[d_cache.scala 281:31 287:27]
  wire [63:0] _GEN_3408 = state == 3'h3 ? _io_to_axi_araddr_T : {{32'd0}, _GEN_3394}; // @[d_cache.scala 281:31 289:26]
  wire  _GEN_3409 = state == 3'h3 ? io_from_lsu_rready : _GEN_3395; // @[d_cache.scala 281:31 290:26]
  wire [31:0] _GEN_3410 = state == 3'h3 ? 32'h0 : _GEN_3396; // @[d_cache.scala 281:31 291:26]
  wire  _GEN_3411 = state == 3'h3 ? 1'h0 : _GEN_3397; // @[d_cache.scala 281:31 292:27]
  wire [63:0] _GEN_3412 = state == 3'h3 ? 64'h0 : _GEN_3398; // @[d_cache.scala 281:31 293:25]
  wire [7:0] _GEN_3413 = state == 3'h3 ? 8'h0 : _GEN_3399; // @[d_cache.scala 281:31 294:25]
  wire  _GEN_3414 = state == 3'h3 ? 1'h0 : _GEN_3400; // @[d_cache.scala 281:31 295:26]
  wire  _GEN_3415 = state == 3'h3 ? 1'h0 : _GEN_3401; // @[d_cache.scala 281:31 296:26]
  wire  _GEN_3416 = state == 3'h2 ? 1'h0 : _T_25; // @[d_cache.scala 249:33 250:27]
  wire [63:0] _GEN_3417 = state == 3'h2 ? {{32'd0}, io_from_lsu_araddr} : _GEN_3408; // @[d_cache.scala 249:33 251:26]
  wire  _GEN_3418 = state == 3'h2 ? 1'h0 : _GEN_3409; // @[d_cache.scala 249:33 252:26]
  wire [31:0] _GEN_3419 = state == 3'h2 ? 32'h0 : _GEN_3410; // @[d_cache.scala 249:33 253:26]
  wire  _GEN_3420 = state == 3'h2 ? 1'h0 : _GEN_3411; // @[d_cache.scala 249:33 254:27]
  wire [63:0] _GEN_3421 = state == 3'h2 ? 64'h0 : _GEN_3412; // @[d_cache.scala 249:33 255:25]
  wire [7:0] _GEN_3422 = state == 3'h2 ? 8'h0 : _GEN_3413; // @[d_cache.scala 249:33 256:25]
  wire  _GEN_3423 = state == 3'h2 ? 1'h0 : _GEN_3414; // @[d_cache.scala 249:33 257:26]
  wire  _GEN_3424 = state == 3'h2 ? 1'h0 : _GEN_3415; // @[d_cache.scala 249:33 258:26]
  wire  _GEN_3426 = state == 3'h2 ? _GEN_3373 : _GEN_3403; // @[d_cache.scala 249:33]
  wire  _GEN_3427 = state == 3'h2 ? way0_hit : _GEN_3404; // @[d_cache.scala 249:33]
  wire  _GEN_3428 = state == 3'h2 ? way0_hit : _GEN_3406; // @[d_cache.scala 249:33]
  wire  _GEN_3429 = state == 3'h2 ? way0_hit : _GEN_3405; // @[d_cache.scala 249:33]
  wire  _GEN_3430 = state == 3'h1 ? 1'h0 : _GEN_3416; // @[d_cache.scala 217:33 218:27]
  wire [63:0] _GEN_3431 = state == 3'h1 ? {{32'd0}, io_from_lsu_araddr} : _GEN_3417; // @[d_cache.scala 217:33 219:26]
  wire  _GEN_3432 = state == 3'h1 ? io_from_lsu_rready : _GEN_3418; // @[d_cache.scala 217:33 220:26]
  wire [31:0] _GEN_3433 = state == 3'h1 ? 32'h0 : _GEN_3419; // @[d_cache.scala 217:33 221:26]
  wire  _GEN_3434 = state == 3'h1 ? 1'h0 : _GEN_3420; // @[d_cache.scala 217:33 222:27]
  wire [63:0] _GEN_3435 = state == 3'h1 ? 64'h0 : _GEN_3421; // @[d_cache.scala 217:33 223:25]
  wire [7:0] _GEN_3436 = state == 3'h1 ? 8'h0 : _GEN_3422; // @[d_cache.scala 217:33 224:25]
  wire  _GEN_3437 = state == 3'h1 ? 1'h0 : _GEN_3423; // @[d_cache.scala 217:33 225:26]
  wire  _GEN_3438 = state == 3'h1 ? io_from_lsu_bready : _GEN_3424; // @[d_cache.scala 217:33 226:26]
  wire [63:0] _GEN_3439 = state == 3'h1 ? _GEN_3369 : 64'h0; // @[d_cache.scala 217:33]
  wire  _GEN_3440 = state == 3'h1 | _GEN_3426; // @[d_cache.scala 217:33]
  wire  _GEN_3441 = state == 3'h1 & way0_hit; // @[d_cache.scala 217:33]
  wire  _GEN_3442 = state == 3'h1 ? 1'h0 : _GEN_3427; // @[d_cache.scala 217:33]
  wire  _GEN_3443 = state == 3'h1 ? 1'h0 : _GEN_3428; // @[d_cache.scala 217:33]
  wire  _GEN_3444 = state == 3'h1 ? 1'h0 : _GEN_3429; // @[d_cache.scala 217:33]
  wire [63:0] _GEN_3452 = state == 3'h0 ? {{32'd0}, io_from_lsu_araddr} : _GEN_3431; // @[d_cache.scala 201:23 209:26]
  wire [63:0] _GEN_3456 = state == 3'h0 ? 64'h0 : _GEN_3435; // @[d_cache.scala 201:23 213:25]
  wire [40:0] _GEN_3784 = reset ? 41'h0 : _GEN_3368; // @[d_cache.scala 32:{34,34}]
  assign io_to_lsu_arready = state == 3'h0 ? io_from_axi_arready : _GEN_3440; // @[d_cache.scala 201:23 203:27]
  assign io_to_lsu_rdata = state == 3'h0 ? 64'h0 : _GEN_3439; // @[d_cache.scala 201:23 202:25]
  assign io_to_lsu_rvalid = state == 3'h0 ? 1'h0 : _GEN_3441; // @[d_cache.scala 201:23 204:26]
  assign io_to_lsu_awready = state == 3'h0 ? io_from_axi_awready : _GEN_3443; // @[d_cache.scala 201:23 207:27]
  assign io_to_lsu_wready = state == 3'h0 ? 1'h0 : _GEN_3442; // @[d_cache.scala 201:23 205:26]
  assign io_to_lsu_bvalid = state == 3'h0 ? 1'h0 : _GEN_3444; // @[d_cache.scala 201:23 206:26]
  assign io_to_axi_araddr = _GEN_3452[31:0];
  assign io_to_axi_arvalid = state == 3'h0 ? 1'h0 : _GEN_3430; // @[d_cache.scala 201:23 208:27]
  assign io_to_axi_rready = state == 3'h0 ? io_from_lsu_rready : _GEN_3432; // @[d_cache.scala 201:23 210:26]
  assign io_to_axi_awaddr = state == 3'h0 ? 32'h0 : _GEN_3433; // @[d_cache.scala 201:23 211:26]
  assign io_to_axi_awvalid = state == 3'h0 ? 1'h0 : _GEN_3434; // @[d_cache.scala 201:23 212:27]
  assign io_to_axi_wdata = _GEN_3456[31:0];
  assign io_to_axi_wstrb = state == 3'h0 ? 8'h0 : _GEN_3436; // @[d_cache.scala 201:23 214:25]
  assign io_to_axi_wvalid = state == 3'h0 ? 1'h0 : _GEN_3437; // @[d_cache.scala 201:23 215:26]
  assign io_to_axi_bready = state == 3'h0 ? io_from_lsu_bready : _GEN_3438; // @[d_cache.scala 201:23 216:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_0 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_0 <= _GEN_455;
        end else begin
          ram_0_0 <= _GEN_2331;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_1 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_1 <= _GEN_456;
        end else begin
          ram_0_1 <= _GEN_2332;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_2 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_2 <= _GEN_457;
        end else begin
          ram_0_2 <= _GEN_2333;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_3 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_3 <= _GEN_458;
        end else begin
          ram_0_3 <= _GEN_2334;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_4 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_4 <= _GEN_459;
        end else begin
          ram_0_4 <= _GEN_2335;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_5 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_5 <= _GEN_460;
        end else begin
          ram_0_5 <= _GEN_2336;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_6 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_6 <= _GEN_461;
        end else begin
          ram_0_6 <= _GEN_2337;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_7 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_7 <= _GEN_462;
        end else begin
          ram_0_7 <= _GEN_2338;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_8 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_8 <= _GEN_463;
        end else begin
          ram_0_8 <= _GEN_2339;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_9 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_9 <= _GEN_464;
        end else begin
          ram_0_9 <= _GEN_2340;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_10 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_10 <= _GEN_465;
        end else begin
          ram_0_10 <= _GEN_2341;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_11 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_11 <= _GEN_466;
        end else begin
          ram_0_11 <= _GEN_2342;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_12 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_12 <= _GEN_467;
        end else begin
          ram_0_12 <= _GEN_2343;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_13 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_13 <= _GEN_468;
        end else begin
          ram_0_13 <= _GEN_2344;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_14 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_14 <= _GEN_469;
        end else begin
          ram_0_14 <= _GEN_2345;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_15 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_15 <= _GEN_470;
        end else begin
          ram_0_15 <= _GEN_2346;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_16 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_16 <= _GEN_471;
        end else begin
          ram_0_16 <= _GEN_2347;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_17 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_17 <= _GEN_472;
        end else begin
          ram_0_17 <= _GEN_2348;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_18 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_18 <= _GEN_473;
        end else begin
          ram_0_18 <= _GEN_2349;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_19 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_19 <= _GEN_474;
        end else begin
          ram_0_19 <= _GEN_2350;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_20 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_20 <= _GEN_475;
        end else begin
          ram_0_20 <= _GEN_2351;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_21 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_21 <= _GEN_476;
        end else begin
          ram_0_21 <= _GEN_2352;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_22 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_22 <= _GEN_477;
        end else begin
          ram_0_22 <= _GEN_2353;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_23 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_23 <= _GEN_478;
        end else begin
          ram_0_23 <= _GEN_2354;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_24 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_24 <= _GEN_479;
        end else begin
          ram_0_24 <= _GEN_2355;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_25 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_25 <= _GEN_480;
        end else begin
          ram_0_25 <= _GEN_2356;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_26 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_26 <= _GEN_481;
        end else begin
          ram_0_26 <= _GEN_2357;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_27 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_27 <= _GEN_482;
        end else begin
          ram_0_27 <= _GEN_2358;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_28 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_28 <= _GEN_483;
        end else begin
          ram_0_28 <= _GEN_2359;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_29 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_29 <= _GEN_484;
        end else begin
          ram_0_29 <= _GEN_2360;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_30 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_30 <= _GEN_485;
        end else begin
          ram_0_30 <= _GEN_2361;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_31 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_31 <= _GEN_486;
        end else begin
          ram_0_31 <= _GEN_2362;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_32 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_32 <= _GEN_487;
        end else begin
          ram_0_32 <= _GEN_2363;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_33 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_33 <= _GEN_488;
        end else begin
          ram_0_33 <= _GEN_2364;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_34 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_34 <= _GEN_489;
        end else begin
          ram_0_34 <= _GEN_2365;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_35 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_35 <= _GEN_490;
        end else begin
          ram_0_35 <= _GEN_2366;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_36 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_36 <= _GEN_491;
        end else begin
          ram_0_36 <= _GEN_2367;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_37 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_37 <= _GEN_492;
        end else begin
          ram_0_37 <= _GEN_2368;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_38 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_38 <= _GEN_493;
        end else begin
          ram_0_38 <= _GEN_2369;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_39 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_39 <= _GEN_494;
        end else begin
          ram_0_39 <= _GEN_2370;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_40 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_40 <= _GEN_495;
        end else begin
          ram_0_40 <= _GEN_2371;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_41 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_41 <= _GEN_496;
        end else begin
          ram_0_41 <= _GEN_2372;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_42 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_42 <= _GEN_497;
        end else begin
          ram_0_42 <= _GEN_2373;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_43 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_43 <= _GEN_498;
        end else begin
          ram_0_43 <= _GEN_2374;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_44 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_44 <= _GEN_499;
        end else begin
          ram_0_44 <= _GEN_2375;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_45 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_45 <= _GEN_500;
        end else begin
          ram_0_45 <= _GEN_2376;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_46 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_46 <= _GEN_501;
        end else begin
          ram_0_46 <= _GEN_2377;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_47 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_47 <= _GEN_502;
        end else begin
          ram_0_47 <= _GEN_2378;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_48 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_48 <= _GEN_503;
        end else begin
          ram_0_48 <= _GEN_2379;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_49 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_49 <= _GEN_504;
        end else begin
          ram_0_49 <= _GEN_2380;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_50 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_50 <= _GEN_505;
        end else begin
          ram_0_50 <= _GEN_2381;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_51 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_51 <= _GEN_506;
        end else begin
          ram_0_51 <= _GEN_2382;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_52 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_52 <= _GEN_507;
        end else begin
          ram_0_52 <= _GEN_2383;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_53 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_53 <= _GEN_508;
        end else begin
          ram_0_53 <= _GEN_2384;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_54 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_54 <= _GEN_509;
        end else begin
          ram_0_54 <= _GEN_2385;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_55 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_55 <= _GEN_510;
        end else begin
          ram_0_55 <= _GEN_2386;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_56 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_56 <= _GEN_511;
        end else begin
          ram_0_56 <= _GEN_2387;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_57 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_57 <= _GEN_512;
        end else begin
          ram_0_57 <= _GEN_2388;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_58 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_58 <= _GEN_513;
        end else begin
          ram_0_58 <= _GEN_2389;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_59 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_59 <= _GEN_514;
        end else begin
          ram_0_59 <= _GEN_2390;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_60 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_60 <= _GEN_515;
        end else begin
          ram_0_60 <= _GEN_2391;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_61 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_61 <= _GEN_516;
        end else begin
          ram_0_61 <= _GEN_2392;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_62 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_62 <= _GEN_517;
        end else begin
          ram_0_62 <= _GEN_2393;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_63 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          ram_0_63 <= _GEN_518;
        end else begin
          ram_0_63 <= _GEN_2394;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_0 <= _GEN_2395;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_1 <= _GEN_2396;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_2 <= _GEN_2397;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_3 <= _GEN_2398;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_4 <= _GEN_2399;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_5 <= _GEN_2400;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_6 <= _GEN_2401;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_7 <= _GEN_2402;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_8 <= _GEN_2403;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_9 <= _GEN_2404;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_10 <= _GEN_2405;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_11 <= _GEN_2406;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_12 <= _GEN_2407;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_13 <= _GEN_2408;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_14 <= _GEN_2409;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_15 <= _GEN_2410;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_16 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_16 <= _GEN_2411;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_17 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_17 <= _GEN_2412;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_18 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_18 <= _GEN_2413;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_19 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_19 <= _GEN_2414;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_20 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_20 <= _GEN_2415;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_21 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_21 <= _GEN_2416;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_22 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_22 <= _GEN_2417;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_23 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_23 <= _GEN_2418;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_24 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_24 <= _GEN_2419;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_25 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_25 <= _GEN_2420;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_26 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_26 <= _GEN_2421;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_27 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_27 <= _GEN_2422;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_28 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_28 <= _GEN_2423;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_29 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_29 <= _GEN_2424;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_30 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_30 <= _GEN_2425;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_31 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_31 <= _GEN_2426;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_32 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_32 <= _GEN_2427;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_33 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_33 <= _GEN_2428;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_34 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_34 <= _GEN_2429;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_35 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_35 <= _GEN_2430;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_36 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_36 <= _GEN_2431;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_37 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_37 <= _GEN_2432;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_38 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_38 <= _GEN_2433;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_39 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_39 <= _GEN_2434;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_40 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_40 <= _GEN_2435;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_41 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_41 <= _GEN_2436;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_42 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_42 <= _GEN_2437;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_43 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_43 <= _GEN_2438;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_44 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_44 <= _GEN_2439;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_45 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_45 <= _GEN_2440;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_46 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_46 <= _GEN_2441;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_47 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_47 <= _GEN_2442;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_48 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_48 <= _GEN_2443;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_49 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_49 <= _GEN_2444;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_50 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_50 <= _GEN_2445;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_51 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_51 <= _GEN_2446;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_52 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_52 <= _GEN_2447;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_53 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_53 <= _GEN_2448;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_54 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_54 <= _GEN_2449;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_55 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_55 <= _GEN_2450;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_56 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_56 <= _GEN_2451;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_57 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_57 <= _GEN_2452;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_58 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_58 <= _GEN_2453;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_59 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_59 <= _GEN_2454;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_60 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_60 <= _GEN_2455;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_61 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_61 <= _GEN_2456;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_62 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_62 <= _GEN_2457;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_63 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          tag_0_63 <= _GEN_2458;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_0 <= _GEN_519;
        end else begin
          valid_0_0 <= _GEN_2459;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_1 <= _GEN_520;
        end else begin
          valid_0_1 <= _GEN_2460;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_2 <= _GEN_521;
        end else begin
          valid_0_2 <= _GEN_2461;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_3 <= _GEN_522;
        end else begin
          valid_0_3 <= _GEN_2462;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_4 <= _GEN_523;
        end else begin
          valid_0_4 <= _GEN_2463;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_5 <= _GEN_524;
        end else begin
          valid_0_5 <= _GEN_2464;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_6 <= _GEN_525;
        end else begin
          valid_0_6 <= _GEN_2465;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_7 <= _GEN_526;
        end else begin
          valid_0_7 <= _GEN_2466;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_8 <= _GEN_527;
        end else begin
          valid_0_8 <= _GEN_2467;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_9 <= _GEN_528;
        end else begin
          valid_0_9 <= _GEN_2468;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_10 <= _GEN_529;
        end else begin
          valid_0_10 <= _GEN_2469;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_11 <= _GEN_530;
        end else begin
          valid_0_11 <= _GEN_2470;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_12 <= _GEN_531;
        end else begin
          valid_0_12 <= _GEN_2471;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_13 <= _GEN_532;
        end else begin
          valid_0_13 <= _GEN_2472;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_14 <= _GEN_533;
        end else begin
          valid_0_14 <= _GEN_2473;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_15 <= _GEN_534;
        end else begin
          valid_0_15 <= _GEN_2474;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_16 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_16 <= _GEN_535;
        end else begin
          valid_0_16 <= _GEN_2475;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_17 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_17 <= _GEN_536;
        end else begin
          valid_0_17 <= _GEN_2476;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_18 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_18 <= _GEN_537;
        end else begin
          valid_0_18 <= _GEN_2477;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_19 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_19 <= _GEN_538;
        end else begin
          valid_0_19 <= _GEN_2478;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_20 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_20 <= _GEN_539;
        end else begin
          valid_0_20 <= _GEN_2479;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_21 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_21 <= _GEN_540;
        end else begin
          valid_0_21 <= _GEN_2480;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_22 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_22 <= _GEN_541;
        end else begin
          valid_0_22 <= _GEN_2481;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_23 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_23 <= _GEN_542;
        end else begin
          valid_0_23 <= _GEN_2482;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_24 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_24 <= _GEN_543;
        end else begin
          valid_0_24 <= _GEN_2483;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_25 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_25 <= _GEN_544;
        end else begin
          valid_0_25 <= _GEN_2484;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_26 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_26 <= _GEN_545;
        end else begin
          valid_0_26 <= _GEN_2485;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_27 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_27 <= _GEN_546;
        end else begin
          valid_0_27 <= _GEN_2486;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_28 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_28 <= _GEN_547;
        end else begin
          valid_0_28 <= _GEN_2487;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_29 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_29 <= _GEN_548;
        end else begin
          valid_0_29 <= _GEN_2488;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_30 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_30 <= _GEN_549;
        end else begin
          valid_0_30 <= _GEN_2489;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_31 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_31 <= _GEN_550;
        end else begin
          valid_0_31 <= _GEN_2490;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_32 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_32 <= _GEN_551;
        end else begin
          valid_0_32 <= _GEN_2491;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_33 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_33 <= _GEN_552;
        end else begin
          valid_0_33 <= _GEN_2492;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_34 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_34 <= _GEN_553;
        end else begin
          valid_0_34 <= _GEN_2493;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_35 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_35 <= _GEN_554;
        end else begin
          valid_0_35 <= _GEN_2494;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_36 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_36 <= _GEN_555;
        end else begin
          valid_0_36 <= _GEN_2495;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_37 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_37 <= _GEN_556;
        end else begin
          valid_0_37 <= _GEN_2496;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_38 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_38 <= _GEN_557;
        end else begin
          valid_0_38 <= _GEN_2497;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_39 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_39 <= _GEN_558;
        end else begin
          valid_0_39 <= _GEN_2498;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_40 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_40 <= _GEN_559;
        end else begin
          valid_0_40 <= _GEN_2499;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_41 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_41 <= _GEN_560;
        end else begin
          valid_0_41 <= _GEN_2500;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_42 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_42 <= _GEN_561;
        end else begin
          valid_0_42 <= _GEN_2501;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_43 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_43 <= _GEN_562;
        end else begin
          valid_0_43 <= _GEN_2502;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_44 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_44 <= _GEN_563;
        end else begin
          valid_0_44 <= _GEN_2503;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_45 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_45 <= _GEN_564;
        end else begin
          valid_0_45 <= _GEN_2504;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_46 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_46 <= _GEN_565;
        end else begin
          valid_0_46 <= _GEN_2505;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_47 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_47 <= _GEN_566;
        end else begin
          valid_0_47 <= _GEN_2506;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_48 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_48 <= _GEN_567;
        end else begin
          valid_0_48 <= _GEN_2507;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_49 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_49 <= _GEN_568;
        end else begin
          valid_0_49 <= _GEN_2508;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_50 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_50 <= _GEN_569;
        end else begin
          valid_0_50 <= _GEN_2509;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_51 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_51 <= _GEN_570;
        end else begin
          valid_0_51 <= _GEN_2510;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_52 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_52 <= _GEN_571;
        end else begin
          valid_0_52 <= _GEN_2511;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_53 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_53 <= _GEN_572;
        end else begin
          valid_0_53 <= _GEN_2512;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_54 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_54 <= _GEN_573;
        end else begin
          valid_0_54 <= _GEN_2513;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_55 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_55 <= _GEN_574;
        end else begin
          valid_0_55 <= _GEN_2514;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_56 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_56 <= _GEN_575;
        end else begin
          valid_0_56 <= _GEN_2515;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_57 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_57 <= _GEN_576;
        end else begin
          valid_0_57 <= _GEN_2516;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_58 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_58 <= _GEN_577;
        end else begin
          valid_0_58 <= _GEN_2517;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_59 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_59 <= _GEN_578;
        end else begin
          valid_0_59 <= _GEN_2518;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_60 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_60 <= _GEN_579;
        end else begin
          valid_0_60 <= _GEN_2519;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_61 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_61 <= _GEN_580;
        end else begin
          valid_0_61 <= _GEN_2520;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_62 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_62 <= _GEN_581;
        end else begin
          valid_0_62 <= _GEN_2521;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_63 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          valid_0_63 <= _GEN_582;
        end else begin
          valid_0_63 <= _GEN_2522;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_0 <= _GEN_583;
        end else begin
          dirty_0_0 <= _GEN_2525;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_1 <= _GEN_584;
        end else begin
          dirty_0_1 <= _GEN_2526;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_2 <= _GEN_585;
        end else begin
          dirty_0_2 <= _GEN_2527;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_3 <= _GEN_586;
        end else begin
          dirty_0_3 <= _GEN_2528;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_4 <= _GEN_587;
        end else begin
          dirty_0_4 <= _GEN_2529;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_5 <= _GEN_588;
        end else begin
          dirty_0_5 <= _GEN_2530;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_6 <= _GEN_589;
        end else begin
          dirty_0_6 <= _GEN_2531;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_7 <= _GEN_590;
        end else begin
          dirty_0_7 <= _GEN_2532;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_8 <= _GEN_591;
        end else begin
          dirty_0_8 <= _GEN_2533;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_9 <= _GEN_592;
        end else begin
          dirty_0_9 <= _GEN_2534;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_10 <= _GEN_593;
        end else begin
          dirty_0_10 <= _GEN_2535;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_11 <= _GEN_594;
        end else begin
          dirty_0_11 <= _GEN_2536;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_12 <= _GEN_595;
        end else begin
          dirty_0_12 <= _GEN_2537;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_13 <= _GEN_596;
        end else begin
          dirty_0_13 <= _GEN_2538;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_14 <= _GEN_597;
        end else begin
          dirty_0_14 <= _GEN_2539;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_15 <= _GEN_598;
        end else begin
          dirty_0_15 <= _GEN_2540;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_16 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_16 <= _GEN_599;
        end else begin
          dirty_0_16 <= _GEN_2541;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_17 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_17 <= _GEN_600;
        end else begin
          dirty_0_17 <= _GEN_2542;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_18 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_18 <= _GEN_601;
        end else begin
          dirty_0_18 <= _GEN_2543;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_19 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_19 <= _GEN_602;
        end else begin
          dirty_0_19 <= _GEN_2544;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_20 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_20 <= _GEN_603;
        end else begin
          dirty_0_20 <= _GEN_2545;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_21 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_21 <= _GEN_604;
        end else begin
          dirty_0_21 <= _GEN_2546;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_22 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_22 <= _GEN_605;
        end else begin
          dirty_0_22 <= _GEN_2547;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_23 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_23 <= _GEN_606;
        end else begin
          dirty_0_23 <= _GEN_2548;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_24 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_24 <= _GEN_607;
        end else begin
          dirty_0_24 <= _GEN_2549;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_25 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_25 <= _GEN_608;
        end else begin
          dirty_0_25 <= _GEN_2550;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_26 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_26 <= _GEN_609;
        end else begin
          dirty_0_26 <= _GEN_2551;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_27 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_27 <= _GEN_610;
        end else begin
          dirty_0_27 <= _GEN_2552;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_28 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_28 <= _GEN_611;
        end else begin
          dirty_0_28 <= _GEN_2553;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_29 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_29 <= _GEN_612;
        end else begin
          dirty_0_29 <= _GEN_2554;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_30 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_30 <= _GEN_613;
        end else begin
          dirty_0_30 <= _GEN_2555;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_31 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_31 <= _GEN_614;
        end else begin
          dirty_0_31 <= _GEN_2556;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_32 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_32 <= _GEN_615;
        end else begin
          dirty_0_32 <= _GEN_2557;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_33 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_33 <= _GEN_616;
        end else begin
          dirty_0_33 <= _GEN_2558;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_34 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_34 <= _GEN_617;
        end else begin
          dirty_0_34 <= _GEN_2559;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_35 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_35 <= _GEN_618;
        end else begin
          dirty_0_35 <= _GEN_2560;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_36 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_36 <= _GEN_619;
        end else begin
          dirty_0_36 <= _GEN_2561;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_37 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_37 <= _GEN_620;
        end else begin
          dirty_0_37 <= _GEN_2562;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_38 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_38 <= _GEN_621;
        end else begin
          dirty_0_38 <= _GEN_2563;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_39 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_39 <= _GEN_622;
        end else begin
          dirty_0_39 <= _GEN_2564;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_40 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_40 <= _GEN_623;
        end else begin
          dirty_0_40 <= _GEN_2565;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_41 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_41 <= _GEN_624;
        end else begin
          dirty_0_41 <= _GEN_2566;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_42 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_42 <= _GEN_625;
        end else begin
          dirty_0_42 <= _GEN_2567;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_43 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_43 <= _GEN_626;
        end else begin
          dirty_0_43 <= _GEN_2568;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_44 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_44 <= _GEN_627;
        end else begin
          dirty_0_44 <= _GEN_2569;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_45 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_45 <= _GEN_628;
        end else begin
          dirty_0_45 <= _GEN_2570;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_46 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_46 <= _GEN_629;
        end else begin
          dirty_0_46 <= _GEN_2571;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_47 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_47 <= _GEN_630;
        end else begin
          dirty_0_47 <= _GEN_2572;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_48 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_48 <= _GEN_631;
        end else begin
          dirty_0_48 <= _GEN_2573;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_49 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_49 <= _GEN_632;
        end else begin
          dirty_0_49 <= _GEN_2574;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_50 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_50 <= _GEN_633;
        end else begin
          dirty_0_50 <= _GEN_2575;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_51 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_51 <= _GEN_634;
        end else begin
          dirty_0_51 <= _GEN_2576;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_52 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_52 <= _GEN_635;
        end else begin
          dirty_0_52 <= _GEN_2577;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_53 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_53 <= _GEN_636;
        end else begin
          dirty_0_53 <= _GEN_2578;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_54 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_54 <= _GEN_637;
        end else begin
          dirty_0_54 <= _GEN_2579;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_55 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_55 <= _GEN_638;
        end else begin
          dirty_0_55 <= _GEN_2580;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_56 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_56 <= _GEN_639;
        end else begin
          dirty_0_56 <= _GEN_2581;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_57 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_57 <= _GEN_640;
        end else begin
          dirty_0_57 <= _GEN_2582;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_58 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_58 <= _GEN_641;
        end else begin
          dirty_0_58 <= _GEN_2583;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_59 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_59 <= _GEN_642;
        end else begin
          dirty_0_59 <= _GEN_2584;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_60 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_60 <= _GEN_643;
        end else begin
          dirty_0_60 <= _GEN_2585;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_61 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_61 <= _GEN_644;
        end else begin
          dirty_0_61 <= _GEN_2586;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_62 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_62 <= _GEN_645;
        end else begin
          dirty_0_62 <= _GEN_2587;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_63 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (3'h2 == state) begin // @[d_cache.scala 81:18]
          dirty_0_63 <= _GEN_646;
        end else begin
          dirty_0_63 <= _GEN_2588;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 28:27]
      way0_hit <= 1'h0; // @[d_cache.scala 28:27]
    end else begin
      way0_hit <= _T_4;
    end
    if (reset) begin // @[d_cache.scala 31:34]
      write_back_data <= 64'h0; // @[d_cache.scala 31:34]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          write_back_data <= _GEN_2523;
        end
      end
    end
    write_back_addr <= _GEN_3784[31:0]; // @[d_cache.scala 32:{34,34}]
    if (reset) begin // @[d_cache.scala 35:28]
      unuse_way <= 2'h0; // @[d_cache.scala 35:28]
    end else begin
      unuse_way <= {{1'd0}, _T_5};
    end
    if (reset) begin // @[d_cache.scala 36:31]
      receive_data <= 64'h0; // @[d_cache.scala 36:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 81:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 81:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 81:18]
          receive_data <= _GEN_2330;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 76:24]
      state <= 3'h0; // @[d_cache.scala 76:24]
    end else if (3'h0 == state) begin // @[d_cache.scala 81:18]
      if (io_from_lsu_arvalid) begin // @[d_cache.scala 83:38]
        state <= 3'h1; // @[d_cache.scala 84:23]
      end else if (io_from_lsu_awvalid) begin // @[d_cache.scala 85:44]
        state <= 3'h2; // @[d_cache.scala 86:23]
      end
    end else if (3'h1 == state) begin // @[d_cache.scala 81:18]
      if (way0_hit) begin // @[d_cache.scala 91:27]
        state <= _GEN_196;
      end else begin
        state <= 3'h3; // @[d_cache.scala 103:23]
      end
    end else if (3'h2 == state) begin // @[d_cache.scala 81:18]
      state <= _GEN_454;
    end else begin
      state <= _GEN_2329;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"read addr : %x  write addr : %x\n",io_from_lsu_araddr,io_from_lsu_awaddr); // @[d_cache.scala 15:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"d_cache state:%d\n",state); // @[d_cache.scala 77:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"receive data:%x\n",receive_data); // @[d_cache.scala 79:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_10 & _T_11 & way0_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_0:%d\n",6'h3f == index ? dirty_0_63 : _GEN_194); // @[d_cache.scala 93:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"cacheline0:%x  \n",_GEN_261); // @[d_cache.scala 364:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {1{`RANDOM}};
  tag_0_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  tag_0_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  tag_0_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  tag_0_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  tag_0_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  tag_0_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  tag_0_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  tag_0_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  tag_0_8 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  tag_0_9 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  tag_0_10 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  tag_0_11 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  tag_0_12 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  tag_0_13 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  tag_0_14 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  tag_0_15 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  tag_0_16 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  tag_0_17 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  tag_0_18 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  tag_0_19 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  tag_0_20 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  tag_0_21 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  tag_0_22 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  tag_0_23 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  tag_0_24 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  tag_0_25 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  tag_0_26 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  tag_0_27 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  tag_0_28 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  tag_0_29 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  tag_0_30 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  tag_0_31 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  tag_0_32 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  tag_0_33 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  tag_0_34 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  tag_0_35 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  tag_0_36 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  tag_0_37 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  tag_0_38 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  tag_0_39 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  tag_0_40 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  tag_0_41 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  tag_0_42 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  tag_0_43 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  tag_0_44 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  tag_0_45 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  tag_0_46 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  tag_0_47 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  tag_0_48 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  tag_0_49 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  tag_0_50 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  tag_0_51 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  tag_0_52 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  tag_0_53 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  tag_0_54 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  tag_0_55 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  tag_0_56 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  tag_0_57 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  tag_0_58 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  tag_0_59 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  tag_0_60 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  tag_0_61 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  tag_0_62 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  tag_0_63 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_0_16 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_0_17 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_0_18 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_0_19 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_0_20 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_0_21 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_0_22 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_0_23 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_0_24 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_0_25 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_0_26 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_0_27 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_0_28 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_0_29 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_0_30 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_0_31 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_0_32 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_0_33 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_0_34 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_0_35 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_0_36 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_0_37 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_0_38 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_0_39 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_0_40 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_0_41 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_0_42 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_0_43 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_0_44 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_0_45 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_0_46 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_0_47 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_0_48 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_0_49 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_0_50 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_0_51 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_0_52 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_0_53 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_0_54 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_0_55 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_0_56 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_0_57 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_0_58 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_0_59 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_0_60 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_0_61 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_0_62 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_0_63 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  dirty_0_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  dirty_0_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dirty_0_2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  dirty_0_3 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  dirty_0_4 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  dirty_0_5 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  dirty_0_6 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  dirty_0_7 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dirty_0_8 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  dirty_0_9 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  dirty_0_10 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  dirty_0_11 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  dirty_0_12 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  dirty_0_13 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dirty_0_14 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  dirty_0_15 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  dirty_0_16 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  dirty_0_17 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  dirty_0_18 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  dirty_0_19 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dirty_0_20 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  dirty_0_21 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  dirty_0_22 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  dirty_0_23 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  dirty_0_24 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  dirty_0_25 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  dirty_0_26 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  dirty_0_27 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  dirty_0_28 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  dirty_0_29 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  dirty_0_30 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  dirty_0_31 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  dirty_0_32 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  dirty_0_33 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  dirty_0_34 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  dirty_0_35 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  dirty_0_36 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  dirty_0_37 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  dirty_0_38 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  dirty_0_39 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  dirty_0_40 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  dirty_0_41 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  dirty_0_42 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  dirty_0_43 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  dirty_0_44 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  dirty_0_45 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  dirty_0_46 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  dirty_0_47 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  dirty_0_48 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  dirty_0_49 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  dirty_0_50 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  dirty_0_51 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  dirty_0_52 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  dirty_0_53 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  dirty_0_54 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  dirty_0_55 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  dirty_0_56 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  dirty_0_57 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  dirty_0_58 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  dirty_0_59 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  dirty_0_60 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  dirty_0_61 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  dirty_0_62 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  dirty_0_63 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  way0_hit = _RAND_256[0:0];
  _RAND_257 = {2{`RANDOM}};
  write_back_data = _RAND_257[63:0];
  _RAND_258 = {1{`RANDOM}};
  write_back_addr = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  unuse_way = _RAND_259[1:0];
  _RAND_260 = {2{`RANDOM}};
  receive_data = _RAND_260[63:0];
  _RAND_261 = {1{`RANDOM}};
  state = _RAND_261[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
