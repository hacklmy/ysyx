module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input         io_from_lsu_rready,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [31:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  input         io_from_lsu_bready,
  output        io_to_lsu_arready,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_awready,
  output        io_to_lsu_wready,
  output        io_to_lsu_bvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output        io_to_axi_awvalid,
  output [31:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input         io_from_axi_arready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid,
  input         io_from_axi_awready,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [63:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [63:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = ~reset; // @[d_cache.scala 15:11]
  reg [63:0] ram_0_0; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_1; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_2; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_3; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_4; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_5; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_6; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_7; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_8; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_9; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_10; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_11; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_12; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_13; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_14; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_15; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_16; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_17; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_18; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_19; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_20; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_21; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_22; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_23; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_24; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_25; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_26; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_27; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_28; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_29; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_30; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_31; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_32; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_33; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_34; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_35; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_36; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_37; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_38; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_39; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_40; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_41; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_42; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_43; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_44; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_45; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_46; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_47; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_48; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_49; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_50; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_51; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_52; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_53; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_54; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_55; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_56; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_57; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_58; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_59; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_60; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_61; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_62; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_63; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_64; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_65; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_66; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_67; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_68; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_69; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_70; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_71; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_72; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_73; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_74; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_75; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_76; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_77; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_78; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_79; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_80; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_81; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_82; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_83; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_84; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_85; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_86; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_87; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_88; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_89; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_90; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_91; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_92; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_93; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_94; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_95; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_96; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_97; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_98; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_99; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_100; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_101; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_102; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_103; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_104; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_105; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_106; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_107; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_108; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_109; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_110; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_111; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_112; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_113; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_114; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_115; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_116; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_117; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_118; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_119; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_120; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_121; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_122; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_123; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_124; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_125; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_126; // @[d_cache.scala 18:24]
  reg [63:0] ram_0_127; // @[d_cache.scala 18:24]
  reg [63:0] ram_1_0; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_1; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_2; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_3; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_4; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_5; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_6; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_7; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_8; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_9; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_10; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_11; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_12; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_13; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_14; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_15; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_16; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_17; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_18; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_19; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_20; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_21; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_22; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_23; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_24; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_25; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_26; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_27; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_28; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_29; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_30; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_31; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_32; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_33; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_34; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_35; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_36; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_37; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_38; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_39; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_40; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_41; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_42; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_43; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_44; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_45; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_46; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_47; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_48; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_49; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_50; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_51; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_52; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_53; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_54; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_55; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_56; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_57; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_58; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_59; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_60; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_61; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_62; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_63; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_64; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_65; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_66; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_67; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_68; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_69; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_70; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_71; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_72; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_73; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_74; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_75; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_76; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_77; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_78; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_79; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_80; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_81; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_82; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_83; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_84; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_85; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_86; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_87; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_88; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_89; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_90; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_91; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_92; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_93; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_94; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_95; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_96; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_97; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_98; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_99; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_100; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_101; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_102; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_103; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_104; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_105; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_106; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_107; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_108; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_109; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_110; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_111; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_112; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_113; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_114; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_115; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_116; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_117; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_118; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_119; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_120; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_121; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_122; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_123; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_124; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_125; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_126; // @[d_cache.scala 19:24]
  reg [63:0] ram_1_127; // @[d_cache.scala 19:24]
  reg [31:0] tag_0_0; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_16; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_17; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_18; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_19; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_20; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_21; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_22; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_23; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_24; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_25; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_26; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_27; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_28; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_29; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_30; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_31; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_32; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_33; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_34; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_35; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_36; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_37; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_38; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_39; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_40; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_41; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_42; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_43; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_44; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_45; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_46; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_47; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_48; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_49; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_50; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_51; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_52; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_53; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_54; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_55; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_56; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_57; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_58; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_59; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_60; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_61; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_62; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_63; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_64; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_65; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_66; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_67; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_68; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_69; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_70; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_71; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_72; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_73; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_74; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_75; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_76; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_77; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_78; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_79; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_80; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_81; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_82; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_83; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_84; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_85; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_86; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_87; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_88; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_89; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_90; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_91; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_92; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_93; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_94; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_95; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_96; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_97; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_98; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_99; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_100; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_101; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_102; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_103; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_104; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_105; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_106; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_107; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_108; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_109; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_110; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_111; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_112; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_113; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_114; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_115; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_116; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_117; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_118; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_119; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_120; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_121; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_122; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_123; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_124; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_125; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_126; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_127; // @[d_cache.scala 20:24]
  reg [31:0] tag_1_0; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_1; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_2; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_3; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_4; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_5; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_6; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_7; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_8; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_9; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_10; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_11; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_12; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_13; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_14; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_15; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_16; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_17; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_18; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_19; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_20; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_21; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_22; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_23; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_24; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_25; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_26; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_27; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_28; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_29; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_30; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_31; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_32; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_33; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_34; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_35; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_36; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_37; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_38; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_39; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_40; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_41; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_42; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_43; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_44; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_45; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_46; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_47; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_48; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_49; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_50; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_51; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_52; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_53; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_54; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_55; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_56; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_57; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_58; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_59; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_60; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_61; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_62; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_63; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_64; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_65; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_66; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_67; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_68; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_69; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_70; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_71; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_72; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_73; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_74; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_75; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_76; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_77; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_78; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_79; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_80; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_81; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_82; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_83; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_84; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_85; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_86; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_87; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_88; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_89; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_90; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_91; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_92; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_93; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_94; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_95; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_96; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_97; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_98; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_99; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_100; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_101; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_102; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_103; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_104; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_105; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_106; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_107; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_108; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_109; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_110; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_111; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_112; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_113; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_114; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_115; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_116; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_117; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_118; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_119; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_120; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_121; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_122; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_123; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_124; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_125; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_126; // @[d_cache.scala 21:24]
  reg [31:0] tag_1_127; // @[d_cache.scala 21:24]
  reg  valid_0_0; // @[d_cache.scala 22:26]
  reg  valid_0_1; // @[d_cache.scala 22:26]
  reg  valid_0_2; // @[d_cache.scala 22:26]
  reg  valid_0_3; // @[d_cache.scala 22:26]
  reg  valid_0_4; // @[d_cache.scala 22:26]
  reg  valid_0_5; // @[d_cache.scala 22:26]
  reg  valid_0_6; // @[d_cache.scala 22:26]
  reg  valid_0_7; // @[d_cache.scala 22:26]
  reg  valid_0_8; // @[d_cache.scala 22:26]
  reg  valid_0_9; // @[d_cache.scala 22:26]
  reg  valid_0_10; // @[d_cache.scala 22:26]
  reg  valid_0_11; // @[d_cache.scala 22:26]
  reg  valid_0_12; // @[d_cache.scala 22:26]
  reg  valid_0_13; // @[d_cache.scala 22:26]
  reg  valid_0_14; // @[d_cache.scala 22:26]
  reg  valid_0_15; // @[d_cache.scala 22:26]
  reg  valid_0_16; // @[d_cache.scala 22:26]
  reg  valid_0_17; // @[d_cache.scala 22:26]
  reg  valid_0_18; // @[d_cache.scala 22:26]
  reg  valid_0_19; // @[d_cache.scala 22:26]
  reg  valid_0_20; // @[d_cache.scala 22:26]
  reg  valid_0_21; // @[d_cache.scala 22:26]
  reg  valid_0_22; // @[d_cache.scala 22:26]
  reg  valid_0_23; // @[d_cache.scala 22:26]
  reg  valid_0_24; // @[d_cache.scala 22:26]
  reg  valid_0_25; // @[d_cache.scala 22:26]
  reg  valid_0_26; // @[d_cache.scala 22:26]
  reg  valid_0_27; // @[d_cache.scala 22:26]
  reg  valid_0_28; // @[d_cache.scala 22:26]
  reg  valid_0_29; // @[d_cache.scala 22:26]
  reg  valid_0_30; // @[d_cache.scala 22:26]
  reg  valid_0_31; // @[d_cache.scala 22:26]
  reg  valid_0_32; // @[d_cache.scala 22:26]
  reg  valid_0_33; // @[d_cache.scala 22:26]
  reg  valid_0_34; // @[d_cache.scala 22:26]
  reg  valid_0_35; // @[d_cache.scala 22:26]
  reg  valid_0_36; // @[d_cache.scala 22:26]
  reg  valid_0_37; // @[d_cache.scala 22:26]
  reg  valid_0_38; // @[d_cache.scala 22:26]
  reg  valid_0_39; // @[d_cache.scala 22:26]
  reg  valid_0_40; // @[d_cache.scala 22:26]
  reg  valid_0_41; // @[d_cache.scala 22:26]
  reg  valid_0_42; // @[d_cache.scala 22:26]
  reg  valid_0_43; // @[d_cache.scala 22:26]
  reg  valid_0_44; // @[d_cache.scala 22:26]
  reg  valid_0_45; // @[d_cache.scala 22:26]
  reg  valid_0_46; // @[d_cache.scala 22:26]
  reg  valid_0_47; // @[d_cache.scala 22:26]
  reg  valid_0_48; // @[d_cache.scala 22:26]
  reg  valid_0_49; // @[d_cache.scala 22:26]
  reg  valid_0_50; // @[d_cache.scala 22:26]
  reg  valid_0_51; // @[d_cache.scala 22:26]
  reg  valid_0_52; // @[d_cache.scala 22:26]
  reg  valid_0_53; // @[d_cache.scala 22:26]
  reg  valid_0_54; // @[d_cache.scala 22:26]
  reg  valid_0_55; // @[d_cache.scala 22:26]
  reg  valid_0_56; // @[d_cache.scala 22:26]
  reg  valid_0_57; // @[d_cache.scala 22:26]
  reg  valid_0_58; // @[d_cache.scala 22:26]
  reg  valid_0_59; // @[d_cache.scala 22:26]
  reg  valid_0_60; // @[d_cache.scala 22:26]
  reg  valid_0_61; // @[d_cache.scala 22:26]
  reg  valid_0_62; // @[d_cache.scala 22:26]
  reg  valid_0_63; // @[d_cache.scala 22:26]
  reg  valid_0_64; // @[d_cache.scala 22:26]
  reg  valid_0_65; // @[d_cache.scala 22:26]
  reg  valid_0_66; // @[d_cache.scala 22:26]
  reg  valid_0_67; // @[d_cache.scala 22:26]
  reg  valid_0_68; // @[d_cache.scala 22:26]
  reg  valid_0_69; // @[d_cache.scala 22:26]
  reg  valid_0_70; // @[d_cache.scala 22:26]
  reg  valid_0_71; // @[d_cache.scala 22:26]
  reg  valid_0_72; // @[d_cache.scala 22:26]
  reg  valid_0_73; // @[d_cache.scala 22:26]
  reg  valid_0_74; // @[d_cache.scala 22:26]
  reg  valid_0_75; // @[d_cache.scala 22:26]
  reg  valid_0_76; // @[d_cache.scala 22:26]
  reg  valid_0_77; // @[d_cache.scala 22:26]
  reg  valid_0_78; // @[d_cache.scala 22:26]
  reg  valid_0_79; // @[d_cache.scala 22:26]
  reg  valid_0_80; // @[d_cache.scala 22:26]
  reg  valid_0_81; // @[d_cache.scala 22:26]
  reg  valid_0_82; // @[d_cache.scala 22:26]
  reg  valid_0_83; // @[d_cache.scala 22:26]
  reg  valid_0_84; // @[d_cache.scala 22:26]
  reg  valid_0_85; // @[d_cache.scala 22:26]
  reg  valid_0_86; // @[d_cache.scala 22:26]
  reg  valid_0_87; // @[d_cache.scala 22:26]
  reg  valid_0_88; // @[d_cache.scala 22:26]
  reg  valid_0_89; // @[d_cache.scala 22:26]
  reg  valid_0_90; // @[d_cache.scala 22:26]
  reg  valid_0_91; // @[d_cache.scala 22:26]
  reg  valid_0_92; // @[d_cache.scala 22:26]
  reg  valid_0_93; // @[d_cache.scala 22:26]
  reg  valid_0_94; // @[d_cache.scala 22:26]
  reg  valid_0_95; // @[d_cache.scala 22:26]
  reg  valid_0_96; // @[d_cache.scala 22:26]
  reg  valid_0_97; // @[d_cache.scala 22:26]
  reg  valid_0_98; // @[d_cache.scala 22:26]
  reg  valid_0_99; // @[d_cache.scala 22:26]
  reg  valid_0_100; // @[d_cache.scala 22:26]
  reg  valid_0_101; // @[d_cache.scala 22:26]
  reg  valid_0_102; // @[d_cache.scala 22:26]
  reg  valid_0_103; // @[d_cache.scala 22:26]
  reg  valid_0_104; // @[d_cache.scala 22:26]
  reg  valid_0_105; // @[d_cache.scala 22:26]
  reg  valid_0_106; // @[d_cache.scala 22:26]
  reg  valid_0_107; // @[d_cache.scala 22:26]
  reg  valid_0_108; // @[d_cache.scala 22:26]
  reg  valid_0_109; // @[d_cache.scala 22:26]
  reg  valid_0_110; // @[d_cache.scala 22:26]
  reg  valid_0_111; // @[d_cache.scala 22:26]
  reg  valid_0_112; // @[d_cache.scala 22:26]
  reg  valid_0_113; // @[d_cache.scala 22:26]
  reg  valid_0_114; // @[d_cache.scala 22:26]
  reg  valid_0_115; // @[d_cache.scala 22:26]
  reg  valid_0_116; // @[d_cache.scala 22:26]
  reg  valid_0_117; // @[d_cache.scala 22:26]
  reg  valid_0_118; // @[d_cache.scala 22:26]
  reg  valid_0_119; // @[d_cache.scala 22:26]
  reg  valid_0_120; // @[d_cache.scala 22:26]
  reg  valid_0_121; // @[d_cache.scala 22:26]
  reg  valid_0_122; // @[d_cache.scala 22:26]
  reg  valid_0_123; // @[d_cache.scala 22:26]
  reg  valid_0_124; // @[d_cache.scala 22:26]
  reg  valid_0_125; // @[d_cache.scala 22:26]
  reg  valid_0_126; // @[d_cache.scala 22:26]
  reg  valid_0_127; // @[d_cache.scala 22:26]
  reg  valid_1_0; // @[d_cache.scala 23:26]
  reg  valid_1_1; // @[d_cache.scala 23:26]
  reg  valid_1_2; // @[d_cache.scala 23:26]
  reg  valid_1_3; // @[d_cache.scala 23:26]
  reg  valid_1_4; // @[d_cache.scala 23:26]
  reg  valid_1_5; // @[d_cache.scala 23:26]
  reg  valid_1_6; // @[d_cache.scala 23:26]
  reg  valid_1_7; // @[d_cache.scala 23:26]
  reg  valid_1_8; // @[d_cache.scala 23:26]
  reg  valid_1_9; // @[d_cache.scala 23:26]
  reg  valid_1_10; // @[d_cache.scala 23:26]
  reg  valid_1_11; // @[d_cache.scala 23:26]
  reg  valid_1_12; // @[d_cache.scala 23:26]
  reg  valid_1_13; // @[d_cache.scala 23:26]
  reg  valid_1_14; // @[d_cache.scala 23:26]
  reg  valid_1_15; // @[d_cache.scala 23:26]
  reg  valid_1_16; // @[d_cache.scala 23:26]
  reg  valid_1_17; // @[d_cache.scala 23:26]
  reg  valid_1_18; // @[d_cache.scala 23:26]
  reg  valid_1_19; // @[d_cache.scala 23:26]
  reg  valid_1_20; // @[d_cache.scala 23:26]
  reg  valid_1_21; // @[d_cache.scala 23:26]
  reg  valid_1_22; // @[d_cache.scala 23:26]
  reg  valid_1_23; // @[d_cache.scala 23:26]
  reg  valid_1_24; // @[d_cache.scala 23:26]
  reg  valid_1_25; // @[d_cache.scala 23:26]
  reg  valid_1_26; // @[d_cache.scala 23:26]
  reg  valid_1_27; // @[d_cache.scala 23:26]
  reg  valid_1_28; // @[d_cache.scala 23:26]
  reg  valid_1_29; // @[d_cache.scala 23:26]
  reg  valid_1_30; // @[d_cache.scala 23:26]
  reg  valid_1_31; // @[d_cache.scala 23:26]
  reg  valid_1_32; // @[d_cache.scala 23:26]
  reg  valid_1_33; // @[d_cache.scala 23:26]
  reg  valid_1_34; // @[d_cache.scala 23:26]
  reg  valid_1_35; // @[d_cache.scala 23:26]
  reg  valid_1_36; // @[d_cache.scala 23:26]
  reg  valid_1_37; // @[d_cache.scala 23:26]
  reg  valid_1_38; // @[d_cache.scala 23:26]
  reg  valid_1_39; // @[d_cache.scala 23:26]
  reg  valid_1_40; // @[d_cache.scala 23:26]
  reg  valid_1_41; // @[d_cache.scala 23:26]
  reg  valid_1_42; // @[d_cache.scala 23:26]
  reg  valid_1_43; // @[d_cache.scala 23:26]
  reg  valid_1_44; // @[d_cache.scala 23:26]
  reg  valid_1_45; // @[d_cache.scala 23:26]
  reg  valid_1_46; // @[d_cache.scala 23:26]
  reg  valid_1_47; // @[d_cache.scala 23:26]
  reg  valid_1_48; // @[d_cache.scala 23:26]
  reg  valid_1_49; // @[d_cache.scala 23:26]
  reg  valid_1_50; // @[d_cache.scala 23:26]
  reg  valid_1_51; // @[d_cache.scala 23:26]
  reg  valid_1_52; // @[d_cache.scala 23:26]
  reg  valid_1_53; // @[d_cache.scala 23:26]
  reg  valid_1_54; // @[d_cache.scala 23:26]
  reg  valid_1_55; // @[d_cache.scala 23:26]
  reg  valid_1_56; // @[d_cache.scala 23:26]
  reg  valid_1_57; // @[d_cache.scala 23:26]
  reg  valid_1_58; // @[d_cache.scala 23:26]
  reg  valid_1_59; // @[d_cache.scala 23:26]
  reg  valid_1_60; // @[d_cache.scala 23:26]
  reg  valid_1_61; // @[d_cache.scala 23:26]
  reg  valid_1_62; // @[d_cache.scala 23:26]
  reg  valid_1_63; // @[d_cache.scala 23:26]
  reg  valid_1_64; // @[d_cache.scala 23:26]
  reg  valid_1_65; // @[d_cache.scala 23:26]
  reg  valid_1_66; // @[d_cache.scala 23:26]
  reg  valid_1_67; // @[d_cache.scala 23:26]
  reg  valid_1_68; // @[d_cache.scala 23:26]
  reg  valid_1_69; // @[d_cache.scala 23:26]
  reg  valid_1_70; // @[d_cache.scala 23:26]
  reg  valid_1_71; // @[d_cache.scala 23:26]
  reg  valid_1_72; // @[d_cache.scala 23:26]
  reg  valid_1_73; // @[d_cache.scala 23:26]
  reg  valid_1_74; // @[d_cache.scala 23:26]
  reg  valid_1_75; // @[d_cache.scala 23:26]
  reg  valid_1_76; // @[d_cache.scala 23:26]
  reg  valid_1_77; // @[d_cache.scala 23:26]
  reg  valid_1_78; // @[d_cache.scala 23:26]
  reg  valid_1_79; // @[d_cache.scala 23:26]
  reg  valid_1_80; // @[d_cache.scala 23:26]
  reg  valid_1_81; // @[d_cache.scala 23:26]
  reg  valid_1_82; // @[d_cache.scala 23:26]
  reg  valid_1_83; // @[d_cache.scala 23:26]
  reg  valid_1_84; // @[d_cache.scala 23:26]
  reg  valid_1_85; // @[d_cache.scala 23:26]
  reg  valid_1_86; // @[d_cache.scala 23:26]
  reg  valid_1_87; // @[d_cache.scala 23:26]
  reg  valid_1_88; // @[d_cache.scala 23:26]
  reg  valid_1_89; // @[d_cache.scala 23:26]
  reg  valid_1_90; // @[d_cache.scala 23:26]
  reg  valid_1_91; // @[d_cache.scala 23:26]
  reg  valid_1_92; // @[d_cache.scala 23:26]
  reg  valid_1_93; // @[d_cache.scala 23:26]
  reg  valid_1_94; // @[d_cache.scala 23:26]
  reg  valid_1_95; // @[d_cache.scala 23:26]
  reg  valid_1_96; // @[d_cache.scala 23:26]
  reg  valid_1_97; // @[d_cache.scala 23:26]
  reg  valid_1_98; // @[d_cache.scala 23:26]
  reg  valid_1_99; // @[d_cache.scala 23:26]
  reg  valid_1_100; // @[d_cache.scala 23:26]
  reg  valid_1_101; // @[d_cache.scala 23:26]
  reg  valid_1_102; // @[d_cache.scala 23:26]
  reg  valid_1_103; // @[d_cache.scala 23:26]
  reg  valid_1_104; // @[d_cache.scala 23:26]
  reg  valid_1_105; // @[d_cache.scala 23:26]
  reg  valid_1_106; // @[d_cache.scala 23:26]
  reg  valid_1_107; // @[d_cache.scala 23:26]
  reg  valid_1_108; // @[d_cache.scala 23:26]
  reg  valid_1_109; // @[d_cache.scala 23:26]
  reg  valid_1_110; // @[d_cache.scala 23:26]
  reg  valid_1_111; // @[d_cache.scala 23:26]
  reg  valid_1_112; // @[d_cache.scala 23:26]
  reg  valid_1_113; // @[d_cache.scala 23:26]
  reg  valid_1_114; // @[d_cache.scala 23:26]
  reg  valid_1_115; // @[d_cache.scala 23:26]
  reg  valid_1_116; // @[d_cache.scala 23:26]
  reg  valid_1_117; // @[d_cache.scala 23:26]
  reg  valid_1_118; // @[d_cache.scala 23:26]
  reg  valid_1_119; // @[d_cache.scala 23:26]
  reg  valid_1_120; // @[d_cache.scala 23:26]
  reg  valid_1_121; // @[d_cache.scala 23:26]
  reg  valid_1_122; // @[d_cache.scala 23:26]
  reg  valid_1_123; // @[d_cache.scala 23:26]
  reg  valid_1_124; // @[d_cache.scala 23:26]
  reg  valid_1_125; // @[d_cache.scala 23:26]
  reg  valid_1_126; // @[d_cache.scala 23:26]
  reg  valid_1_127; // @[d_cache.scala 23:26]
  reg  dirty_0_0; // @[d_cache.scala 24:26]
  reg  dirty_0_1; // @[d_cache.scala 24:26]
  reg  dirty_0_2; // @[d_cache.scala 24:26]
  reg  dirty_0_3; // @[d_cache.scala 24:26]
  reg  dirty_0_4; // @[d_cache.scala 24:26]
  reg  dirty_0_5; // @[d_cache.scala 24:26]
  reg  dirty_0_6; // @[d_cache.scala 24:26]
  reg  dirty_0_7; // @[d_cache.scala 24:26]
  reg  dirty_0_8; // @[d_cache.scala 24:26]
  reg  dirty_0_9; // @[d_cache.scala 24:26]
  reg  dirty_0_10; // @[d_cache.scala 24:26]
  reg  dirty_0_11; // @[d_cache.scala 24:26]
  reg  dirty_0_12; // @[d_cache.scala 24:26]
  reg  dirty_0_13; // @[d_cache.scala 24:26]
  reg  dirty_0_14; // @[d_cache.scala 24:26]
  reg  dirty_0_15; // @[d_cache.scala 24:26]
  reg  dirty_0_16; // @[d_cache.scala 24:26]
  reg  dirty_0_17; // @[d_cache.scala 24:26]
  reg  dirty_0_18; // @[d_cache.scala 24:26]
  reg  dirty_0_19; // @[d_cache.scala 24:26]
  reg  dirty_0_20; // @[d_cache.scala 24:26]
  reg  dirty_0_21; // @[d_cache.scala 24:26]
  reg  dirty_0_22; // @[d_cache.scala 24:26]
  reg  dirty_0_23; // @[d_cache.scala 24:26]
  reg  dirty_0_24; // @[d_cache.scala 24:26]
  reg  dirty_0_25; // @[d_cache.scala 24:26]
  reg  dirty_0_26; // @[d_cache.scala 24:26]
  reg  dirty_0_27; // @[d_cache.scala 24:26]
  reg  dirty_0_28; // @[d_cache.scala 24:26]
  reg  dirty_0_29; // @[d_cache.scala 24:26]
  reg  dirty_0_30; // @[d_cache.scala 24:26]
  reg  dirty_0_31; // @[d_cache.scala 24:26]
  reg  dirty_0_32; // @[d_cache.scala 24:26]
  reg  dirty_0_33; // @[d_cache.scala 24:26]
  reg  dirty_0_34; // @[d_cache.scala 24:26]
  reg  dirty_0_35; // @[d_cache.scala 24:26]
  reg  dirty_0_36; // @[d_cache.scala 24:26]
  reg  dirty_0_37; // @[d_cache.scala 24:26]
  reg  dirty_0_38; // @[d_cache.scala 24:26]
  reg  dirty_0_39; // @[d_cache.scala 24:26]
  reg  dirty_0_40; // @[d_cache.scala 24:26]
  reg  dirty_0_41; // @[d_cache.scala 24:26]
  reg  dirty_0_42; // @[d_cache.scala 24:26]
  reg  dirty_0_43; // @[d_cache.scala 24:26]
  reg  dirty_0_44; // @[d_cache.scala 24:26]
  reg  dirty_0_45; // @[d_cache.scala 24:26]
  reg  dirty_0_46; // @[d_cache.scala 24:26]
  reg  dirty_0_47; // @[d_cache.scala 24:26]
  reg  dirty_0_48; // @[d_cache.scala 24:26]
  reg  dirty_0_49; // @[d_cache.scala 24:26]
  reg  dirty_0_50; // @[d_cache.scala 24:26]
  reg  dirty_0_51; // @[d_cache.scala 24:26]
  reg  dirty_0_52; // @[d_cache.scala 24:26]
  reg  dirty_0_53; // @[d_cache.scala 24:26]
  reg  dirty_0_54; // @[d_cache.scala 24:26]
  reg  dirty_0_55; // @[d_cache.scala 24:26]
  reg  dirty_0_56; // @[d_cache.scala 24:26]
  reg  dirty_0_57; // @[d_cache.scala 24:26]
  reg  dirty_0_58; // @[d_cache.scala 24:26]
  reg  dirty_0_59; // @[d_cache.scala 24:26]
  reg  dirty_0_60; // @[d_cache.scala 24:26]
  reg  dirty_0_61; // @[d_cache.scala 24:26]
  reg  dirty_0_62; // @[d_cache.scala 24:26]
  reg  dirty_0_63; // @[d_cache.scala 24:26]
  reg  dirty_0_64; // @[d_cache.scala 24:26]
  reg  dirty_0_65; // @[d_cache.scala 24:26]
  reg  dirty_0_66; // @[d_cache.scala 24:26]
  reg  dirty_0_67; // @[d_cache.scala 24:26]
  reg  dirty_0_68; // @[d_cache.scala 24:26]
  reg  dirty_0_69; // @[d_cache.scala 24:26]
  reg  dirty_0_70; // @[d_cache.scala 24:26]
  reg  dirty_0_71; // @[d_cache.scala 24:26]
  reg  dirty_0_72; // @[d_cache.scala 24:26]
  reg  dirty_0_73; // @[d_cache.scala 24:26]
  reg  dirty_0_74; // @[d_cache.scala 24:26]
  reg  dirty_0_75; // @[d_cache.scala 24:26]
  reg  dirty_0_76; // @[d_cache.scala 24:26]
  reg  dirty_0_77; // @[d_cache.scala 24:26]
  reg  dirty_0_78; // @[d_cache.scala 24:26]
  reg  dirty_0_79; // @[d_cache.scala 24:26]
  reg  dirty_0_80; // @[d_cache.scala 24:26]
  reg  dirty_0_81; // @[d_cache.scala 24:26]
  reg  dirty_0_82; // @[d_cache.scala 24:26]
  reg  dirty_0_83; // @[d_cache.scala 24:26]
  reg  dirty_0_84; // @[d_cache.scala 24:26]
  reg  dirty_0_85; // @[d_cache.scala 24:26]
  reg  dirty_0_86; // @[d_cache.scala 24:26]
  reg  dirty_0_87; // @[d_cache.scala 24:26]
  reg  dirty_0_88; // @[d_cache.scala 24:26]
  reg  dirty_0_89; // @[d_cache.scala 24:26]
  reg  dirty_0_90; // @[d_cache.scala 24:26]
  reg  dirty_0_91; // @[d_cache.scala 24:26]
  reg  dirty_0_92; // @[d_cache.scala 24:26]
  reg  dirty_0_93; // @[d_cache.scala 24:26]
  reg  dirty_0_94; // @[d_cache.scala 24:26]
  reg  dirty_0_95; // @[d_cache.scala 24:26]
  reg  dirty_0_96; // @[d_cache.scala 24:26]
  reg  dirty_0_97; // @[d_cache.scala 24:26]
  reg  dirty_0_98; // @[d_cache.scala 24:26]
  reg  dirty_0_99; // @[d_cache.scala 24:26]
  reg  dirty_0_100; // @[d_cache.scala 24:26]
  reg  dirty_0_101; // @[d_cache.scala 24:26]
  reg  dirty_0_102; // @[d_cache.scala 24:26]
  reg  dirty_0_103; // @[d_cache.scala 24:26]
  reg  dirty_0_104; // @[d_cache.scala 24:26]
  reg  dirty_0_105; // @[d_cache.scala 24:26]
  reg  dirty_0_106; // @[d_cache.scala 24:26]
  reg  dirty_0_107; // @[d_cache.scala 24:26]
  reg  dirty_0_108; // @[d_cache.scala 24:26]
  reg  dirty_0_109; // @[d_cache.scala 24:26]
  reg  dirty_0_110; // @[d_cache.scala 24:26]
  reg  dirty_0_111; // @[d_cache.scala 24:26]
  reg  dirty_0_112; // @[d_cache.scala 24:26]
  reg  dirty_0_113; // @[d_cache.scala 24:26]
  reg  dirty_0_114; // @[d_cache.scala 24:26]
  reg  dirty_0_115; // @[d_cache.scala 24:26]
  reg  dirty_0_116; // @[d_cache.scala 24:26]
  reg  dirty_0_117; // @[d_cache.scala 24:26]
  reg  dirty_0_118; // @[d_cache.scala 24:26]
  reg  dirty_0_119; // @[d_cache.scala 24:26]
  reg  dirty_0_120; // @[d_cache.scala 24:26]
  reg  dirty_0_121; // @[d_cache.scala 24:26]
  reg  dirty_0_122; // @[d_cache.scala 24:26]
  reg  dirty_0_123; // @[d_cache.scala 24:26]
  reg  dirty_0_124; // @[d_cache.scala 24:26]
  reg  dirty_0_125; // @[d_cache.scala 24:26]
  reg  dirty_0_126; // @[d_cache.scala 24:26]
  reg  dirty_0_127; // @[d_cache.scala 24:26]
  reg  dirty_1_0; // @[d_cache.scala 25:26]
  reg  dirty_1_1; // @[d_cache.scala 25:26]
  reg  dirty_1_2; // @[d_cache.scala 25:26]
  reg  dirty_1_3; // @[d_cache.scala 25:26]
  reg  dirty_1_4; // @[d_cache.scala 25:26]
  reg  dirty_1_5; // @[d_cache.scala 25:26]
  reg  dirty_1_6; // @[d_cache.scala 25:26]
  reg  dirty_1_7; // @[d_cache.scala 25:26]
  reg  dirty_1_8; // @[d_cache.scala 25:26]
  reg  dirty_1_9; // @[d_cache.scala 25:26]
  reg  dirty_1_10; // @[d_cache.scala 25:26]
  reg  dirty_1_11; // @[d_cache.scala 25:26]
  reg  dirty_1_12; // @[d_cache.scala 25:26]
  reg  dirty_1_13; // @[d_cache.scala 25:26]
  reg  dirty_1_14; // @[d_cache.scala 25:26]
  reg  dirty_1_15; // @[d_cache.scala 25:26]
  reg  dirty_1_16; // @[d_cache.scala 25:26]
  reg  dirty_1_17; // @[d_cache.scala 25:26]
  reg  dirty_1_18; // @[d_cache.scala 25:26]
  reg  dirty_1_19; // @[d_cache.scala 25:26]
  reg  dirty_1_20; // @[d_cache.scala 25:26]
  reg  dirty_1_21; // @[d_cache.scala 25:26]
  reg  dirty_1_22; // @[d_cache.scala 25:26]
  reg  dirty_1_23; // @[d_cache.scala 25:26]
  reg  dirty_1_24; // @[d_cache.scala 25:26]
  reg  dirty_1_25; // @[d_cache.scala 25:26]
  reg  dirty_1_26; // @[d_cache.scala 25:26]
  reg  dirty_1_27; // @[d_cache.scala 25:26]
  reg  dirty_1_28; // @[d_cache.scala 25:26]
  reg  dirty_1_29; // @[d_cache.scala 25:26]
  reg  dirty_1_30; // @[d_cache.scala 25:26]
  reg  dirty_1_31; // @[d_cache.scala 25:26]
  reg  dirty_1_32; // @[d_cache.scala 25:26]
  reg  dirty_1_33; // @[d_cache.scala 25:26]
  reg  dirty_1_34; // @[d_cache.scala 25:26]
  reg  dirty_1_35; // @[d_cache.scala 25:26]
  reg  dirty_1_36; // @[d_cache.scala 25:26]
  reg  dirty_1_37; // @[d_cache.scala 25:26]
  reg  dirty_1_38; // @[d_cache.scala 25:26]
  reg  dirty_1_39; // @[d_cache.scala 25:26]
  reg  dirty_1_40; // @[d_cache.scala 25:26]
  reg  dirty_1_41; // @[d_cache.scala 25:26]
  reg  dirty_1_42; // @[d_cache.scala 25:26]
  reg  dirty_1_43; // @[d_cache.scala 25:26]
  reg  dirty_1_44; // @[d_cache.scala 25:26]
  reg  dirty_1_45; // @[d_cache.scala 25:26]
  reg  dirty_1_46; // @[d_cache.scala 25:26]
  reg  dirty_1_47; // @[d_cache.scala 25:26]
  reg  dirty_1_48; // @[d_cache.scala 25:26]
  reg  dirty_1_49; // @[d_cache.scala 25:26]
  reg  dirty_1_50; // @[d_cache.scala 25:26]
  reg  dirty_1_51; // @[d_cache.scala 25:26]
  reg  dirty_1_52; // @[d_cache.scala 25:26]
  reg  dirty_1_53; // @[d_cache.scala 25:26]
  reg  dirty_1_54; // @[d_cache.scala 25:26]
  reg  dirty_1_55; // @[d_cache.scala 25:26]
  reg  dirty_1_56; // @[d_cache.scala 25:26]
  reg  dirty_1_57; // @[d_cache.scala 25:26]
  reg  dirty_1_58; // @[d_cache.scala 25:26]
  reg  dirty_1_59; // @[d_cache.scala 25:26]
  reg  dirty_1_60; // @[d_cache.scala 25:26]
  reg  dirty_1_61; // @[d_cache.scala 25:26]
  reg  dirty_1_62; // @[d_cache.scala 25:26]
  reg  dirty_1_63; // @[d_cache.scala 25:26]
  reg  dirty_1_64; // @[d_cache.scala 25:26]
  reg  dirty_1_65; // @[d_cache.scala 25:26]
  reg  dirty_1_66; // @[d_cache.scala 25:26]
  reg  dirty_1_67; // @[d_cache.scala 25:26]
  reg  dirty_1_68; // @[d_cache.scala 25:26]
  reg  dirty_1_69; // @[d_cache.scala 25:26]
  reg  dirty_1_70; // @[d_cache.scala 25:26]
  reg  dirty_1_71; // @[d_cache.scala 25:26]
  reg  dirty_1_72; // @[d_cache.scala 25:26]
  reg  dirty_1_73; // @[d_cache.scala 25:26]
  reg  dirty_1_74; // @[d_cache.scala 25:26]
  reg  dirty_1_75; // @[d_cache.scala 25:26]
  reg  dirty_1_76; // @[d_cache.scala 25:26]
  reg  dirty_1_77; // @[d_cache.scala 25:26]
  reg  dirty_1_78; // @[d_cache.scala 25:26]
  reg  dirty_1_79; // @[d_cache.scala 25:26]
  reg  dirty_1_80; // @[d_cache.scala 25:26]
  reg  dirty_1_81; // @[d_cache.scala 25:26]
  reg  dirty_1_82; // @[d_cache.scala 25:26]
  reg  dirty_1_83; // @[d_cache.scala 25:26]
  reg  dirty_1_84; // @[d_cache.scala 25:26]
  reg  dirty_1_85; // @[d_cache.scala 25:26]
  reg  dirty_1_86; // @[d_cache.scala 25:26]
  reg  dirty_1_87; // @[d_cache.scala 25:26]
  reg  dirty_1_88; // @[d_cache.scala 25:26]
  reg  dirty_1_89; // @[d_cache.scala 25:26]
  reg  dirty_1_90; // @[d_cache.scala 25:26]
  reg  dirty_1_91; // @[d_cache.scala 25:26]
  reg  dirty_1_92; // @[d_cache.scala 25:26]
  reg  dirty_1_93; // @[d_cache.scala 25:26]
  reg  dirty_1_94; // @[d_cache.scala 25:26]
  reg  dirty_1_95; // @[d_cache.scala 25:26]
  reg  dirty_1_96; // @[d_cache.scala 25:26]
  reg  dirty_1_97; // @[d_cache.scala 25:26]
  reg  dirty_1_98; // @[d_cache.scala 25:26]
  reg  dirty_1_99; // @[d_cache.scala 25:26]
  reg  dirty_1_100; // @[d_cache.scala 25:26]
  reg  dirty_1_101; // @[d_cache.scala 25:26]
  reg  dirty_1_102; // @[d_cache.scala 25:26]
  reg  dirty_1_103; // @[d_cache.scala 25:26]
  reg  dirty_1_104; // @[d_cache.scala 25:26]
  reg  dirty_1_105; // @[d_cache.scala 25:26]
  reg  dirty_1_106; // @[d_cache.scala 25:26]
  reg  dirty_1_107; // @[d_cache.scala 25:26]
  reg  dirty_1_108; // @[d_cache.scala 25:26]
  reg  dirty_1_109; // @[d_cache.scala 25:26]
  reg  dirty_1_110; // @[d_cache.scala 25:26]
  reg  dirty_1_111; // @[d_cache.scala 25:26]
  reg  dirty_1_112; // @[d_cache.scala 25:26]
  reg  dirty_1_113; // @[d_cache.scala 25:26]
  reg  dirty_1_114; // @[d_cache.scala 25:26]
  reg  dirty_1_115; // @[d_cache.scala 25:26]
  reg  dirty_1_116; // @[d_cache.scala 25:26]
  reg  dirty_1_117; // @[d_cache.scala 25:26]
  reg  dirty_1_118; // @[d_cache.scala 25:26]
  reg  dirty_1_119; // @[d_cache.scala 25:26]
  reg  dirty_1_120; // @[d_cache.scala 25:26]
  reg  dirty_1_121; // @[d_cache.scala 25:26]
  reg  dirty_1_122; // @[d_cache.scala 25:26]
  reg  dirty_1_123; // @[d_cache.scala 25:26]
  reg  dirty_1_124; // @[d_cache.scala 25:26]
  reg  dirty_1_125; // @[d_cache.scala 25:26]
  reg  dirty_1_126; // @[d_cache.scala 25:26]
  reg  dirty_1_127; // @[d_cache.scala 25:26]
  reg  way0_hit; // @[d_cache.scala 26:27]
  reg  way1_hit; // @[d_cache.scala 27:27]
  reg [63:0] write_back_data; // @[d_cache.scala 29:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 30:34]
  reg [1:0] unuse_way; // @[d_cache.scala 33:28]
  reg [63:0] receive_data; // @[d_cache.scala 34:31]
  reg  quene; // @[d_cache.scala 35:24]
  wire [2:0] offset = io_from_lsu_araddr[2:0]; // @[d_cache.scala 37:36]
  wire [21:0] tag = io_from_lsu_araddr[31:10]; // @[d_cache.scala 39:33]
  wire [5:0] _shift_bit_T_8 = offset == 3'h7 ? 6'h38 : 6'h0; // @[d_cache.scala 47:24]
  wire [5:0] _shift_bit_T_9 = offset == 3'h6 ? 6'h30 : _shift_bit_T_8; // @[d_cache.scala 46:24]
  wire [5:0] _shift_bit_T_10 = offset == 3'h5 ? 6'h28 : _shift_bit_T_9; // @[d_cache.scala 45:24]
  wire [5:0] _shift_bit_T_11 = offset == 3'h4 ? 6'h20 : _shift_bit_T_10; // @[d_cache.scala 44:24]
  wire [5:0] _shift_bit_T_12 = offset == 3'h3 ? 6'h18 : _shift_bit_T_11; // @[d_cache.scala 43:24]
  wire [5:0] _shift_bit_T_13 = offset == 3'h2 ? 6'h10 : _shift_bit_T_12; // @[d_cache.scala 42:24]
  wire [5:0] _shift_bit_T_14 = offset == 3'h1 ? 6'h8 : _shift_bit_T_13; // @[d_cache.scala 41:24]
  wire [5:0] shift_bit = offset == 3'h0 ? 6'h0 : _shift_bit_T_14; // @[d_cache.scala 40:24]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 52:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 51:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 50:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 49:20]
  wire [31:0] index = {{25'd0}, io_from_lsu_araddr[9:3]}; // @[d_cache.scala 36:21 38:11]
  wire [31:0] _GEN_1 = 7'h1 == index[6:0] ? tag_0_1 : tag_0_0; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_2 = 7'h2 == index[6:0] ? tag_0_2 : _GEN_1; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_3 = 7'h3 == index[6:0] ? tag_0_3 : _GEN_2; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_4 = 7'h4 == index[6:0] ? tag_0_4 : _GEN_3; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_5 = 7'h5 == index[6:0] ? tag_0_5 : _GEN_4; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_6 = 7'h6 == index[6:0] ? tag_0_6 : _GEN_5; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_7 = 7'h7 == index[6:0] ? tag_0_7 : _GEN_6; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_8 = 7'h8 == index[6:0] ? tag_0_8 : _GEN_7; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_9 = 7'h9 == index[6:0] ? tag_0_9 : _GEN_8; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_10 = 7'ha == index[6:0] ? tag_0_10 : _GEN_9; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_11 = 7'hb == index[6:0] ? tag_0_11 : _GEN_10; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_12 = 7'hc == index[6:0] ? tag_0_12 : _GEN_11; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_13 = 7'hd == index[6:0] ? tag_0_13 : _GEN_12; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_14 = 7'he == index[6:0] ? tag_0_14 : _GEN_13; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_15 = 7'hf == index[6:0] ? tag_0_15 : _GEN_14; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_16 = 7'h10 == index[6:0] ? tag_0_16 : _GEN_15; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_17 = 7'h11 == index[6:0] ? tag_0_17 : _GEN_16; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_18 = 7'h12 == index[6:0] ? tag_0_18 : _GEN_17; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_19 = 7'h13 == index[6:0] ? tag_0_19 : _GEN_18; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_20 = 7'h14 == index[6:0] ? tag_0_20 : _GEN_19; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_21 = 7'h15 == index[6:0] ? tag_0_21 : _GEN_20; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_22 = 7'h16 == index[6:0] ? tag_0_22 : _GEN_21; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_23 = 7'h17 == index[6:0] ? tag_0_23 : _GEN_22; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_24 = 7'h18 == index[6:0] ? tag_0_24 : _GEN_23; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_25 = 7'h19 == index[6:0] ? tag_0_25 : _GEN_24; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_26 = 7'h1a == index[6:0] ? tag_0_26 : _GEN_25; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_27 = 7'h1b == index[6:0] ? tag_0_27 : _GEN_26; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_28 = 7'h1c == index[6:0] ? tag_0_28 : _GEN_27; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_29 = 7'h1d == index[6:0] ? tag_0_29 : _GEN_28; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_30 = 7'h1e == index[6:0] ? tag_0_30 : _GEN_29; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_31 = 7'h1f == index[6:0] ? tag_0_31 : _GEN_30; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_32 = 7'h20 == index[6:0] ? tag_0_32 : _GEN_31; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_33 = 7'h21 == index[6:0] ? tag_0_33 : _GEN_32; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_34 = 7'h22 == index[6:0] ? tag_0_34 : _GEN_33; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_35 = 7'h23 == index[6:0] ? tag_0_35 : _GEN_34; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_36 = 7'h24 == index[6:0] ? tag_0_36 : _GEN_35; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_37 = 7'h25 == index[6:0] ? tag_0_37 : _GEN_36; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_38 = 7'h26 == index[6:0] ? tag_0_38 : _GEN_37; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_39 = 7'h27 == index[6:0] ? tag_0_39 : _GEN_38; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_40 = 7'h28 == index[6:0] ? tag_0_40 : _GEN_39; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_41 = 7'h29 == index[6:0] ? tag_0_41 : _GEN_40; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_42 = 7'h2a == index[6:0] ? tag_0_42 : _GEN_41; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_43 = 7'h2b == index[6:0] ? tag_0_43 : _GEN_42; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_44 = 7'h2c == index[6:0] ? tag_0_44 : _GEN_43; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_45 = 7'h2d == index[6:0] ? tag_0_45 : _GEN_44; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_46 = 7'h2e == index[6:0] ? tag_0_46 : _GEN_45; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_47 = 7'h2f == index[6:0] ? tag_0_47 : _GEN_46; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_48 = 7'h30 == index[6:0] ? tag_0_48 : _GEN_47; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_49 = 7'h31 == index[6:0] ? tag_0_49 : _GEN_48; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_50 = 7'h32 == index[6:0] ? tag_0_50 : _GEN_49; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_51 = 7'h33 == index[6:0] ? tag_0_51 : _GEN_50; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_52 = 7'h34 == index[6:0] ? tag_0_52 : _GEN_51; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_53 = 7'h35 == index[6:0] ? tag_0_53 : _GEN_52; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_54 = 7'h36 == index[6:0] ? tag_0_54 : _GEN_53; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_55 = 7'h37 == index[6:0] ? tag_0_55 : _GEN_54; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_56 = 7'h38 == index[6:0] ? tag_0_56 : _GEN_55; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_57 = 7'h39 == index[6:0] ? tag_0_57 : _GEN_56; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_58 = 7'h3a == index[6:0] ? tag_0_58 : _GEN_57; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_59 = 7'h3b == index[6:0] ? tag_0_59 : _GEN_58; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_60 = 7'h3c == index[6:0] ? tag_0_60 : _GEN_59; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_61 = 7'h3d == index[6:0] ? tag_0_61 : _GEN_60; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_62 = 7'h3e == index[6:0] ? tag_0_62 : _GEN_61; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_63 = 7'h3f == index[6:0] ? tag_0_63 : _GEN_62; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_64 = 7'h40 == index[6:0] ? tag_0_64 : _GEN_63; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_65 = 7'h41 == index[6:0] ? tag_0_65 : _GEN_64; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_66 = 7'h42 == index[6:0] ? tag_0_66 : _GEN_65; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_67 = 7'h43 == index[6:0] ? tag_0_67 : _GEN_66; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_68 = 7'h44 == index[6:0] ? tag_0_68 : _GEN_67; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_69 = 7'h45 == index[6:0] ? tag_0_69 : _GEN_68; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_70 = 7'h46 == index[6:0] ? tag_0_70 : _GEN_69; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_71 = 7'h47 == index[6:0] ? tag_0_71 : _GEN_70; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_72 = 7'h48 == index[6:0] ? tag_0_72 : _GEN_71; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_73 = 7'h49 == index[6:0] ? tag_0_73 : _GEN_72; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_74 = 7'h4a == index[6:0] ? tag_0_74 : _GEN_73; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_75 = 7'h4b == index[6:0] ? tag_0_75 : _GEN_74; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_76 = 7'h4c == index[6:0] ? tag_0_76 : _GEN_75; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_77 = 7'h4d == index[6:0] ? tag_0_77 : _GEN_76; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_78 = 7'h4e == index[6:0] ? tag_0_78 : _GEN_77; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_79 = 7'h4f == index[6:0] ? tag_0_79 : _GEN_78; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_80 = 7'h50 == index[6:0] ? tag_0_80 : _GEN_79; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_81 = 7'h51 == index[6:0] ? tag_0_81 : _GEN_80; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_82 = 7'h52 == index[6:0] ? tag_0_82 : _GEN_81; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_83 = 7'h53 == index[6:0] ? tag_0_83 : _GEN_82; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_84 = 7'h54 == index[6:0] ? tag_0_84 : _GEN_83; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_85 = 7'h55 == index[6:0] ? tag_0_85 : _GEN_84; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_86 = 7'h56 == index[6:0] ? tag_0_86 : _GEN_85; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_87 = 7'h57 == index[6:0] ? tag_0_87 : _GEN_86; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_88 = 7'h58 == index[6:0] ? tag_0_88 : _GEN_87; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_89 = 7'h59 == index[6:0] ? tag_0_89 : _GEN_88; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_90 = 7'h5a == index[6:0] ? tag_0_90 : _GEN_89; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_91 = 7'h5b == index[6:0] ? tag_0_91 : _GEN_90; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_92 = 7'h5c == index[6:0] ? tag_0_92 : _GEN_91; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_93 = 7'h5d == index[6:0] ? tag_0_93 : _GEN_92; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_94 = 7'h5e == index[6:0] ? tag_0_94 : _GEN_93; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_95 = 7'h5f == index[6:0] ? tag_0_95 : _GEN_94; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_96 = 7'h60 == index[6:0] ? tag_0_96 : _GEN_95; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_97 = 7'h61 == index[6:0] ? tag_0_97 : _GEN_96; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_98 = 7'h62 == index[6:0] ? tag_0_98 : _GEN_97; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_99 = 7'h63 == index[6:0] ? tag_0_99 : _GEN_98; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_100 = 7'h64 == index[6:0] ? tag_0_100 : _GEN_99; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_101 = 7'h65 == index[6:0] ? tag_0_101 : _GEN_100; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_102 = 7'h66 == index[6:0] ? tag_0_102 : _GEN_101; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_103 = 7'h67 == index[6:0] ? tag_0_103 : _GEN_102; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_104 = 7'h68 == index[6:0] ? tag_0_104 : _GEN_103; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_105 = 7'h69 == index[6:0] ? tag_0_105 : _GEN_104; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_106 = 7'h6a == index[6:0] ? tag_0_106 : _GEN_105; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_107 = 7'h6b == index[6:0] ? tag_0_107 : _GEN_106; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_108 = 7'h6c == index[6:0] ? tag_0_108 : _GEN_107; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_109 = 7'h6d == index[6:0] ? tag_0_109 : _GEN_108; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_110 = 7'h6e == index[6:0] ? tag_0_110 : _GEN_109; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_111 = 7'h6f == index[6:0] ? tag_0_111 : _GEN_110; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_112 = 7'h70 == index[6:0] ? tag_0_112 : _GEN_111; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_113 = 7'h71 == index[6:0] ? tag_0_113 : _GEN_112; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_114 = 7'h72 == index[6:0] ? tag_0_114 : _GEN_113; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_115 = 7'h73 == index[6:0] ? tag_0_115 : _GEN_114; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_116 = 7'h74 == index[6:0] ? tag_0_116 : _GEN_115; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_117 = 7'h75 == index[6:0] ? tag_0_117 : _GEN_116; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_118 = 7'h76 == index[6:0] ? tag_0_118 : _GEN_117; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_119 = 7'h77 == index[6:0] ? tag_0_119 : _GEN_118; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_120 = 7'h78 == index[6:0] ? tag_0_120 : _GEN_119; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_121 = 7'h79 == index[6:0] ? tag_0_121 : _GEN_120; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_122 = 7'h7a == index[6:0] ? tag_0_122 : _GEN_121; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_123 = 7'h7b == index[6:0] ? tag_0_123 : _GEN_122; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_124 = 7'h7c == index[6:0] ? tag_0_124 : _GEN_123; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_125 = 7'h7d == index[6:0] ? tag_0_125 : _GEN_124; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_126 = 7'h7e == index[6:0] ? tag_0_126 : _GEN_125; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_127 = 7'h7f == index[6:0] ? tag_0_127 : _GEN_126; // @[d_cache.scala 54:{24,24}]
  wire [31:0] _GEN_16801 = {{10'd0}, tag}; // @[d_cache.scala 54:24]
  wire  _GEN_129 = 7'h1 == index[6:0] ? valid_0_1 : valid_0_0; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_130 = 7'h2 == index[6:0] ? valid_0_2 : _GEN_129; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_131 = 7'h3 == index[6:0] ? valid_0_3 : _GEN_130; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_132 = 7'h4 == index[6:0] ? valid_0_4 : _GEN_131; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_133 = 7'h5 == index[6:0] ? valid_0_5 : _GEN_132; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_134 = 7'h6 == index[6:0] ? valid_0_6 : _GEN_133; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_135 = 7'h7 == index[6:0] ? valid_0_7 : _GEN_134; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_136 = 7'h8 == index[6:0] ? valid_0_8 : _GEN_135; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_137 = 7'h9 == index[6:0] ? valid_0_9 : _GEN_136; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_138 = 7'ha == index[6:0] ? valid_0_10 : _GEN_137; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_139 = 7'hb == index[6:0] ? valid_0_11 : _GEN_138; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_140 = 7'hc == index[6:0] ? valid_0_12 : _GEN_139; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_141 = 7'hd == index[6:0] ? valid_0_13 : _GEN_140; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_142 = 7'he == index[6:0] ? valid_0_14 : _GEN_141; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_143 = 7'hf == index[6:0] ? valid_0_15 : _GEN_142; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_144 = 7'h10 == index[6:0] ? valid_0_16 : _GEN_143; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_145 = 7'h11 == index[6:0] ? valid_0_17 : _GEN_144; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_146 = 7'h12 == index[6:0] ? valid_0_18 : _GEN_145; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_147 = 7'h13 == index[6:0] ? valid_0_19 : _GEN_146; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_148 = 7'h14 == index[6:0] ? valid_0_20 : _GEN_147; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_149 = 7'h15 == index[6:0] ? valid_0_21 : _GEN_148; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_150 = 7'h16 == index[6:0] ? valid_0_22 : _GEN_149; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_151 = 7'h17 == index[6:0] ? valid_0_23 : _GEN_150; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_152 = 7'h18 == index[6:0] ? valid_0_24 : _GEN_151; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_153 = 7'h19 == index[6:0] ? valid_0_25 : _GEN_152; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_154 = 7'h1a == index[6:0] ? valid_0_26 : _GEN_153; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_155 = 7'h1b == index[6:0] ? valid_0_27 : _GEN_154; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_156 = 7'h1c == index[6:0] ? valid_0_28 : _GEN_155; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_157 = 7'h1d == index[6:0] ? valid_0_29 : _GEN_156; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_158 = 7'h1e == index[6:0] ? valid_0_30 : _GEN_157; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_159 = 7'h1f == index[6:0] ? valid_0_31 : _GEN_158; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_160 = 7'h20 == index[6:0] ? valid_0_32 : _GEN_159; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_161 = 7'h21 == index[6:0] ? valid_0_33 : _GEN_160; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_162 = 7'h22 == index[6:0] ? valid_0_34 : _GEN_161; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_163 = 7'h23 == index[6:0] ? valid_0_35 : _GEN_162; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_164 = 7'h24 == index[6:0] ? valid_0_36 : _GEN_163; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_165 = 7'h25 == index[6:0] ? valid_0_37 : _GEN_164; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_166 = 7'h26 == index[6:0] ? valid_0_38 : _GEN_165; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_167 = 7'h27 == index[6:0] ? valid_0_39 : _GEN_166; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_168 = 7'h28 == index[6:0] ? valid_0_40 : _GEN_167; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_169 = 7'h29 == index[6:0] ? valid_0_41 : _GEN_168; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_170 = 7'h2a == index[6:0] ? valid_0_42 : _GEN_169; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_171 = 7'h2b == index[6:0] ? valid_0_43 : _GEN_170; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_172 = 7'h2c == index[6:0] ? valid_0_44 : _GEN_171; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_173 = 7'h2d == index[6:0] ? valid_0_45 : _GEN_172; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_174 = 7'h2e == index[6:0] ? valid_0_46 : _GEN_173; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_175 = 7'h2f == index[6:0] ? valid_0_47 : _GEN_174; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_176 = 7'h30 == index[6:0] ? valid_0_48 : _GEN_175; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_177 = 7'h31 == index[6:0] ? valid_0_49 : _GEN_176; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_178 = 7'h32 == index[6:0] ? valid_0_50 : _GEN_177; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_179 = 7'h33 == index[6:0] ? valid_0_51 : _GEN_178; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_180 = 7'h34 == index[6:0] ? valid_0_52 : _GEN_179; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_181 = 7'h35 == index[6:0] ? valid_0_53 : _GEN_180; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_182 = 7'h36 == index[6:0] ? valid_0_54 : _GEN_181; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_183 = 7'h37 == index[6:0] ? valid_0_55 : _GEN_182; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_184 = 7'h38 == index[6:0] ? valid_0_56 : _GEN_183; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_185 = 7'h39 == index[6:0] ? valid_0_57 : _GEN_184; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_186 = 7'h3a == index[6:0] ? valid_0_58 : _GEN_185; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_187 = 7'h3b == index[6:0] ? valid_0_59 : _GEN_186; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_188 = 7'h3c == index[6:0] ? valid_0_60 : _GEN_187; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_189 = 7'h3d == index[6:0] ? valid_0_61 : _GEN_188; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_190 = 7'h3e == index[6:0] ? valid_0_62 : _GEN_189; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_191 = 7'h3f == index[6:0] ? valid_0_63 : _GEN_190; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_192 = 7'h40 == index[6:0] ? valid_0_64 : _GEN_191; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_193 = 7'h41 == index[6:0] ? valid_0_65 : _GEN_192; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_194 = 7'h42 == index[6:0] ? valid_0_66 : _GEN_193; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_195 = 7'h43 == index[6:0] ? valid_0_67 : _GEN_194; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_196 = 7'h44 == index[6:0] ? valid_0_68 : _GEN_195; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_197 = 7'h45 == index[6:0] ? valid_0_69 : _GEN_196; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_198 = 7'h46 == index[6:0] ? valid_0_70 : _GEN_197; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_199 = 7'h47 == index[6:0] ? valid_0_71 : _GEN_198; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_200 = 7'h48 == index[6:0] ? valid_0_72 : _GEN_199; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_201 = 7'h49 == index[6:0] ? valid_0_73 : _GEN_200; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_202 = 7'h4a == index[6:0] ? valid_0_74 : _GEN_201; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_203 = 7'h4b == index[6:0] ? valid_0_75 : _GEN_202; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_204 = 7'h4c == index[6:0] ? valid_0_76 : _GEN_203; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_205 = 7'h4d == index[6:0] ? valid_0_77 : _GEN_204; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_206 = 7'h4e == index[6:0] ? valid_0_78 : _GEN_205; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_207 = 7'h4f == index[6:0] ? valid_0_79 : _GEN_206; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_208 = 7'h50 == index[6:0] ? valid_0_80 : _GEN_207; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_209 = 7'h51 == index[6:0] ? valid_0_81 : _GEN_208; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_210 = 7'h52 == index[6:0] ? valid_0_82 : _GEN_209; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_211 = 7'h53 == index[6:0] ? valid_0_83 : _GEN_210; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_212 = 7'h54 == index[6:0] ? valid_0_84 : _GEN_211; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_213 = 7'h55 == index[6:0] ? valid_0_85 : _GEN_212; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_214 = 7'h56 == index[6:0] ? valid_0_86 : _GEN_213; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_215 = 7'h57 == index[6:0] ? valid_0_87 : _GEN_214; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_216 = 7'h58 == index[6:0] ? valid_0_88 : _GEN_215; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_217 = 7'h59 == index[6:0] ? valid_0_89 : _GEN_216; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_218 = 7'h5a == index[6:0] ? valid_0_90 : _GEN_217; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_219 = 7'h5b == index[6:0] ? valid_0_91 : _GEN_218; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_220 = 7'h5c == index[6:0] ? valid_0_92 : _GEN_219; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_221 = 7'h5d == index[6:0] ? valid_0_93 : _GEN_220; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_222 = 7'h5e == index[6:0] ? valid_0_94 : _GEN_221; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_223 = 7'h5f == index[6:0] ? valid_0_95 : _GEN_222; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_224 = 7'h60 == index[6:0] ? valid_0_96 : _GEN_223; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_225 = 7'h61 == index[6:0] ? valid_0_97 : _GEN_224; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_226 = 7'h62 == index[6:0] ? valid_0_98 : _GEN_225; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_227 = 7'h63 == index[6:0] ? valid_0_99 : _GEN_226; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_228 = 7'h64 == index[6:0] ? valid_0_100 : _GEN_227; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_229 = 7'h65 == index[6:0] ? valid_0_101 : _GEN_228; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_230 = 7'h66 == index[6:0] ? valid_0_102 : _GEN_229; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_231 = 7'h67 == index[6:0] ? valid_0_103 : _GEN_230; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_232 = 7'h68 == index[6:0] ? valid_0_104 : _GEN_231; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_233 = 7'h69 == index[6:0] ? valid_0_105 : _GEN_232; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_234 = 7'h6a == index[6:0] ? valid_0_106 : _GEN_233; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_235 = 7'h6b == index[6:0] ? valid_0_107 : _GEN_234; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_236 = 7'h6c == index[6:0] ? valid_0_108 : _GEN_235; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_237 = 7'h6d == index[6:0] ? valid_0_109 : _GEN_236; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_238 = 7'h6e == index[6:0] ? valid_0_110 : _GEN_237; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_239 = 7'h6f == index[6:0] ? valid_0_111 : _GEN_238; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_240 = 7'h70 == index[6:0] ? valid_0_112 : _GEN_239; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_241 = 7'h71 == index[6:0] ? valid_0_113 : _GEN_240; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_242 = 7'h72 == index[6:0] ? valid_0_114 : _GEN_241; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_243 = 7'h73 == index[6:0] ? valid_0_115 : _GEN_242; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_244 = 7'h74 == index[6:0] ? valid_0_116 : _GEN_243; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_245 = 7'h75 == index[6:0] ? valid_0_117 : _GEN_244; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_246 = 7'h76 == index[6:0] ? valid_0_118 : _GEN_245; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_247 = 7'h77 == index[6:0] ? valid_0_119 : _GEN_246; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_248 = 7'h78 == index[6:0] ? valid_0_120 : _GEN_247; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_249 = 7'h79 == index[6:0] ? valid_0_121 : _GEN_248; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_250 = 7'h7a == index[6:0] ? valid_0_122 : _GEN_249; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_251 = 7'h7b == index[6:0] ? valid_0_123 : _GEN_250; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_252 = 7'h7c == index[6:0] ? valid_0_124 : _GEN_251; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_253 = 7'h7d == index[6:0] ? valid_0_125 : _GEN_252; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_254 = 7'h7e == index[6:0] ? valid_0_126 : _GEN_253; // @[d_cache.scala 54:{50,50}]
  wire  _GEN_255 = 7'h7f == index[6:0] ? valid_0_127 : _GEN_254; // @[d_cache.scala 54:{50,50}]
  wire  _T_6 = _GEN_127 == _GEN_16801 & _GEN_255; // @[d_cache.scala 54:33]
  wire [31:0] _GEN_258 = 7'h1 == index[6:0] ? tag_1_1 : tag_1_0; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_259 = 7'h2 == index[6:0] ? tag_1_2 : _GEN_258; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_260 = 7'h3 == index[6:0] ? tag_1_3 : _GEN_259; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_261 = 7'h4 == index[6:0] ? tag_1_4 : _GEN_260; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_262 = 7'h5 == index[6:0] ? tag_1_5 : _GEN_261; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_263 = 7'h6 == index[6:0] ? tag_1_6 : _GEN_262; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_264 = 7'h7 == index[6:0] ? tag_1_7 : _GEN_263; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_265 = 7'h8 == index[6:0] ? tag_1_8 : _GEN_264; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_266 = 7'h9 == index[6:0] ? tag_1_9 : _GEN_265; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_267 = 7'ha == index[6:0] ? tag_1_10 : _GEN_266; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_268 = 7'hb == index[6:0] ? tag_1_11 : _GEN_267; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_269 = 7'hc == index[6:0] ? tag_1_12 : _GEN_268; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_270 = 7'hd == index[6:0] ? tag_1_13 : _GEN_269; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_271 = 7'he == index[6:0] ? tag_1_14 : _GEN_270; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_272 = 7'hf == index[6:0] ? tag_1_15 : _GEN_271; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_273 = 7'h10 == index[6:0] ? tag_1_16 : _GEN_272; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_274 = 7'h11 == index[6:0] ? tag_1_17 : _GEN_273; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_275 = 7'h12 == index[6:0] ? tag_1_18 : _GEN_274; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_276 = 7'h13 == index[6:0] ? tag_1_19 : _GEN_275; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_277 = 7'h14 == index[6:0] ? tag_1_20 : _GEN_276; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_278 = 7'h15 == index[6:0] ? tag_1_21 : _GEN_277; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_279 = 7'h16 == index[6:0] ? tag_1_22 : _GEN_278; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_280 = 7'h17 == index[6:0] ? tag_1_23 : _GEN_279; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_281 = 7'h18 == index[6:0] ? tag_1_24 : _GEN_280; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_282 = 7'h19 == index[6:0] ? tag_1_25 : _GEN_281; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_283 = 7'h1a == index[6:0] ? tag_1_26 : _GEN_282; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_284 = 7'h1b == index[6:0] ? tag_1_27 : _GEN_283; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_285 = 7'h1c == index[6:0] ? tag_1_28 : _GEN_284; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_286 = 7'h1d == index[6:0] ? tag_1_29 : _GEN_285; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_287 = 7'h1e == index[6:0] ? tag_1_30 : _GEN_286; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_288 = 7'h1f == index[6:0] ? tag_1_31 : _GEN_287; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_289 = 7'h20 == index[6:0] ? tag_1_32 : _GEN_288; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_290 = 7'h21 == index[6:0] ? tag_1_33 : _GEN_289; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_291 = 7'h22 == index[6:0] ? tag_1_34 : _GEN_290; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_292 = 7'h23 == index[6:0] ? tag_1_35 : _GEN_291; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_293 = 7'h24 == index[6:0] ? tag_1_36 : _GEN_292; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_294 = 7'h25 == index[6:0] ? tag_1_37 : _GEN_293; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_295 = 7'h26 == index[6:0] ? tag_1_38 : _GEN_294; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_296 = 7'h27 == index[6:0] ? tag_1_39 : _GEN_295; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_297 = 7'h28 == index[6:0] ? tag_1_40 : _GEN_296; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_298 = 7'h29 == index[6:0] ? tag_1_41 : _GEN_297; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_299 = 7'h2a == index[6:0] ? tag_1_42 : _GEN_298; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_300 = 7'h2b == index[6:0] ? tag_1_43 : _GEN_299; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_301 = 7'h2c == index[6:0] ? tag_1_44 : _GEN_300; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_302 = 7'h2d == index[6:0] ? tag_1_45 : _GEN_301; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_303 = 7'h2e == index[6:0] ? tag_1_46 : _GEN_302; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_304 = 7'h2f == index[6:0] ? tag_1_47 : _GEN_303; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_305 = 7'h30 == index[6:0] ? tag_1_48 : _GEN_304; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_306 = 7'h31 == index[6:0] ? tag_1_49 : _GEN_305; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_307 = 7'h32 == index[6:0] ? tag_1_50 : _GEN_306; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_308 = 7'h33 == index[6:0] ? tag_1_51 : _GEN_307; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_309 = 7'h34 == index[6:0] ? tag_1_52 : _GEN_308; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_310 = 7'h35 == index[6:0] ? tag_1_53 : _GEN_309; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_311 = 7'h36 == index[6:0] ? tag_1_54 : _GEN_310; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_312 = 7'h37 == index[6:0] ? tag_1_55 : _GEN_311; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_313 = 7'h38 == index[6:0] ? tag_1_56 : _GEN_312; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_314 = 7'h39 == index[6:0] ? tag_1_57 : _GEN_313; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_315 = 7'h3a == index[6:0] ? tag_1_58 : _GEN_314; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_316 = 7'h3b == index[6:0] ? tag_1_59 : _GEN_315; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_317 = 7'h3c == index[6:0] ? tag_1_60 : _GEN_316; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_318 = 7'h3d == index[6:0] ? tag_1_61 : _GEN_317; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_319 = 7'h3e == index[6:0] ? tag_1_62 : _GEN_318; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_320 = 7'h3f == index[6:0] ? tag_1_63 : _GEN_319; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_321 = 7'h40 == index[6:0] ? tag_1_64 : _GEN_320; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_322 = 7'h41 == index[6:0] ? tag_1_65 : _GEN_321; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_323 = 7'h42 == index[6:0] ? tag_1_66 : _GEN_322; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_324 = 7'h43 == index[6:0] ? tag_1_67 : _GEN_323; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_325 = 7'h44 == index[6:0] ? tag_1_68 : _GEN_324; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_326 = 7'h45 == index[6:0] ? tag_1_69 : _GEN_325; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_327 = 7'h46 == index[6:0] ? tag_1_70 : _GEN_326; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_328 = 7'h47 == index[6:0] ? tag_1_71 : _GEN_327; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_329 = 7'h48 == index[6:0] ? tag_1_72 : _GEN_328; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_330 = 7'h49 == index[6:0] ? tag_1_73 : _GEN_329; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_331 = 7'h4a == index[6:0] ? tag_1_74 : _GEN_330; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_332 = 7'h4b == index[6:0] ? tag_1_75 : _GEN_331; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_333 = 7'h4c == index[6:0] ? tag_1_76 : _GEN_332; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_334 = 7'h4d == index[6:0] ? tag_1_77 : _GEN_333; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_335 = 7'h4e == index[6:0] ? tag_1_78 : _GEN_334; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_336 = 7'h4f == index[6:0] ? tag_1_79 : _GEN_335; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_337 = 7'h50 == index[6:0] ? tag_1_80 : _GEN_336; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_338 = 7'h51 == index[6:0] ? tag_1_81 : _GEN_337; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_339 = 7'h52 == index[6:0] ? tag_1_82 : _GEN_338; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_340 = 7'h53 == index[6:0] ? tag_1_83 : _GEN_339; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_341 = 7'h54 == index[6:0] ? tag_1_84 : _GEN_340; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_342 = 7'h55 == index[6:0] ? tag_1_85 : _GEN_341; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_343 = 7'h56 == index[6:0] ? tag_1_86 : _GEN_342; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_344 = 7'h57 == index[6:0] ? tag_1_87 : _GEN_343; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_345 = 7'h58 == index[6:0] ? tag_1_88 : _GEN_344; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_346 = 7'h59 == index[6:0] ? tag_1_89 : _GEN_345; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_347 = 7'h5a == index[6:0] ? tag_1_90 : _GEN_346; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_348 = 7'h5b == index[6:0] ? tag_1_91 : _GEN_347; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_349 = 7'h5c == index[6:0] ? tag_1_92 : _GEN_348; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_350 = 7'h5d == index[6:0] ? tag_1_93 : _GEN_349; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_351 = 7'h5e == index[6:0] ? tag_1_94 : _GEN_350; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_352 = 7'h5f == index[6:0] ? tag_1_95 : _GEN_351; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_353 = 7'h60 == index[6:0] ? tag_1_96 : _GEN_352; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_354 = 7'h61 == index[6:0] ? tag_1_97 : _GEN_353; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_355 = 7'h62 == index[6:0] ? tag_1_98 : _GEN_354; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_356 = 7'h63 == index[6:0] ? tag_1_99 : _GEN_355; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_357 = 7'h64 == index[6:0] ? tag_1_100 : _GEN_356; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_358 = 7'h65 == index[6:0] ? tag_1_101 : _GEN_357; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_359 = 7'h66 == index[6:0] ? tag_1_102 : _GEN_358; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_360 = 7'h67 == index[6:0] ? tag_1_103 : _GEN_359; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_361 = 7'h68 == index[6:0] ? tag_1_104 : _GEN_360; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_362 = 7'h69 == index[6:0] ? tag_1_105 : _GEN_361; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_363 = 7'h6a == index[6:0] ? tag_1_106 : _GEN_362; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_364 = 7'h6b == index[6:0] ? tag_1_107 : _GEN_363; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_365 = 7'h6c == index[6:0] ? tag_1_108 : _GEN_364; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_366 = 7'h6d == index[6:0] ? tag_1_109 : _GEN_365; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_367 = 7'h6e == index[6:0] ? tag_1_110 : _GEN_366; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_368 = 7'h6f == index[6:0] ? tag_1_111 : _GEN_367; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_369 = 7'h70 == index[6:0] ? tag_1_112 : _GEN_368; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_370 = 7'h71 == index[6:0] ? tag_1_113 : _GEN_369; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_371 = 7'h72 == index[6:0] ? tag_1_114 : _GEN_370; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_372 = 7'h73 == index[6:0] ? tag_1_115 : _GEN_371; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_373 = 7'h74 == index[6:0] ? tag_1_116 : _GEN_372; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_374 = 7'h75 == index[6:0] ? tag_1_117 : _GEN_373; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_375 = 7'h76 == index[6:0] ? tag_1_118 : _GEN_374; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_376 = 7'h77 == index[6:0] ? tag_1_119 : _GEN_375; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_377 = 7'h78 == index[6:0] ? tag_1_120 : _GEN_376; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_378 = 7'h79 == index[6:0] ? tag_1_121 : _GEN_377; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_379 = 7'h7a == index[6:0] ? tag_1_122 : _GEN_378; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_380 = 7'h7b == index[6:0] ? tag_1_123 : _GEN_379; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_381 = 7'h7c == index[6:0] ? tag_1_124 : _GEN_380; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_382 = 7'h7d == index[6:0] ? tag_1_125 : _GEN_381; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_383 = 7'h7e == index[6:0] ? tag_1_126 : _GEN_382; // @[d_cache.scala 59:{24,24}]
  wire [31:0] _GEN_384 = 7'h7f == index[6:0] ? tag_1_127 : _GEN_383; // @[d_cache.scala 59:{24,24}]
  wire  _GEN_386 = 7'h1 == index[6:0] ? valid_1_1 : valid_1_0; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_387 = 7'h2 == index[6:0] ? valid_1_2 : _GEN_386; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_388 = 7'h3 == index[6:0] ? valid_1_3 : _GEN_387; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_389 = 7'h4 == index[6:0] ? valid_1_4 : _GEN_388; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_390 = 7'h5 == index[6:0] ? valid_1_5 : _GEN_389; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_391 = 7'h6 == index[6:0] ? valid_1_6 : _GEN_390; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_392 = 7'h7 == index[6:0] ? valid_1_7 : _GEN_391; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_393 = 7'h8 == index[6:0] ? valid_1_8 : _GEN_392; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_394 = 7'h9 == index[6:0] ? valid_1_9 : _GEN_393; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_395 = 7'ha == index[6:0] ? valid_1_10 : _GEN_394; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_396 = 7'hb == index[6:0] ? valid_1_11 : _GEN_395; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_397 = 7'hc == index[6:0] ? valid_1_12 : _GEN_396; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_398 = 7'hd == index[6:0] ? valid_1_13 : _GEN_397; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_399 = 7'he == index[6:0] ? valid_1_14 : _GEN_398; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_400 = 7'hf == index[6:0] ? valid_1_15 : _GEN_399; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_401 = 7'h10 == index[6:0] ? valid_1_16 : _GEN_400; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_402 = 7'h11 == index[6:0] ? valid_1_17 : _GEN_401; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_403 = 7'h12 == index[6:0] ? valid_1_18 : _GEN_402; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_404 = 7'h13 == index[6:0] ? valid_1_19 : _GEN_403; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_405 = 7'h14 == index[6:0] ? valid_1_20 : _GEN_404; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_406 = 7'h15 == index[6:0] ? valid_1_21 : _GEN_405; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_407 = 7'h16 == index[6:0] ? valid_1_22 : _GEN_406; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_408 = 7'h17 == index[6:0] ? valid_1_23 : _GEN_407; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_409 = 7'h18 == index[6:0] ? valid_1_24 : _GEN_408; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_410 = 7'h19 == index[6:0] ? valid_1_25 : _GEN_409; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_411 = 7'h1a == index[6:0] ? valid_1_26 : _GEN_410; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_412 = 7'h1b == index[6:0] ? valid_1_27 : _GEN_411; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_413 = 7'h1c == index[6:0] ? valid_1_28 : _GEN_412; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_414 = 7'h1d == index[6:0] ? valid_1_29 : _GEN_413; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_415 = 7'h1e == index[6:0] ? valid_1_30 : _GEN_414; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_416 = 7'h1f == index[6:0] ? valid_1_31 : _GEN_415; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_417 = 7'h20 == index[6:0] ? valid_1_32 : _GEN_416; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_418 = 7'h21 == index[6:0] ? valid_1_33 : _GEN_417; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_419 = 7'h22 == index[6:0] ? valid_1_34 : _GEN_418; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_420 = 7'h23 == index[6:0] ? valid_1_35 : _GEN_419; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_421 = 7'h24 == index[6:0] ? valid_1_36 : _GEN_420; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_422 = 7'h25 == index[6:0] ? valid_1_37 : _GEN_421; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_423 = 7'h26 == index[6:0] ? valid_1_38 : _GEN_422; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_424 = 7'h27 == index[6:0] ? valid_1_39 : _GEN_423; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_425 = 7'h28 == index[6:0] ? valid_1_40 : _GEN_424; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_426 = 7'h29 == index[6:0] ? valid_1_41 : _GEN_425; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_427 = 7'h2a == index[6:0] ? valid_1_42 : _GEN_426; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_428 = 7'h2b == index[6:0] ? valid_1_43 : _GEN_427; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_429 = 7'h2c == index[6:0] ? valid_1_44 : _GEN_428; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_430 = 7'h2d == index[6:0] ? valid_1_45 : _GEN_429; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_431 = 7'h2e == index[6:0] ? valid_1_46 : _GEN_430; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_432 = 7'h2f == index[6:0] ? valid_1_47 : _GEN_431; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_433 = 7'h30 == index[6:0] ? valid_1_48 : _GEN_432; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_434 = 7'h31 == index[6:0] ? valid_1_49 : _GEN_433; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_435 = 7'h32 == index[6:0] ? valid_1_50 : _GEN_434; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_436 = 7'h33 == index[6:0] ? valid_1_51 : _GEN_435; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_437 = 7'h34 == index[6:0] ? valid_1_52 : _GEN_436; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_438 = 7'h35 == index[6:0] ? valid_1_53 : _GEN_437; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_439 = 7'h36 == index[6:0] ? valid_1_54 : _GEN_438; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_440 = 7'h37 == index[6:0] ? valid_1_55 : _GEN_439; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_441 = 7'h38 == index[6:0] ? valid_1_56 : _GEN_440; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_442 = 7'h39 == index[6:0] ? valid_1_57 : _GEN_441; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_443 = 7'h3a == index[6:0] ? valid_1_58 : _GEN_442; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_444 = 7'h3b == index[6:0] ? valid_1_59 : _GEN_443; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_445 = 7'h3c == index[6:0] ? valid_1_60 : _GEN_444; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_446 = 7'h3d == index[6:0] ? valid_1_61 : _GEN_445; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_447 = 7'h3e == index[6:0] ? valid_1_62 : _GEN_446; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_448 = 7'h3f == index[6:0] ? valid_1_63 : _GEN_447; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_449 = 7'h40 == index[6:0] ? valid_1_64 : _GEN_448; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_450 = 7'h41 == index[6:0] ? valid_1_65 : _GEN_449; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_451 = 7'h42 == index[6:0] ? valid_1_66 : _GEN_450; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_452 = 7'h43 == index[6:0] ? valid_1_67 : _GEN_451; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_453 = 7'h44 == index[6:0] ? valid_1_68 : _GEN_452; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_454 = 7'h45 == index[6:0] ? valid_1_69 : _GEN_453; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_455 = 7'h46 == index[6:0] ? valid_1_70 : _GEN_454; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_456 = 7'h47 == index[6:0] ? valid_1_71 : _GEN_455; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_457 = 7'h48 == index[6:0] ? valid_1_72 : _GEN_456; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_458 = 7'h49 == index[6:0] ? valid_1_73 : _GEN_457; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_459 = 7'h4a == index[6:0] ? valid_1_74 : _GEN_458; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_460 = 7'h4b == index[6:0] ? valid_1_75 : _GEN_459; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_461 = 7'h4c == index[6:0] ? valid_1_76 : _GEN_460; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_462 = 7'h4d == index[6:0] ? valid_1_77 : _GEN_461; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_463 = 7'h4e == index[6:0] ? valid_1_78 : _GEN_462; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_464 = 7'h4f == index[6:0] ? valid_1_79 : _GEN_463; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_465 = 7'h50 == index[6:0] ? valid_1_80 : _GEN_464; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_466 = 7'h51 == index[6:0] ? valid_1_81 : _GEN_465; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_467 = 7'h52 == index[6:0] ? valid_1_82 : _GEN_466; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_468 = 7'h53 == index[6:0] ? valid_1_83 : _GEN_467; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_469 = 7'h54 == index[6:0] ? valid_1_84 : _GEN_468; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_470 = 7'h55 == index[6:0] ? valid_1_85 : _GEN_469; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_471 = 7'h56 == index[6:0] ? valid_1_86 : _GEN_470; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_472 = 7'h57 == index[6:0] ? valid_1_87 : _GEN_471; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_473 = 7'h58 == index[6:0] ? valid_1_88 : _GEN_472; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_474 = 7'h59 == index[6:0] ? valid_1_89 : _GEN_473; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_475 = 7'h5a == index[6:0] ? valid_1_90 : _GEN_474; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_476 = 7'h5b == index[6:0] ? valid_1_91 : _GEN_475; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_477 = 7'h5c == index[6:0] ? valid_1_92 : _GEN_476; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_478 = 7'h5d == index[6:0] ? valid_1_93 : _GEN_477; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_479 = 7'h5e == index[6:0] ? valid_1_94 : _GEN_478; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_480 = 7'h5f == index[6:0] ? valid_1_95 : _GEN_479; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_481 = 7'h60 == index[6:0] ? valid_1_96 : _GEN_480; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_482 = 7'h61 == index[6:0] ? valid_1_97 : _GEN_481; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_483 = 7'h62 == index[6:0] ? valid_1_98 : _GEN_482; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_484 = 7'h63 == index[6:0] ? valid_1_99 : _GEN_483; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_485 = 7'h64 == index[6:0] ? valid_1_100 : _GEN_484; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_486 = 7'h65 == index[6:0] ? valid_1_101 : _GEN_485; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_487 = 7'h66 == index[6:0] ? valid_1_102 : _GEN_486; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_488 = 7'h67 == index[6:0] ? valid_1_103 : _GEN_487; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_489 = 7'h68 == index[6:0] ? valid_1_104 : _GEN_488; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_490 = 7'h69 == index[6:0] ? valid_1_105 : _GEN_489; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_491 = 7'h6a == index[6:0] ? valid_1_106 : _GEN_490; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_492 = 7'h6b == index[6:0] ? valid_1_107 : _GEN_491; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_493 = 7'h6c == index[6:0] ? valid_1_108 : _GEN_492; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_494 = 7'h6d == index[6:0] ? valid_1_109 : _GEN_493; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_495 = 7'h6e == index[6:0] ? valid_1_110 : _GEN_494; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_496 = 7'h6f == index[6:0] ? valid_1_111 : _GEN_495; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_497 = 7'h70 == index[6:0] ? valid_1_112 : _GEN_496; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_498 = 7'h71 == index[6:0] ? valid_1_113 : _GEN_497; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_499 = 7'h72 == index[6:0] ? valid_1_114 : _GEN_498; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_500 = 7'h73 == index[6:0] ? valid_1_115 : _GEN_499; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_501 = 7'h74 == index[6:0] ? valid_1_116 : _GEN_500; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_502 = 7'h75 == index[6:0] ? valid_1_117 : _GEN_501; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_503 = 7'h76 == index[6:0] ? valid_1_118 : _GEN_502; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_504 = 7'h77 == index[6:0] ? valid_1_119 : _GEN_503; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_505 = 7'h78 == index[6:0] ? valid_1_120 : _GEN_504; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_506 = 7'h79 == index[6:0] ? valid_1_121 : _GEN_505; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_507 = 7'h7a == index[6:0] ? valid_1_122 : _GEN_506; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_508 = 7'h7b == index[6:0] ? valid_1_123 : _GEN_507; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_509 = 7'h7c == index[6:0] ? valid_1_124 : _GEN_508; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_510 = 7'h7d == index[6:0] ? valid_1_125 : _GEN_509; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_511 = 7'h7e == index[6:0] ? valid_1_126 : _GEN_510; // @[d_cache.scala 59:{50,50}]
  wire  _GEN_512 = 7'h7f == index[6:0] ? valid_1_127 : _GEN_511; // @[d_cache.scala 59:{50,50}]
  wire  _T_11 = _GEN_384 == _GEN_16801 & _GEN_512; // @[d_cache.scala 59:33]
  reg [2:0] state; // @[d_cache.scala 73:24]
  wire  _T_24 = 3'h0 == state; // @[d_cache.scala 78:18]
  wire  _T_25 = 3'h1 == state; // @[d_cache.scala 78:18]
  wire  _GEN_775 = 7'h1 == index[6:0] ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_776 = 7'h2 == index[6:0] ? dirty_0_2 : _GEN_775; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_777 = 7'h3 == index[6:0] ? dirty_0_3 : _GEN_776; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_778 = 7'h4 == index[6:0] ? dirty_0_4 : _GEN_777; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_779 = 7'h5 == index[6:0] ? dirty_0_5 : _GEN_778; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_780 = 7'h6 == index[6:0] ? dirty_0_6 : _GEN_779; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_781 = 7'h7 == index[6:0] ? dirty_0_7 : _GEN_780; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_782 = 7'h8 == index[6:0] ? dirty_0_8 : _GEN_781; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_783 = 7'h9 == index[6:0] ? dirty_0_9 : _GEN_782; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_784 = 7'ha == index[6:0] ? dirty_0_10 : _GEN_783; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_785 = 7'hb == index[6:0] ? dirty_0_11 : _GEN_784; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_786 = 7'hc == index[6:0] ? dirty_0_12 : _GEN_785; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_787 = 7'hd == index[6:0] ? dirty_0_13 : _GEN_786; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_788 = 7'he == index[6:0] ? dirty_0_14 : _GEN_787; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_789 = 7'hf == index[6:0] ? dirty_0_15 : _GEN_788; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_790 = 7'h10 == index[6:0] ? dirty_0_16 : _GEN_789; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_791 = 7'h11 == index[6:0] ? dirty_0_17 : _GEN_790; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_792 = 7'h12 == index[6:0] ? dirty_0_18 : _GEN_791; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_793 = 7'h13 == index[6:0] ? dirty_0_19 : _GEN_792; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_794 = 7'h14 == index[6:0] ? dirty_0_20 : _GEN_793; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_795 = 7'h15 == index[6:0] ? dirty_0_21 : _GEN_794; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_796 = 7'h16 == index[6:0] ? dirty_0_22 : _GEN_795; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_797 = 7'h17 == index[6:0] ? dirty_0_23 : _GEN_796; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_798 = 7'h18 == index[6:0] ? dirty_0_24 : _GEN_797; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_799 = 7'h19 == index[6:0] ? dirty_0_25 : _GEN_798; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_800 = 7'h1a == index[6:0] ? dirty_0_26 : _GEN_799; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_801 = 7'h1b == index[6:0] ? dirty_0_27 : _GEN_800; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_802 = 7'h1c == index[6:0] ? dirty_0_28 : _GEN_801; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_803 = 7'h1d == index[6:0] ? dirty_0_29 : _GEN_802; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_804 = 7'h1e == index[6:0] ? dirty_0_30 : _GEN_803; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_805 = 7'h1f == index[6:0] ? dirty_0_31 : _GEN_804; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_806 = 7'h20 == index[6:0] ? dirty_0_32 : _GEN_805; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_807 = 7'h21 == index[6:0] ? dirty_0_33 : _GEN_806; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_808 = 7'h22 == index[6:0] ? dirty_0_34 : _GEN_807; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_809 = 7'h23 == index[6:0] ? dirty_0_35 : _GEN_808; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_810 = 7'h24 == index[6:0] ? dirty_0_36 : _GEN_809; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_811 = 7'h25 == index[6:0] ? dirty_0_37 : _GEN_810; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_812 = 7'h26 == index[6:0] ? dirty_0_38 : _GEN_811; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_813 = 7'h27 == index[6:0] ? dirty_0_39 : _GEN_812; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_814 = 7'h28 == index[6:0] ? dirty_0_40 : _GEN_813; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_815 = 7'h29 == index[6:0] ? dirty_0_41 : _GEN_814; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_816 = 7'h2a == index[6:0] ? dirty_0_42 : _GEN_815; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_817 = 7'h2b == index[6:0] ? dirty_0_43 : _GEN_816; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_818 = 7'h2c == index[6:0] ? dirty_0_44 : _GEN_817; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_819 = 7'h2d == index[6:0] ? dirty_0_45 : _GEN_818; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_820 = 7'h2e == index[6:0] ? dirty_0_46 : _GEN_819; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_821 = 7'h2f == index[6:0] ? dirty_0_47 : _GEN_820; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_822 = 7'h30 == index[6:0] ? dirty_0_48 : _GEN_821; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_823 = 7'h31 == index[6:0] ? dirty_0_49 : _GEN_822; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_824 = 7'h32 == index[6:0] ? dirty_0_50 : _GEN_823; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_825 = 7'h33 == index[6:0] ? dirty_0_51 : _GEN_824; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_826 = 7'h34 == index[6:0] ? dirty_0_52 : _GEN_825; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_827 = 7'h35 == index[6:0] ? dirty_0_53 : _GEN_826; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_828 = 7'h36 == index[6:0] ? dirty_0_54 : _GEN_827; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_829 = 7'h37 == index[6:0] ? dirty_0_55 : _GEN_828; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_830 = 7'h38 == index[6:0] ? dirty_0_56 : _GEN_829; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_831 = 7'h39 == index[6:0] ? dirty_0_57 : _GEN_830; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_832 = 7'h3a == index[6:0] ? dirty_0_58 : _GEN_831; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_833 = 7'h3b == index[6:0] ? dirty_0_59 : _GEN_832; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_834 = 7'h3c == index[6:0] ? dirty_0_60 : _GEN_833; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_835 = 7'h3d == index[6:0] ? dirty_0_61 : _GEN_834; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_836 = 7'h3e == index[6:0] ? dirty_0_62 : _GEN_835; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_837 = 7'h3f == index[6:0] ? dirty_0_63 : _GEN_836; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_838 = 7'h40 == index[6:0] ? dirty_0_64 : _GEN_837; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_839 = 7'h41 == index[6:0] ? dirty_0_65 : _GEN_838; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_840 = 7'h42 == index[6:0] ? dirty_0_66 : _GEN_839; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_841 = 7'h43 == index[6:0] ? dirty_0_67 : _GEN_840; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_842 = 7'h44 == index[6:0] ? dirty_0_68 : _GEN_841; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_843 = 7'h45 == index[6:0] ? dirty_0_69 : _GEN_842; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_844 = 7'h46 == index[6:0] ? dirty_0_70 : _GEN_843; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_845 = 7'h47 == index[6:0] ? dirty_0_71 : _GEN_844; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_846 = 7'h48 == index[6:0] ? dirty_0_72 : _GEN_845; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_847 = 7'h49 == index[6:0] ? dirty_0_73 : _GEN_846; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_848 = 7'h4a == index[6:0] ? dirty_0_74 : _GEN_847; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_849 = 7'h4b == index[6:0] ? dirty_0_75 : _GEN_848; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_850 = 7'h4c == index[6:0] ? dirty_0_76 : _GEN_849; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_851 = 7'h4d == index[6:0] ? dirty_0_77 : _GEN_850; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_852 = 7'h4e == index[6:0] ? dirty_0_78 : _GEN_851; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_853 = 7'h4f == index[6:0] ? dirty_0_79 : _GEN_852; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_854 = 7'h50 == index[6:0] ? dirty_0_80 : _GEN_853; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_855 = 7'h51 == index[6:0] ? dirty_0_81 : _GEN_854; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_856 = 7'h52 == index[6:0] ? dirty_0_82 : _GEN_855; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_857 = 7'h53 == index[6:0] ? dirty_0_83 : _GEN_856; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_858 = 7'h54 == index[6:0] ? dirty_0_84 : _GEN_857; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_859 = 7'h55 == index[6:0] ? dirty_0_85 : _GEN_858; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_860 = 7'h56 == index[6:0] ? dirty_0_86 : _GEN_859; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_861 = 7'h57 == index[6:0] ? dirty_0_87 : _GEN_860; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_862 = 7'h58 == index[6:0] ? dirty_0_88 : _GEN_861; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_863 = 7'h59 == index[6:0] ? dirty_0_89 : _GEN_862; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_864 = 7'h5a == index[6:0] ? dirty_0_90 : _GEN_863; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_865 = 7'h5b == index[6:0] ? dirty_0_91 : _GEN_864; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_866 = 7'h5c == index[6:0] ? dirty_0_92 : _GEN_865; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_867 = 7'h5d == index[6:0] ? dirty_0_93 : _GEN_866; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_868 = 7'h5e == index[6:0] ? dirty_0_94 : _GEN_867; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_869 = 7'h5f == index[6:0] ? dirty_0_95 : _GEN_868; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_870 = 7'h60 == index[6:0] ? dirty_0_96 : _GEN_869; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_871 = 7'h61 == index[6:0] ? dirty_0_97 : _GEN_870; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_872 = 7'h62 == index[6:0] ? dirty_0_98 : _GEN_871; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_873 = 7'h63 == index[6:0] ? dirty_0_99 : _GEN_872; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_874 = 7'h64 == index[6:0] ? dirty_0_100 : _GEN_873; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_875 = 7'h65 == index[6:0] ? dirty_0_101 : _GEN_874; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_876 = 7'h66 == index[6:0] ? dirty_0_102 : _GEN_875; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_877 = 7'h67 == index[6:0] ? dirty_0_103 : _GEN_876; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_878 = 7'h68 == index[6:0] ? dirty_0_104 : _GEN_877; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_879 = 7'h69 == index[6:0] ? dirty_0_105 : _GEN_878; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_880 = 7'h6a == index[6:0] ? dirty_0_106 : _GEN_879; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_881 = 7'h6b == index[6:0] ? dirty_0_107 : _GEN_880; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_882 = 7'h6c == index[6:0] ? dirty_0_108 : _GEN_881; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_883 = 7'h6d == index[6:0] ? dirty_0_109 : _GEN_882; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_884 = 7'h6e == index[6:0] ? dirty_0_110 : _GEN_883; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_885 = 7'h6f == index[6:0] ? dirty_0_111 : _GEN_884; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_886 = 7'h70 == index[6:0] ? dirty_0_112 : _GEN_885; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_887 = 7'h71 == index[6:0] ? dirty_0_113 : _GEN_886; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_888 = 7'h72 == index[6:0] ? dirty_0_114 : _GEN_887; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_889 = 7'h73 == index[6:0] ? dirty_0_115 : _GEN_888; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_890 = 7'h74 == index[6:0] ? dirty_0_116 : _GEN_889; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_891 = 7'h75 == index[6:0] ? dirty_0_117 : _GEN_890; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_892 = 7'h76 == index[6:0] ? dirty_0_118 : _GEN_891; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_893 = 7'h77 == index[6:0] ? dirty_0_119 : _GEN_892; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_894 = 7'h78 == index[6:0] ? dirty_0_120 : _GEN_893; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_895 = 7'h79 == index[6:0] ? dirty_0_121 : _GEN_894; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_896 = 7'h7a == index[6:0] ? dirty_0_122 : _GEN_895; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_897 = 7'h7b == index[6:0] ? dirty_0_123 : _GEN_896; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_898 = 7'h7c == index[6:0] ? dirty_0_124 : _GEN_897; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_899 = 7'h7d == index[6:0] ? dirty_0_125 : _GEN_898; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_900 = 7'h7e == index[6:0] ? dirty_0_126 : _GEN_899; // @[d_cache.scala 90:{27,27}]
  wire  _GEN_901 = 7'h7f == index[6:0] ? dirty_0_127 : _GEN_900; // @[d_cache.scala 90:{27,27}]
  wire [2:0] _GEN_902 = io_from_lsu_rready ? 3'h0 : state; // @[d_cache.scala 73:24 89:41 91:27]
  wire  _GEN_904 = 7'h1 == index[6:0] ? dirty_1_1 : dirty_1_0; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_905 = 7'h2 == index[6:0] ? dirty_1_2 : _GEN_904; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_906 = 7'h3 == index[6:0] ? dirty_1_3 : _GEN_905; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_907 = 7'h4 == index[6:0] ? dirty_1_4 : _GEN_906; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_908 = 7'h5 == index[6:0] ? dirty_1_5 : _GEN_907; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_909 = 7'h6 == index[6:0] ? dirty_1_6 : _GEN_908; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_910 = 7'h7 == index[6:0] ? dirty_1_7 : _GEN_909; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_911 = 7'h8 == index[6:0] ? dirty_1_8 : _GEN_910; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_912 = 7'h9 == index[6:0] ? dirty_1_9 : _GEN_911; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_913 = 7'ha == index[6:0] ? dirty_1_10 : _GEN_912; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_914 = 7'hb == index[6:0] ? dirty_1_11 : _GEN_913; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_915 = 7'hc == index[6:0] ? dirty_1_12 : _GEN_914; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_916 = 7'hd == index[6:0] ? dirty_1_13 : _GEN_915; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_917 = 7'he == index[6:0] ? dirty_1_14 : _GEN_916; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_918 = 7'hf == index[6:0] ? dirty_1_15 : _GEN_917; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_919 = 7'h10 == index[6:0] ? dirty_1_16 : _GEN_918; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_920 = 7'h11 == index[6:0] ? dirty_1_17 : _GEN_919; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_921 = 7'h12 == index[6:0] ? dirty_1_18 : _GEN_920; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_922 = 7'h13 == index[6:0] ? dirty_1_19 : _GEN_921; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_923 = 7'h14 == index[6:0] ? dirty_1_20 : _GEN_922; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_924 = 7'h15 == index[6:0] ? dirty_1_21 : _GEN_923; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_925 = 7'h16 == index[6:0] ? dirty_1_22 : _GEN_924; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_926 = 7'h17 == index[6:0] ? dirty_1_23 : _GEN_925; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_927 = 7'h18 == index[6:0] ? dirty_1_24 : _GEN_926; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_928 = 7'h19 == index[6:0] ? dirty_1_25 : _GEN_927; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_929 = 7'h1a == index[6:0] ? dirty_1_26 : _GEN_928; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_930 = 7'h1b == index[6:0] ? dirty_1_27 : _GEN_929; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_931 = 7'h1c == index[6:0] ? dirty_1_28 : _GEN_930; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_932 = 7'h1d == index[6:0] ? dirty_1_29 : _GEN_931; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_933 = 7'h1e == index[6:0] ? dirty_1_30 : _GEN_932; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_934 = 7'h1f == index[6:0] ? dirty_1_31 : _GEN_933; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_935 = 7'h20 == index[6:0] ? dirty_1_32 : _GEN_934; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_936 = 7'h21 == index[6:0] ? dirty_1_33 : _GEN_935; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_937 = 7'h22 == index[6:0] ? dirty_1_34 : _GEN_936; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_938 = 7'h23 == index[6:0] ? dirty_1_35 : _GEN_937; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_939 = 7'h24 == index[6:0] ? dirty_1_36 : _GEN_938; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_940 = 7'h25 == index[6:0] ? dirty_1_37 : _GEN_939; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_941 = 7'h26 == index[6:0] ? dirty_1_38 : _GEN_940; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_942 = 7'h27 == index[6:0] ? dirty_1_39 : _GEN_941; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_943 = 7'h28 == index[6:0] ? dirty_1_40 : _GEN_942; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_944 = 7'h29 == index[6:0] ? dirty_1_41 : _GEN_943; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_945 = 7'h2a == index[6:0] ? dirty_1_42 : _GEN_944; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_946 = 7'h2b == index[6:0] ? dirty_1_43 : _GEN_945; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_947 = 7'h2c == index[6:0] ? dirty_1_44 : _GEN_946; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_948 = 7'h2d == index[6:0] ? dirty_1_45 : _GEN_947; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_949 = 7'h2e == index[6:0] ? dirty_1_46 : _GEN_948; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_950 = 7'h2f == index[6:0] ? dirty_1_47 : _GEN_949; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_951 = 7'h30 == index[6:0] ? dirty_1_48 : _GEN_950; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_952 = 7'h31 == index[6:0] ? dirty_1_49 : _GEN_951; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_953 = 7'h32 == index[6:0] ? dirty_1_50 : _GEN_952; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_954 = 7'h33 == index[6:0] ? dirty_1_51 : _GEN_953; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_955 = 7'h34 == index[6:0] ? dirty_1_52 : _GEN_954; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_956 = 7'h35 == index[6:0] ? dirty_1_53 : _GEN_955; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_957 = 7'h36 == index[6:0] ? dirty_1_54 : _GEN_956; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_958 = 7'h37 == index[6:0] ? dirty_1_55 : _GEN_957; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_959 = 7'h38 == index[6:0] ? dirty_1_56 : _GEN_958; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_960 = 7'h39 == index[6:0] ? dirty_1_57 : _GEN_959; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_961 = 7'h3a == index[6:0] ? dirty_1_58 : _GEN_960; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_962 = 7'h3b == index[6:0] ? dirty_1_59 : _GEN_961; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_963 = 7'h3c == index[6:0] ? dirty_1_60 : _GEN_962; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_964 = 7'h3d == index[6:0] ? dirty_1_61 : _GEN_963; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_965 = 7'h3e == index[6:0] ? dirty_1_62 : _GEN_964; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_966 = 7'h3f == index[6:0] ? dirty_1_63 : _GEN_965; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_967 = 7'h40 == index[6:0] ? dirty_1_64 : _GEN_966; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_968 = 7'h41 == index[6:0] ? dirty_1_65 : _GEN_967; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_969 = 7'h42 == index[6:0] ? dirty_1_66 : _GEN_968; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_970 = 7'h43 == index[6:0] ? dirty_1_67 : _GEN_969; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_971 = 7'h44 == index[6:0] ? dirty_1_68 : _GEN_970; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_972 = 7'h45 == index[6:0] ? dirty_1_69 : _GEN_971; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_973 = 7'h46 == index[6:0] ? dirty_1_70 : _GEN_972; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_974 = 7'h47 == index[6:0] ? dirty_1_71 : _GEN_973; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_975 = 7'h48 == index[6:0] ? dirty_1_72 : _GEN_974; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_976 = 7'h49 == index[6:0] ? dirty_1_73 : _GEN_975; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_977 = 7'h4a == index[6:0] ? dirty_1_74 : _GEN_976; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_978 = 7'h4b == index[6:0] ? dirty_1_75 : _GEN_977; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_979 = 7'h4c == index[6:0] ? dirty_1_76 : _GEN_978; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_980 = 7'h4d == index[6:0] ? dirty_1_77 : _GEN_979; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_981 = 7'h4e == index[6:0] ? dirty_1_78 : _GEN_980; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_982 = 7'h4f == index[6:0] ? dirty_1_79 : _GEN_981; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_983 = 7'h50 == index[6:0] ? dirty_1_80 : _GEN_982; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_984 = 7'h51 == index[6:0] ? dirty_1_81 : _GEN_983; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_985 = 7'h52 == index[6:0] ? dirty_1_82 : _GEN_984; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_986 = 7'h53 == index[6:0] ? dirty_1_83 : _GEN_985; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_987 = 7'h54 == index[6:0] ? dirty_1_84 : _GEN_986; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_988 = 7'h55 == index[6:0] ? dirty_1_85 : _GEN_987; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_989 = 7'h56 == index[6:0] ? dirty_1_86 : _GEN_988; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_990 = 7'h57 == index[6:0] ? dirty_1_87 : _GEN_989; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_991 = 7'h58 == index[6:0] ? dirty_1_88 : _GEN_990; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_992 = 7'h59 == index[6:0] ? dirty_1_89 : _GEN_991; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_993 = 7'h5a == index[6:0] ? dirty_1_90 : _GEN_992; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_994 = 7'h5b == index[6:0] ? dirty_1_91 : _GEN_993; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_995 = 7'h5c == index[6:0] ? dirty_1_92 : _GEN_994; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_996 = 7'h5d == index[6:0] ? dirty_1_93 : _GEN_995; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_997 = 7'h5e == index[6:0] ? dirty_1_94 : _GEN_996; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_998 = 7'h5f == index[6:0] ? dirty_1_95 : _GEN_997; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_999 = 7'h60 == index[6:0] ? dirty_1_96 : _GEN_998; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1000 = 7'h61 == index[6:0] ? dirty_1_97 : _GEN_999; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1001 = 7'h62 == index[6:0] ? dirty_1_98 : _GEN_1000; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1002 = 7'h63 == index[6:0] ? dirty_1_99 : _GEN_1001; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1003 = 7'h64 == index[6:0] ? dirty_1_100 : _GEN_1002; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1004 = 7'h65 == index[6:0] ? dirty_1_101 : _GEN_1003; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1005 = 7'h66 == index[6:0] ? dirty_1_102 : _GEN_1004; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1006 = 7'h67 == index[6:0] ? dirty_1_103 : _GEN_1005; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1007 = 7'h68 == index[6:0] ? dirty_1_104 : _GEN_1006; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1008 = 7'h69 == index[6:0] ? dirty_1_105 : _GEN_1007; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1009 = 7'h6a == index[6:0] ? dirty_1_106 : _GEN_1008; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1010 = 7'h6b == index[6:0] ? dirty_1_107 : _GEN_1009; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1011 = 7'h6c == index[6:0] ? dirty_1_108 : _GEN_1010; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1012 = 7'h6d == index[6:0] ? dirty_1_109 : _GEN_1011; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1013 = 7'h6e == index[6:0] ? dirty_1_110 : _GEN_1012; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1014 = 7'h6f == index[6:0] ? dirty_1_111 : _GEN_1013; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1015 = 7'h70 == index[6:0] ? dirty_1_112 : _GEN_1014; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1016 = 7'h71 == index[6:0] ? dirty_1_113 : _GEN_1015; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1017 = 7'h72 == index[6:0] ? dirty_1_114 : _GEN_1016; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1018 = 7'h73 == index[6:0] ? dirty_1_115 : _GEN_1017; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1019 = 7'h74 == index[6:0] ? dirty_1_116 : _GEN_1018; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1020 = 7'h75 == index[6:0] ? dirty_1_117 : _GEN_1019; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1021 = 7'h76 == index[6:0] ? dirty_1_118 : _GEN_1020; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1022 = 7'h77 == index[6:0] ? dirty_1_119 : _GEN_1021; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1023 = 7'h78 == index[6:0] ? dirty_1_120 : _GEN_1022; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1024 = 7'h79 == index[6:0] ? dirty_1_121 : _GEN_1023; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1025 = 7'h7a == index[6:0] ? dirty_1_122 : _GEN_1024; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1026 = 7'h7b == index[6:0] ? dirty_1_123 : _GEN_1025; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1027 = 7'h7c == index[6:0] ? dirty_1_124 : _GEN_1026; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1028 = 7'h7d == index[6:0] ? dirty_1_125 : _GEN_1027; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1029 = 7'h7e == index[6:0] ? dirty_1_126 : _GEN_1028; // @[d_cache.scala 96:{27,27}]
  wire  _GEN_1030 = 7'h7f == index[6:0] ? dirty_1_127 : _GEN_1029; // @[d_cache.scala 96:{27,27}]
  wire [2:0] _GEN_1031 = way1_hit ? _GEN_902 : 3'h3; // @[d_cache.scala 100:23 94:33]
  wire [63:0] _GEN_16803 = {{32'd0}, io_from_lsu_wdata}; // @[d_cache.scala 106:53]
  wire [63:0] _ram_0_T = _GEN_16803 & wmask; // @[d_cache.scala 106:53]
  wire [126:0] _GEN_17844 = {{63'd0}, _ram_0_T}; // @[d_cache.scala 106:62]
  wire [126:0] _ram_0_T_1 = _GEN_17844 << shift_bit; // @[d_cache.scala 106:62]
  wire [126:0] _GEN_17845 = {{63'd0}, wmask}; // @[d_cache.scala 106:102]
  wire [126:0] _ram_0_T_3 = _GEN_17845 << shift_bit; // @[d_cache.scala 106:102]
  wire [126:0] _ram_0_T_4 = ~_ram_0_T_3; // @[d_cache.scala 106:94]
  wire [63:0] _GEN_1034 = 7'h1 == index[6:0] ? ram_0_1 : ram_0_0; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1035 = 7'h2 == index[6:0] ? ram_0_2 : _GEN_1034; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1036 = 7'h3 == index[6:0] ? ram_0_3 : _GEN_1035; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1037 = 7'h4 == index[6:0] ? ram_0_4 : _GEN_1036; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1038 = 7'h5 == index[6:0] ? ram_0_5 : _GEN_1037; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1039 = 7'h6 == index[6:0] ? ram_0_6 : _GEN_1038; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1040 = 7'h7 == index[6:0] ? ram_0_7 : _GEN_1039; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1041 = 7'h8 == index[6:0] ? ram_0_8 : _GEN_1040; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1042 = 7'h9 == index[6:0] ? ram_0_9 : _GEN_1041; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1043 = 7'ha == index[6:0] ? ram_0_10 : _GEN_1042; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1044 = 7'hb == index[6:0] ? ram_0_11 : _GEN_1043; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1045 = 7'hc == index[6:0] ? ram_0_12 : _GEN_1044; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1046 = 7'hd == index[6:0] ? ram_0_13 : _GEN_1045; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1047 = 7'he == index[6:0] ? ram_0_14 : _GEN_1046; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1048 = 7'hf == index[6:0] ? ram_0_15 : _GEN_1047; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1049 = 7'h10 == index[6:0] ? ram_0_16 : _GEN_1048; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1050 = 7'h11 == index[6:0] ? ram_0_17 : _GEN_1049; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1051 = 7'h12 == index[6:0] ? ram_0_18 : _GEN_1050; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1052 = 7'h13 == index[6:0] ? ram_0_19 : _GEN_1051; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1053 = 7'h14 == index[6:0] ? ram_0_20 : _GEN_1052; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1054 = 7'h15 == index[6:0] ? ram_0_21 : _GEN_1053; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1055 = 7'h16 == index[6:0] ? ram_0_22 : _GEN_1054; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1056 = 7'h17 == index[6:0] ? ram_0_23 : _GEN_1055; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1057 = 7'h18 == index[6:0] ? ram_0_24 : _GEN_1056; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1058 = 7'h19 == index[6:0] ? ram_0_25 : _GEN_1057; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1059 = 7'h1a == index[6:0] ? ram_0_26 : _GEN_1058; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1060 = 7'h1b == index[6:0] ? ram_0_27 : _GEN_1059; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1061 = 7'h1c == index[6:0] ? ram_0_28 : _GEN_1060; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1062 = 7'h1d == index[6:0] ? ram_0_29 : _GEN_1061; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1063 = 7'h1e == index[6:0] ? ram_0_30 : _GEN_1062; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1064 = 7'h1f == index[6:0] ? ram_0_31 : _GEN_1063; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1065 = 7'h20 == index[6:0] ? ram_0_32 : _GEN_1064; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1066 = 7'h21 == index[6:0] ? ram_0_33 : _GEN_1065; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1067 = 7'h22 == index[6:0] ? ram_0_34 : _GEN_1066; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1068 = 7'h23 == index[6:0] ? ram_0_35 : _GEN_1067; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1069 = 7'h24 == index[6:0] ? ram_0_36 : _GEN_1068; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1070 = 7'h25 == index[6:0] ? ram_0_37 : _GEN_1069; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1071 = 7'h26 == index[6:0] ? ram_0_38 : _GEN_1070; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1072 = 7'h27 == index[6:0] ? ram_0_39 : _GEN_1071; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1073 = 7'h28 == index[6:0] ? ram_0_40 : _GEN_1072; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1074 = 7'h29 == index[6:0] ? ram_0_41 : _GEN_1073; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1075 = 7'h2a == index[6:0] ? ram_0_42 : _GEN_1074; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1076 = 7'h2b == index[6:0] ? ram_0_43 : _GEN_1075; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1077 = 7'h2c == index[6:0] ? ram_0_44 : _GEN_1076; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1078 = 7'h2d == index[6:0] ? ram_0_45 : _GEN_1077; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1079 = 7'h2e == index[6:0] ? ram_0_46 : _GEN_1078; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1080 = 7'h2f == index[6:0] ? ram_0_47 : _GEN_1079; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1081 = 7'h30 == index[6:0] ? ram_0_48 : _GEN_1080; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1082 = 7'h31 == index[6:0] ? ram_0_49 : _GEN_1081; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1083 = 7'h32 == index[6:0] ? ram_0_50 : _GEN_1082; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1084 = 7'h33 == index[6:0] ? ram_0_51 : _GEN_1083; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1085 = 7'h34 == index[6:0] ? ram_0_52 : _GEN_1084; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1086 = 7'h35 == index[6:0] ? ram_0_53 : _GEN_1085; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1087 = 7'h36 == index[6:0] ? ram_0_54 : _GEN_1086; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1088 = 7'h37 == index[6:0] ? ram_0_55 : _GEN_1087; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1089 = 7'h38 == index[6:0] ? ram_0_56 : _GEN_1088; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1090 = 7'h39 == index[6:0] ? ram_0_57 : _GEN_1089; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1091 = 7'h3a == index[6:0] ? ram_0_58 : _GEN_1090; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1092 = 7'h3b == index[6:0] ? ram_0_59 : _GEN_1091; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1093 = 7'h3c == index[6:0] ? ram_0_60 : _GEN_1092; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1094 = 7'h3d == index[6:0] ? ram_0_61 : _GEN_1093; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1095 = 7'h3e == index[6:0] ? ram_0_62 : _GEN_1094; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1096 = 7'h3f == index[6:0] ? ram_0_63 : _GEN_1095; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1097 = 7'h40 == index[6:0] ? ram_0_64 : _GEN_1096; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1098 = 7'h41 == index[6:0] ? ram_0_65 : _GEN_1097; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1099 = 7'h42 == index[6:0] ? ram_0_66 : _GEN_1098; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1100 = 7'h43 == index[6:0] ? ram_0_67 : _GEN_1099; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1101 = 7'h44 == index[6:0] ? ram_0_68 : _GEN_1100; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1102 = 7'h45 == index[6:0] ? ram_0_69 : _GEN_1101; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1103 = 7'h46 == index[6:0] ? ram_0_70 : _GEN_1102; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1104 = 7'h47 == index[6:0] ? ram_0_71 : _GEN_1103; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1105 = 7'h48 == index[6:0] ? ram_0_72 : _GEN_1104; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1106 = 7'h49 == index[6:0] ? ram_0_73 : _GEN_1105; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1107 = 7'h4a == index[6:0] ? ram_0_74 : _GEN_1106; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1108 = 7'h4b == index[6:0] ? ram_0_75 : _GEN_1107; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1109 = 7'h4c == index[6:0] ? ram_0_76 : _GEN_1108; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1110 = 7'h4d == index[6:0] ? ram_0_77 : _GEN_1109; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1111 = 7'h4e == index[6:0] ? ram_0_78 : _GEN_1110; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1112 = 7'h4f == index[6:0] ? ram_0_79 : _GEN_1111; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1113 = 7'h50 == index[6:0] ? ram_0_80 : _GEN_1112; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1114 = 7'h51 == index[6:0] ? ram_0_81 : _GEN_1113; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1115 = 7'h52 == index[6:0] ? ram_0_82 : _GEN_1114; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1116 = 7'h53 == index[6:0] ? ram_0_83 : _GEN_1115; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1117 = 7'h54 == index[6:0] ? ram_0_84 : _GEN_1116; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1118 = 7'h55 == index[6:0] ? ram_0_85 : _GEN_1117; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1119 = 7'h56 == index[6:0] ? ram_0_86 : _GEN_1118; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1120 = 7'h57 == index[6:0] ? ram_0_87 : _GEN_1119; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1121 = 7'h58 == index[6:0] ? ram_0_88 : _GEN_1120; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1122 = 7'h59 == index[6:0] ? ram_0_89 : _GEN_1121; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1123 = 7'h5a == index[6:0] ? ram_0_90 : _GEN_1122; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1124 = 7'h5b == index[6:0] ? ram_0_91 : _GEN_1123; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1125 = 7'h5c == index[6:0] ? ram_0_92 : _GEN_1124; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1126 = 7'h5d == index[6:0] ? ram_0_93 : _GEN_1125; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1127 = 7'h5e == index[6:0] ? ram_0_94 : _GEN_1126; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1128 = 7'h5f == index[6:0] ? ram_0_95 : _GEN_1127; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1129 = 7'h60 == index[6:0] ? ram_0_96 : _GEN_1128; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1130 = 7'h61 == index[6:0] ? ram_0_97 : _GEN_1129; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1131 = 7'h62 == index[6:0] ? ram_0_98 : _GEN_1130; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1132 = 7'h63 == index[6:0] ? ram_0_99 : _GEN_1131; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1133 = 7'h64 == index[6:0] ? ram_0_100 : _GEN_1132; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1134 = 7'h65 == index[6:0] ? ram_0_101 : _GEN_1133; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1135 = 7'h66 == index[6:0] ? ram_0_102 : _GEN_1134; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1136 = 7'h67 == index[6:0] ? ram_0_103 : _GEN_1135; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1137 = 7'h68 == index[6:0] ? ram_0_104 : _GEN_1136; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1138 = 7'h69 == index[6:0] ? ram_0_105 : _GEN_1137; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1139 = 7'h6a == index[6:0] ? ram_0_106 : _GEN_1138; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1140 = 7'h6b == index[6:0] ? ram_0_107 : _GEN_1139; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1141 = 7'h6c == index[6:0] ? ram_0_108 : _GEN_1140; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1142 = 7'h6d == index[6:0] ? ram_0_109 : _GEN_1141; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1143 = 7'h6e == index[6:0] ? ram_0_110 : _GEN_1142; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1144 = 7'h6f == index[6:0] ? ram_0_111 : _GEN_1143; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1145 = 7'h70 == index[6:0] ? ram_0_112 : _GEN_1144; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1146 = 7'h71 == index[6:0] ? ram_0_113 : _GEN_1145; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1147 = 7'h72 == index[6:0] ? ram_0_114 : _GEN_1146; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1148 = 7'h73 == index[6:0] ? ram_0_115 : _GEN_1147; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1149 = 7'h74 == index[6:0] ? ram_0_116 : _GEN_1148; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1150 = 7'h75 == index[6:0] ? ram_0_117 : _GEN_1149; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1151 = 7'h76 == index[6:0] ? ram_0_118 : _GEN_1150; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1152 = 7'h77 == index[6:0] ? ram_0_119 : _GEN_1151; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1153 = 7'h78 == index[6:0] ? ram_0_120 : _GEN_1152; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1154 = 7'h79 == index[6:0] ? ram_0_121 : _GEN_1153; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1155 = 7'h7a == index[6:0] ? ram_0_122 : _GEN_1154; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1156 = 7'h7b == index[6:0] ? ram_0_123 : _GEN_1155; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1157 = 7'h7c == index[6:0] ? ram_0_124 : _GEN_1156; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1158 = 7'h7d == index[6:0] ? ram_0_125 : _GEN_1157; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1159 = 7'h7e == index[6:0] ? ram_0_126 : _GEN_1158; // @[d_cache.scala 106:{92,92}]
  wire [63:0] _GEN_1160 = 7'h7f == index[6:0] ? ram_0_127 : _GEN_1159; // @[d_cache.scala 106:{92,92}]
  wire [126:0] _GEN_16804 = {{63'd0}, _GEN_1160}; // @[d_cache.scala 106:92]
  wire [126:0] _ram_0_T_5 = _GEN_16804 & _ram_0_T_4; // @[d_cache.scala 106:92]
  wire [126:0] _ram_0_T_6 = _ram_0_T_1 | _ram_0_T_5; // @[d_cache.scala 106:76]
  wire [63:0] _GEN_1161 = 7'h0 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_0; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1162 = 7'h1 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_1; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1163 = 7'h2 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_2; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1164 = 7'h3 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_3; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1165 = 7'h4 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_4; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1166 = 7'h5 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_5; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1167 = 7'h6 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_6; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1168 = 7'h7 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_7; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1169 = 7'h8 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_8; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1170 = 7'h9 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_9; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1171 = 7'ha == index[6:0] ? _ram_0_T_6[63:0] : ram_0_10; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1172 = 7'hb == index[6:0] ? _ram_0_T_6[63:0] : ram_0_11; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1173 = 7'hc == index[6:0] ? _ram_0_T_6[63:0] : ram_0_12; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1174 = 7'hd == index[6:0] ? _ram_0_T_6[63:0] : ram_0_13; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1175 = 7'he == index[6:0] ? _ram_0_T_6[63:0] : ram_0_14; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1176 = 7'hf == index[6:0] ? _ram_0_T_6[63:0] : ram_0_15; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1177 = 7'h10 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_16; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1178 = 7'h11 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_17; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1179 = 7'h12 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_18; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1180 = 7'h13 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_19; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1181 = 7'h14 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_20; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1182 = 7'h15 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_21; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1183 = 7'h16 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_22; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1184 = 7'h17 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_23; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1185 = 7'h18 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_24; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1186 = 7'h19 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_25; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1187 = 7'h1a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_26; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1188 = 7'h1b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_27; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1189 = 7'h1c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_28; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1190 = 7'h1d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_29; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1191 = 7'h1e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_30; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1192 = 7'h1f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_31; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1193 = 7'h20 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_32; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1194 = 7'h21 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_33; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1195 = 7'h22 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_34; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1196 = 7'h23 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_35; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1197 = 7'h24 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_36; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1198 = 7'h25 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_37; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1199 = 7'h26 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_38; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1200 = 7'h27 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_39; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1201 = 7'h28 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_40; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1202 = 7'h29 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_41; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1203 = 7'h2a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_42; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1204 = 7'h2b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_43; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1205 = 7'h2c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_44; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1206 = 7'h2d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_45; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1207 = 7'h2e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_46; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1208 = 7'h2f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_47; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1209 = 7'h30 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_48; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1210 = 7'h31 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_49; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1211 = 7'h32 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_50; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1212 = 7'h33 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_51; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1213 = 7'h34 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_52; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1214 = 7'h35 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_53; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1215 = 7'h36 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_54; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1216 = 7'h37 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_55; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1217 = 7'h38 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_56; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1218 = 7'h39 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_57; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1219 = 7'h3a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_58; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1220 = 7'h3b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_59; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1221 = 7'h3c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_60; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1222 = 7'h3d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_61; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1223 = 7'h3e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_62; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1224 = 7'h3f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_63; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1225 = 7'h40 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_64; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1226 = 7'h41 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_65; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1227 = 7'h42 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_66; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1228 = 7'h43 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_67; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1229 = 7'h44 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_68; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1230 = 7'h45 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_69; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1231 = 7'h46 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_70; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1232 = 7'h47 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_71; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1233 = 7'h48 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_72; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1234 = 7'h49 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_73; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1235 = 7'h4a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_74; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1236 = 7'h4b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_75; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1237 = 7'h4c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_76; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1238 = 7'h4d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_77; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1239 = 7'h4e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_78; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1240 = 7'h4f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_79; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1241 = 7'h50 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_80; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1242 = 7'h51 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_81; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1243 = 7'h52 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_82; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1244 = 7'h53 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_83; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1245 = 7'h54 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_84; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1246 = 7'h55 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_85; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1247 = 7'h56 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_86; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1248 = 7'h57 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_87; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1249 = 7'h58 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_88; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1250 = 7'h59 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_89; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1251 = 7'h5a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_90; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1252 = 7'h5b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_91; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1253 = 7'h5c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_92; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1254 = 7'h5d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_93; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1255 = 7'h5e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_94; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1256 = 7'h5f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_95; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1257 = 7'h60 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_96; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1258 = 7'h61 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_97; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1259 = 7'h62 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_98; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1260 = 7'h63 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_99; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1261 = 7'h64 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_100; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1262 = 7'h65 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_101; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1263 = 7'h66 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_102; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1264 = 7'h67 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_103; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1265 = 7'h68 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_104; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1266 = 7'h69 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_105; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1267 = 7'h6a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_106; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1268 = 7'h6b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_107; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1269 = 7'h6c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_108; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1270 = 7'h6d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_109; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1271 = 7'h6e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_110; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1272 = 7'h6f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_111; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1273 = 7'h70 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_112; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1274 = 7'h71 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_113; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1275 = 7'h72 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_114; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1276 = 7'h73 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_115; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1277 = 7'h74 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_116; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1278 = 7'h75 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_117; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1279 = 7'h76 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_118; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1280 = 7'h77 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_119; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1281 = 7'h78 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_120; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1282 = 7'h79 == index[6:0] ? _ram_0_T_6[63:0] : ram_0_121; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1283 = 7'h7a == index[6:0] ? _ram_0_T_6[63:0] : ram_0_122; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1284 = 7'h7b == index[6:0] ? _ram_0_T_6[63:0] : ram_0_123; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1285 = 7'h7c == index[6:0] ? _ram_0_T_6[63:0] : ram_0_124; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1286 = 7'h7d == index[6:0] ? _ram_0_T_6[63:0] : ram_0_125; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1287 = 7'h7e == index[6:0] ? _ram_0_T_6[63:0] : ram_0_126; // @[d_cache.scala 106:{30,30} 18:24]
  wire [63:0] _GEN_1288 = 7'h7f == index[6:0] ? _ram_0_T_6[63:0] : ram_0_127; // @[d_cache.scala 106:{30,30} 18:24]
  wire  _GEN_16805 = 7'h0 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1289 = 7'h0 == index[6:0] | dirty_0_0; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16806 = 7'h1 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1290 = 7'h1 == index[6:0] | dirty_0_1; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16807 = 7'h2 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1291 = 7'h2 == index[6:0] | dirty_0_2; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16808 = 7'h3 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1292 = 7'h3 == index[6:0] | dirty_0_3; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16809 = 7'h4 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1293 = 7'h4 == index[6:0] | dirty_0_4; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16810 = 7'h5 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1294 = 7'h5 == index[6:0] | dirty_0_5; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16811 = 7'h6 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1295 = 7'h6 == index[6:0] | dirty_0_6; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16812 = 7'h7 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1296 = 7'h7 == index[6:0] | dirty_0_7; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16813 = 7'h8 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1297 = 7'h8 == index[6:0] | dirty_0_8; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16814 = 7'h9 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1298 = 7'h9 == index[6:0] | dirty_0_9; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16815 = 7'ha == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1299 = 7'ha == index[6:0] | dirty_0_10; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16816 = 7'hb == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1300 = 7'hb == index[6:0] | dirty_0_11; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16817 = 7'hc == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1301 = 7'hc == index[6:0] | dirty_0_12; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16818 = 7'hd == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1302 = 7'hd == index[6:0] | dirty_0_13; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16819 = 7'he == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1303 = 7'he == index[6:0] | dirty_0_14; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16820 = 7'hf == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1304 = 7'hf == index[6:0] | dirty_0_15; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16821 = 7'h10 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1305 = 7'h10 == index[6:0] | dirty_0_16; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16822 = 7'h11 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1306 = 7'h11 == index[6:0] | dirty_0_17; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16823 = 7'h12 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1307 = 7'h12 == index[6:0] | dirty_0_18; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16824 = 7'h13 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1308 = 7'h13 == index[6:0] | dirty_0_19; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16825 = 7'h14 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1309 = 7'h14 == index[6:0] | dirty_0_20; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16826 = 7'h15 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1310 = 7'h15 == index[6:0] | dirty_0_21; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16827 = 7'h16 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1311 = 7'h16 == index[6:0] | dirty_0_22; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16828 = 7'h17 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1312 = 7'h17 == index[6:0] | dirty_0_23; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16829 = 7'h18 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1313 = 7'h18 == index[6:0] | dirty_0_24; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16830 = 7'h19 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1314 = 7'h19 == index[6:0] | dirty_0_25; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16831 = 7'h1a == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1315 = 7'h1a == index[6:0] | dirty_0_26; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16832 = 7'h1b == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1316 = 7'h1b == index[6:0] | dirty_0_27; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16833 = 7'h1c == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1317 = 7'h1c == index[6:0] | dirty_0_28; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16834 = 7'h1d == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1318 = 7'h1d == index[6:0] | dirty_0_29; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16835 = 7'h1e == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1319 = 7'h1e == index[6:0] | dirty_0_30; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16836 = 7'h1f == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1320 = 7'h1f == index[6:0] | dirty_0_31; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16837 = 7'h20 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1321 = 7'h20 == index[6:0] | dirty_0_32; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16838 = 7'h21 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1322 = 7'h21 == index[6:0] | dirty_0_33; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16839 = 7'h22 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1323 = 7'h22 == index[6:0] | dirty_0_34; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16840 = 7'h23 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1324 = 7'h23 == index[6:0] | dirty_0_35; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16841 = 7'h24 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1325 = 7'h24 == index[6:0] | dirty_0_36; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16842 = 7'h25 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1326 = 7'h25 == index[6:0] | dirty_0_37; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16843 = 7'h26 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1327 = 7'h26 == index[6:0] | dirty_0_38; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16844 = 7'h27 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1328 = 7'h27 == index[6:0] | dirty_0_39; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16845 = 7'h28 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1329 = 7'h28 == index[6:0] | dirty_0_40; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16846 = 7'h29 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1330 = 7'h29 == index[6:0] | dirty_0_41; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16847 = 7'h2a == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1331 = 7'h2a == index[6:0] | dirty_0_42; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16848 = 7'h2b == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1332 = 7'h2b == index[6:0] | dirty_0_43; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16849 = 7'h2c == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1333 = 7'h2c == index[6:0] | dirty_0_44; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16850 = 7'h2d == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1334 = 7'h2d == index[6:0] | dirty_0_45; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16851 = 7'h2e == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1335 = 7'h2e == index[6:0] | dirty_0_46; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16852 = 7'h2f == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1336 = 7'h2f == index[6:0] | dirty_0_47; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16853 = 7'h30 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1337 = 7'h30 == index[6:0] | dirty_0_48; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16854 = 7'h31 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1338 = 7'h31 == index[6:0] | dirty_0_49; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16855 = 7'h32 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1339 = 7'h32 == index[6:0] | dirty_0_50; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16856 = 7'h33 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1340 = 7'h33 == index[6:0] | dirty_0_51; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16857 = 7'h34 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1341 = 7'h34 == index[6:0] | dirty_0_52; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16858 = 7'h35 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1342 = 7'h35 == index[6:0] | dirty_0_53; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16859 = 7'h36 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1343 = 7'h36 == index[6:0] | dirty_0_54; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16860 = 7'h37 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1344 = 7'h37 == index[6:0] | dirty_0_55; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16861 = 7'h38 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1345 = 7'h38 == index[6:0] | dirty_0_56; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16862 = 7'h39 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1346 = 7'h39 == index[6:0] | dirty_0_57; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16863 = 7'h3a == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1347 = 7'h3a == index[6:0] | dirty_0_58; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16864 = 7'h3b == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1348 = 7'h3b == index[6:0] | dirty_0_59; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16865 = 7'h3c == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1349 = 7'h3c == index[6:0] | dirty_0_60; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16866 = 7'h3d == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1350 = 7'h3d == index[6:0] | dirty_0_61; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16867 = 7'h3e == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1351 = 7'h3e == index[6:0] | dirty_0_62; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16868 = 7'h3f == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1352 = 7'h3f == index[6:0] | dirty_0_63; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16869 = 7'h40 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1353 = 7'h40 == index[6:0] | dirty_0_64; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16870 = 7'h41 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1354 = 7'h41 == index[6:0] | dirty_0_65; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16871 = 7'h42 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1355 = 7'h42 == index[6:0] | dirty_0_66; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16872 = 7'h43 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1356 = 7'h43 == index[6:0] | dirty_0_67; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16873 = 7'h44 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1357 = 7'h44 == index[6:0] | dirty_0_68; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16874 = 7'h45 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1358 = 7'h45 == index[6:0] | dirty_0_69; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16875 = 7'h46 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1359 = 7'h46 == index[6:0] | dirty_0_70; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16876 = 7'h47 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1360 = 7'h47 == index[6:0] | dirty_0_71; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16877 = 7'h48 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1361 = 7'h48 == index[6:0] | dirty_0_72; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16878 = 7'h49 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1362 = 7'h49 == index[6:0] | dirty_0_73; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16879 = 7'h4a == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1363 = 7'h4a == index[6:0] | dirty_0_74; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16880 = 7'h4b == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1364 = 7'h4b == index[6:0] | dirty_0_75; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16881 = 7'h4c == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1365 = 7'h4c == index[6:0] | dirty_0_76; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16882 = 7'h4d == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1366 = 7'h4d == index[6:0] | dirty_0_77; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16883 = 7'h4e == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1367 = 7'h4e == index[6:0] | dirty_0_78; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16884 = 7'h4f == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1368 = 7'h4f == index[6:0] | dirty_0_79; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16885 = 7'h50 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1369 = 7'h50 == index[6:0] | dirty_0_80; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16886 = 7'h51 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1370 = 7'h51 == index[6:0] | dirty_0_81; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16887 = 7'h52 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1371 = 7'h52 == index[6:0] | dirty_0_82; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16888 = 7'h53 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1372 = 7'h53 == index[6:0] | dirty_0_83; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16889 = 7'h54 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1373 = 7'h54 == index[6:0] | dirty_0_84; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16890 = 7'h55 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1374 = 7'h55 == index[6:0] | dirty_0_85; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16891 = 7'h56 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1375 = 7'h56 == index[6:0] | dirty_0_86; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16892 = 7'h57 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1376 = 7'h57 == index[6:0] | dirty_0_87; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16893 = 7'h58 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1377 = 7'h58 == index[6:0] | dirty_0_88; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16894 = 7'h59 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1378 = 7'h59 == index[6:0] | dirty_0_89; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16895 = 7'h5a == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1379 = 7'h5a == index[6:0] | dirty_0_90; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16896 = 7'h5b == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1380 = 7'h5b == index[6:0] | dirty_0_91; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16897 = 7'h5c == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1381 = 7'h5c == index[6:0] | dirty_0_92; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16898 = 7'h5d == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1382 = 7'h5d == index[6:0] | dirty_0_93; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16899 = 7'h5e == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1383 = 7'h5e == index[6:0] | dirty_0_94; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16900 = 7'h5f == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1384 = 7'h5f == index[6:0] | dirty_0_95; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16901 = 7'h60 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1385 = 7'h60 == index[6:0] | dirty_0_96; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16902 = 7'h61 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1386 = 7'h61 == index[6:0] | dirty_0_97; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16903 = 7'h62 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1387 = 7'h62 == index[6:0] | dirty_0_98; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16904 = 7'h63 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1388 = 7'h63 == index[6:0] | dirty_0_99; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16905 = 7'h64 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1389 = 7'h64 == index[6:0] | dirty_0_100; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16906 = 7'h65 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1390 = 7'h65 == index[6:0] | dirty_0_101; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16907 = 7'h66 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1391 = 7'h66 == index[6:0] | dirty_0_102; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16908 = 7'h67 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1392 = 7'h67 == index[6:0] | dirty_0_103; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16909 = 7'h68 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1393 = 7'h68 == index[6:0] | dirty_0_104; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16910 = 7'h69 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1394 = 7'h69 == index[6:0] | dirty_0_105; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16911 = 7'h6a == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1395 = 7'h6a == index[6:0] | dirty_0_106; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16912 = 7'h6b == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1396 = 7'h6b == index[6:0] | dirty_0_107; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16913 = 7'h6c == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1397 = 7'h6c == index[6:0] | dirty_0_108; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16914 = 7'h6d == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1398 = 7'h6d == index[6:0] | dirty_0_109; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16915 = 7'h6e == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1399 = 7'h6e == index[6:0] | dirty_0_110; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16916 = 7'h6f == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1400 = 7'h6f == index[6:0] | dirty_0_111; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16917 = 7'h70 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1401 = 7'h70 == index[6:0] | dirty_0_112; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16918 = 7'h71 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1402 = 7'h71 == index[6:0] | dirty_0_113; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16919 = 7'h72 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1403 = 7'h72 == index[6:0] | dirty_0_114; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16920 = 7'h73 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1404 = 7'h73 == index[6:0] | dirty_0_115; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16921 = 7'h74 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1405 = 7'h74 == index[6:0] | dirty_0_116; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16922 = 7'h75 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1406 = 7'h75 == index[6:0] | dirty_0_117; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16923 = 7'h76 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1407 = 7'h76 == index[6:0] | dirty_0_118; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16924 = 7'h77 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1408 = 7'h77 == index[6:0] | dirty_0_119; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16925 = 7'h78 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1409 = 7'h78 == index[6:0] | dirty_0_120; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16926 = 7'h79 == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1410 = 7'h79 == index[6:0] | dirty_0_121; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16927 = 7'h7a == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1411 = 7'h7a == index[6:0] | dirty_0_122; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16928 = 7'h7b == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1412 = 7'h7b == index[6:0] | dirty_0_123; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16929 = 7'h7c == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1413 = 7'h7c == index[6:0] | dirty_0_124; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16930 = 7'h7d == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1414 = 7'h7d == index[6:0] | dirty_0_125; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16931 = 7'h7e == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1415 = 7'h7e == index[6:0] | dirty_0_126; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_16932 = 7'h7f == index[6:0]; // @[d_cache.scala 109:{32,32} 24:26]
  wire  _GEN_1416 = 7'h7f == index[6:0] | dirty_0_127; // @[d_cache.scala 109:{32,32} 24:26]
  wire [63:0] _GEN_1545 = 7'h0 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_0; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1546 = 7'h1 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_1; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1547 = 7'h2 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_2; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1548 = 7'h3 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_3; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1549 = 7'h4 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_4; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1550 = 7'h5 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_5; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1551 = 7'h6 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_6; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1552 = 7'h7 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_7; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1553 = 7'h8 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_8; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1554 = 7'h9 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_9; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1555 = 7'ha == index[6:0] ? _ram_0_T_6[63:0] : ram_1_10; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1556 = 7'hb == index[6:0] ? _ram_0_T_6[63:0] : ram_1_11; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1557 = 7'hc == index[6:0] ? _ram_0_T_6[63:0] : ram_1_12; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1558 = 7'hd == index[6:0] ? _ram_0_T_6[63:0] : ram_1_13; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1559 = 7'he == index[6:0] ? _ram_0_T_6[63:0] : ram_1_14; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1560 = 7'hf == index[6:0] ? _ram_0_T_6[63:0] : ram_1_15; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1561 = 7'h10 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_16; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1562 = 7'h11 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_17; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1563 = 7'h12 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_18; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1564 = 7'h13 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_19; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1565 = 7'h14 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_20; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1566 = 7'h15 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_21; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1567 = 7'h16 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_22; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1568 = 7'h17 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_23; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1569 = 7'h18 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_24; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1570 = 7'h19 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_25; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1571 = 7'h1a == index[6:0] ? _ram_0_T_6[63:0] : ram_1_26; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1572 = 7'h1b == index[6:0] ? _ram_0_T_6[63:0] : ram_1_27; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1573 = 7'h1c == index[6:0] ? _ram_0_T_6[63:0] : ram_1_28; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1574 = 7'h1d == index[6:0] ? _ram_0_T_6[63:0] : ram_1_29; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1575 = 7'h1e == index[6:0] ? _ram_0_T_6[63:0] : ram_1_30; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1576 = 7'h1f == index[6:0] ? _ram_0_T_6[63:0] : ram_1_31; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1577 = 7'h20 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_32; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1578 = 7'h21 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_33; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1579 = 7'h22 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_34; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1580 = 7'h23 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_35; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1581 = 7'h24 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_36; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1582 = 7'h25 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_37; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1583 = 7'h26 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_38; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1584 = 7'h27 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_39; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1585 = 7'h28 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_40; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1586 = 7'h29 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_41; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1587 = 7'h2a == index[6:0] ? _ram_0_T_6[63:0] : ram_1_42; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1588 = 7'h2b == index[6:0] ? _ram_0_T_6[63:0] : ram_1_43; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1589 = 7'h2c == index[6:0] ? _ram_0_T_6[63:0] : ram_1_44; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1590 = 7'h2d == index[6:0] ? _ram_0_T_6[63:0] : ram_1_45; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1591 = 7'h2e == index[6:0] ? _ram_0_T_6[63:0] : ram_1_46; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1592 = 7'h2f == index[6:0] ? _ram_0_T_6[63:0] : ram_1_47; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1593 = 7'h30 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_48; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1594 = 7'h31 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_49; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1595 = 7'h32 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_50; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1596 = 7'h33 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_51; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1597 = 7'h34 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_52; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1598 = 7'h35 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_53; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1599 = 7'h36 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_54; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1600 = 7'h37 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_55; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1601 = 7'h38 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_56; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1602 = 7'h39 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_57; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1603 = 7'h3a == index[6:0] ? _ram_0_T_6[63:0] : ram_1_58; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1604 = 7'h3b == index[6:0] ? _ram_0_T_6[63:0] : ram_1_59; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1605 = 7'h3c == index[6:0] ? _ram_0_T_6[63:0] : ram_1_60; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1606 = 7'h3d == index[6:0] ? _ram_0_T_6[63:0] : ram_1_61; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1607 = 7'h3e == index[6:0] ? _ram_0_T_6[63:0] : ram_1_62; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1608 = 7'h3f == index[6:0] ? _ram_0_T_6[63:0] : ram_1_63; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1609 = 7'h40 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_64; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1610 = 7'h41 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_65; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1611 = 7'h42 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_66; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1612 = 7'h43 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_67; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1613 = 7'h44 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_68; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1614 = 7'h45 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_69; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1615 = 7'h46 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_70; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1616 = 7'h47 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_71; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1617 = 7'h48 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_72; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1618 = 7'h49 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_73; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1619 = 7'h4a == index[6:0] ? _ram_0_T_6[63:0] : ram_1_74; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1620 = 7'h4b == index[6:0] ? _ram_0_T_6[63:0] : ram_1_75; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1621 = 7'h4c == index[6:0] ? _ram_0_T_6[63:0] : ram_1_76; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1622 = 7'h4d == index[6:0] ? _ram_0_T_6[63:0] : ram_1_77; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1623 = 7'h4e == index[6:0] ? _ram_0_T_6[63:0] : ram_1_78; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1624 = 7'h4f == index[6:0] ? _ram_0_T_6[63:0] : ram_1_79; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1625 = 7'h50 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_80; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1626 = 7'h51 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_81; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1627 = 7'h52 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_82; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1628 = 7'h53 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_83; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1629 = 7'h54 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_84; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1630 = 7'h55 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_85; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1631 = 7'h56 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_86; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1632 = 7'h57 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_87; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1633 = 7'h58 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_88; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1634 = 7'h59 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_89; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1635 = 7'h5a == index[6:0] ? _ram_0_T_6[63:0] : ram_1_90; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1636 = 7'h5b == index[6:0] ? _ram_0_T_6[63:0] : ram_1_91; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1637 = 7'h5c == index[6:0] ? _ram_0_T_6[63:0] : ram_1_92; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1638 = 7'h5d == index[6:0] ? _ram_0_T_6[63:0] : ram_1_93; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1639 = 7'h5e == index[6:0] ? _ram_0_T_6[63:0] : ram_1_94; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1640 = 7'h5f == index[6:0] ? _ram_0_T_6[63:0] : ram_1_95; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1641 = 7'h60 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_96; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1642 = 7'h61 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_97; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1643 = 7'h62 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_98; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1644 = 7'h63 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_99; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1645 = 7'h64 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_100; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1646 = 7'h65 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_101; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1647 = 7'h66 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_102; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1648 = 7'h67 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_103; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1649 = 7'h68 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_104; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1650 = 7'h69 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_105; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1651 = 7'h6a == index[6:0] ? _ram_0_T_6[63:0] : ram_1_106; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1652 = 7'h6b == index[6:0] ? _ram_0_T_6[63:0] : ram_1_107; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1653 = 7'h6c == index[6:0] ? _ram_0_T_6[63:0] : ram_1_108; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1654 = 7'h6d == index[6:0] ? _ram_0_T_6[63:0] : ram_1_109; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1655 = 7'h6e == index[6:0] ? _ram_0_T_6[63:0] : ram_1_110; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1656 = 7'h6f == index[6:0] ? _ram_0_T_6[63:0] : ram_1_111; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1657 = 7'h70 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_112; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1658 = 7'h71 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_113; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1659 = 7'h72 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_114; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1660 = 7'h73 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_115; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1661 = 7'h74 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_116; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1662 = 7'h75 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_117; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1663 = 7'h76 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_118; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1664 = 7'h77 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_119; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1665 = 7'h78 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_120; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1666 = 7'h79 == index[6:0] ? _ram_0_T_6[63:0] : ram_1_121; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1667 = 7'h7a == index[6:0] ? _ram_0_T_6[63:0] : ram_1_122; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1668 = 7'h7b == index[6:0] ? _ram_0_T_6[63:0] : ram_1_123; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1669 = 7'h7c == index[6:0] ? _ram_0_T_6[63:0] : ram_1_124; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1670 = 7'h7d == index[6:0] ? _ram_0_T_6[63:0] : ram_1_125; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1671 = 7'h7e == index[6:0] ? _ram_0_T_6[63:0] : ram_1_126; // @[d_cache.scala 113:{30,30} 19:24]
  wire [63:0] _GEN_1672 = 7'h7f == index[6:0] ? _ram_0_T_6[63:0] : ram_1_127; // @[d_cache.scala 113:{30,30} 19:24]
  wire  _GEN_1673 = _GEN_16805 | dirty_1_0; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1674 = _GEN_16806 | dirty_1_1; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1675 = _GEN_16807 | dirty_1_2; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1676 = _GEN_16808 | dirty_1_3; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1677 = _GEN_16809 | dirty_1_4; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1678 = _GEN_16810 | dirty_1_5; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1679 = _GEN_16811 | dirty_1_6; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1680 = _GEN_16812 | dirty_1_7; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1681 = _GEN_16813 | dirty_1_8; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1682 = _GEN_16814 | dirty_1_9; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1683 = _GEN_16815 | dirty_1_10; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1684 = _GEN_16816 | dirty_1_11; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1685 = _GEN_16817 | dirty_1_12; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1686 = _GEN_16818 | dirty_1_13; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1687 = _GEN_16819 | dirty_1_14; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1688 = _GEN_16820 | dirty_1_15; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1689 = _GEN_16821 | dirty_1_16; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1690 = _GEN_16822 | dirty_1_17; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1691 = _GEN_16823 | dirty_1_18; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1692 = _GEN_16824 | dirty_1_19; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1693 = _GEN_16825 | dirty_1_20; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1694 = _GEN_16826 | dirty_1_21; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1695 = _GEN_16827 | dirty_1_22; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1696 = _GEN_16828 | dirty_1_23; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1697 = _GEN_16829 | dirty_1_24; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1698 = _GEN_16830 | dirty_1_25; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1699 = _GEN_16831 | dirty_1_26; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1700 = _GEN_16832 | dirty_1_27; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1701 = _GEN_16833 | dirty_1_28; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1702 = _GEN_16834 | dirty_1_29; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1703 = _GEN_16835 | dirty_1_30; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1704 = _GEN_16836 | dirty_1_31; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1705 = _GEN_16837 | dirty_1_32; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1706 = _GEN_16838 | dirty_1_33; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1707 = _GEN_16839 | dirty_1_34; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1708 = _GEN_16840 | dirty_1_35; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1709 = _GEN_16841 | dirty_1_36; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1710 = _GEN_16842 | dirty_1_37; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1711 = _GEN_16843 | dirty_1_38; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1712 = _GEN_16844 | dirty_1_39; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1713 = _GEN_16845 | dirty_1_40; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1714 = _GEN_16846 | dirty_1_41; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1715 = _GEN_16847 | dirty_1_42; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1716 = _GEN_16848 | dirty_1_43; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1717 = _GEN_16849 | dirty_1_44; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1718 = _GEN_16850 | dirty_1_45; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1719 = _GEN_16851 | dirty_1_46; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1720 = _GEN_16852 | dirty_1_47; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1721 = _GEN_16853 | dirty_1_48; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1722 = _GEN_16854 | dirty_1_49; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1723 = _GEN_16855 | dirty_1_50; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1724 = _GEN_16856 | dirty_1_51; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1725 = _GEN_16857 | dirty_1_52; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1726 = _GEN_16858 | dirty_1_53; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1727 = _GEN_16859 | dirty_1_54; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1728 = _GEN_16860 | dirty_1_55; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1729 = _GEN_16861 | dirty_1_56; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1730 = _GEN_16862 | dirty_1_57; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1731 = _GEN_16863 | dirty_1_58; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1732 = _GEN_16864 | dirty_1_59; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1733 = _GEN_16865 | dirty_1_60; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1734 = _GEN_16866 | dirty_1_61; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1735 = _GEN_16867 | dirty_1_62; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1736 = _GEN_16868 | dirty_1_63; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1737 = _GEN_16869 | dirty_1_64; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1738 = _GEN_16870 | dirty_1_65; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1739 = _GEN_16871 | dirty_1_66; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1740 = _GEN_16872 | dirty_1_67; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1741 = _GEN_16873 | dirty_1_68; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1742 = _GEN_16874 | dirty_1_69; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1743 = _GEN_16875 | dirty_1_70; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1744 = _GEN_16876 | dirty_1_71; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1745 = _GEN_16877 | dirty_1_72; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1746 = _GEN_16878 | dirty_1_73; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1747 = _GEN_16879 | dirty_1_74; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1748 = _GEN_16880 | dirty_1_75; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1749 = _GEN_16881 | dirty_1_76; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1750 = _GEN_16882 | dirty_1_77; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1751 = _GEN_16883 | dirty_1_78; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1752 = _GEN_16884 | dirty_1_79; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1753 = _GEN_16885 | dirty_1_80; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1754 = _GEN_16886 | dirty_1_81; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1755 = _GEN_16887 | dirty_1_82; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1756 = _GEN_16888 | dirty_1_83; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1757 = _GEN_16889 | dirty_1_84; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1758 = _GEN_16890 | dirty_1_85; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1759 = _GEN_16891 | dirty_1_86; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1760 = _GEN_16892 | dirty_1_87; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1761 = _GEN_16893 | dirty_1_88; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1762 = _GEN_16894 | dirty_1_89; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1763 = _GEN_16895 | dirty_1_90; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1764 = _GEN_16896 | dirty_1_91; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1765 = _GEN_16897 | dirty_1_92; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1766 = _GEN_16898 | dirty_1_93; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1767 = _GEN_16899 | dirty_1_94; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1768 = _GEN_16900 | dirty_1_95; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1769 = _GEN_16901 | dirty_1_96; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1770 = _GEN_16902 | dirty_1_97; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1771 = _GEN_16903 | dirty_1_98; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1772 = _GEN_16904 | dirty_1_99; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1773 = _GEN_16905 | dirty_1_100; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1774 = _GEN_16906 | dirty_1_101; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1775 = _GEN_16907 | dirty_1_102; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1776 = _GEN_16908 | dirty_1_103; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1777 = _GEN_16909 | dirty_1_104; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1778 = _GEN_16910 | dirty_1_105; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1779 = _GEN_16911 | dirty_1_106; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1780 = _GEN_16912 | dirty_1_107; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1781 = _GEN_16913 | dirty_1_108; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1782 = _GEN_16914 | dirty_1_109; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1783 = _GEN_16915 | dirty_1_110; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1784 = _GEN_16916 | dirty_1_111; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1785 = _GEN_16917 | dirty_1_112; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1786 = _GEN_16918 | dirty_1_113; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1787 = _GEN_16919 | dirty_1_114; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1788 = _GEN_16920 | dirty_1_115; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1789 = _GEN_16921 | dirty_1_116; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1790 = _GEN_16922 | dirty_1_117; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1791 = _GEN_16923 | dirty_1_118; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1792 = _GEN_16924 | dirty_1_119; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1793 = _GEN_16925 | dirty_1_120; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1794 = _GEN_16926 | dirty_1_121; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1795 = _GEN_16927 | dirty_1_122; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1796 = _GEN_16928 | dirty_1_123; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1797 = _GEN_16929 | dirty_1_124; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1798 = _GEN_16930 | dirty_1_125; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1799 = _GEN_16931 | dirty_1_126; // @[d_cache.scala 115:{32,32} 25:26]
  wire  _GEN_1800 = _GEN_16932 | dirty_1_127; // @[d_cache.scala 115:{32,32} 25:26]
  wire [2:0] _GEN_1801 = way1_hit ? 3'h0 : 3'h4; // @[d_cache.scala 111:33 112:23 117:23]
  wire [63:0] _GEN_1802 = way1_hit ? _GEN_1545 : ram_1_0; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1803 = way1_hit ? _GEN_1546 : ram_1_1; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1804 = way1_hit ? _GEN_1547 : ram_1_2; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1805 = way1_hit ? _GEN_1548 : ram_1_3; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1806 = way1_hit ? _GEN_1549 : ram_1_4; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1807 = way1_hit ? _GEN_1550 : ram_1_5; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1808 = way1_hit ? _GEN_1551 : ram_1_6; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1809 = way1_hit ? _GEN_1552 : ram_1_7; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1810 = way1_hit ? _GEN_1553 : ram_1_8; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1811 = way1_hit ? _GEN_1554 : ram_1_9; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1812 = way1_hit ? _GEN_1555 : ram_1_10; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1813 = way1_hit ? _GEN_1556 : ram_1_11; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1814 = way1_hit ? _GEN_1557 : ram_1_12; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1815 = way1_hit ? _GEN_1558 : ram_1_13; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1816 = way1_hit ? _GEN_1559 : ram_1_14; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1817 = way1_hit ? _GEN_1560 : ram_1_15; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1818 = way1_hit ? _GEN_1561 : ram_1_16; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1819 = way1_hit ? _GEN_1562 : ram_1_17; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1820 = way1_hit ? _GEN_1563 : ram_1_18; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1821 = way1_hit ? _GEN_1564 : ram_1_19; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1822 = way1_hit ? _GEN_1565 : ram_1_20; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1823 = way1_hit ? _GEN_1566 : ram_1_21; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1824 = way1_hit ? _GEN_1567 : ram_1_22; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1825 = way1_hit ? _GEN_1568 : ram_1_23; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1826 = way1_hit ? _GEN_1569 : ram_1_24; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1827 = way1_hit ? _GEN_1570 : ram_1_25; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1828 = way1_hit ? _GEN_1571 : ram_1_26; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1829 = way1_hit ? _GEN_1572 : ram_1_27; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1830 = way1_hit ? _GEN_1573 : ram_1_28; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1831 = way1_hit ? _GEN_1574 : ram_1_29; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1832 = way1_hit ? _GEN_1575 : ram_1_30; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1833 = way1_hit ? _GEN_1576 : ram_1_31; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1834 = way1_hit ? _GEN_1577 : ram_1_32; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1835 = way1_hit ? _GEN_1578 : ram_1_33; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1836 = way1_hit ? _GEN_1579 : ram_1_34; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1837 = way1_hit ? _GEN_1580 : ram_1_35; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1838 = way1_hit ? _GEN_1581 : ram_1_36; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1839 = way1_hit ? _GEN_1582 : ram_1_37; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1840 = way1_hit ? _GEN_1583 : ram_1_38; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1841 = way1_hit ? _GEN_1584 : ram_1_39; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1842 = way1_hit ? _GEN_1585 : ram_1_40; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1843 = way1_hit ? _GEN_1586 : ram_1_41; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1844 = way1_hit ? _GEN_1587 : ram_1_42; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1845 = way1_hit ? _GEN_1588 : ram_1_43; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1846 = way1_hit ? _GEN_1589 : ram_1_44; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1847 = way1_hit ? _GEN_1590 : ram_1_45; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1848 = way1_hit ? _GEN_1591 : ram_1_46; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1849 = way1_hit ? _GEN_1592 : ram_1_47; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1850 = way1_hit ? _GEN_1593 : ram_1_48; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1851 = way1_hit ? _GEN_1594 : ram_1_49; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1852 = way1_hit ? _GEN_1595 : ram_1_50; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1853 = way1_hit ? _GEN_1596 : ram_1_51; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1854 = way1_hit ? _GEN_1597 : ram_1_52; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1855 = way1_hit ? _GEN_1598 : ram_1_53; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1856 = way1_hit ? _GEN_1599 : ram_1_54; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1857 = way1_hit ? _GEN_1600 : ram_1_55; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1858 = way1_hit ? _GEN_1601 : ram_1_56; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1859 = way1_hit ? _GEN_1602 : ram_1_57; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1860 = way1_hit ? _GEN_1603 : ram_1_58; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1861 = way1_hit ? _GEN_1604 : ram_1_59; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1862 = way1_hit ? _GEN_1605 : ram_1_60; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1863 = way1_hit ? _GEN_1606 : ram_1_61; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1864 = way1_hit ? _GEN_1607 : ram_1_62; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1865 = way1_hit ? _GEN_1608 : ram_1_63; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1866 = way1_hit ? _GEN_1609 : ram_1_64; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1867 = way1_hit ? _GEN_1610 : ram_1_65; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1868 = way1_hit ? _GEN_1611 : ram_1_66; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1869 = way1_hit ? _GEN_1612 : ram_1_67; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1870 = way1_hit ? _GEN_1613 : ram_1_68; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1871 = way1_hit ? _GEN_1614 : ram_1_69; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1872 = way1_hit ? _GEN_1615 : ram_1_70; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1873 = way1_hit ? _GEN_1616 : ram_1_71; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1874 = way1_hit ? _GEN_1617 : ram_1_72; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1875 = way1_hit ? _GEN_1618 : ram_1_73; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1876 = way1_hit ? _GEN_1619 : ram_1_74; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1877 = way1_hit ? _GEN_1620 : ram_1_75; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1878 = way1_hit ? _GEN_1621 : ram_1_76; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1879 = way1_hit ? _GEN_1622 : ram_1_77; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1880 = way1_hit ? _GEN_1623 : ram_1_78; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1881 = way1_hit ? _GEN_1624 : ram_1_79; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1882 = way1_hit ? _GEN_1625 : ram_1_80; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1883 = way1_hit ? _GEN_1626 : ram_1_81; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1884 = way1_hit ? _GEN_1627 : ram_1_82; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1885 = way1_hit ? _GEN_1628 : ram_1_83; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1886 = way1_hit ? _GEN_1629 : ram_1_84; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1887 = way1_hit ? _GEN_1630 : ram_1_85; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1888 = way1_hit ? _GEN_1631 : ram_1_86; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1889 = way1_hit ? _GEN_1632 : ram_1_87; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1890 = way1_hit ? _GEN_1633 : ram_1_88; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1891 = way1_hit ? _GEN_1634 : ram_1_89; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1892 = way1_hit ? _GEN_1635 : ram_1_90; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1893 = way1_hit ? _GEN_1636 : ram_1_91; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1894 = way1_hit ? _GEN_1637 : ram_1_92; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1895 = way1_hit ? _GEN_1638 : ram_1_93; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1896 = way1_hit ? _GEN_1639 : ram_1_94; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1897 = way1_hit ? _GEN_1640 : ram_1_95; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1898 = way1_hit ? _GEN_1641 : ram_1_96; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1899 = way1_hit ? _GEN_1642 : ram_1_97; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1900 = way1_hit ? _GEN_1643 : ram_1_98; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1901 = way1_hit ? _GEN_1644 : ram_1_99; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1902 = way1_hit ? _GEN_1645 : ram_1_100; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1903 = way1_hit ? _GEN_1646 : ram_1_101; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1904 = way1_hit ? _GEN_1647 : ram_1_102; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1905 = way1_hit ? _GEN_1648 : ram_1_103; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1906 = way1_hit ? _GEN_1649 : ram_1_104; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1907 = way1_hit ? _GEN_1650 : ram_1_105; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1908 = way1_hit ? _GEN_1651 : ram_1_106; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1909 = way1_hit ? _GEN_1652 : ram_1_107; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1910 = way1_hit ? _GEN_1653 : ram_1_108; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1911 = way1_hit ? _GEN_1654 : ram_1_109; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1912 = way1_hit ? _GEN_1655 : ram_1_110; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1913 = way1_hit ? _GEN_1656 : ram_1_111; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1914 = way1_hit ? _GEN_1657 : ram_1_112; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1915 = way1_hit ? _GEN_1658 : ram_1_113; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1916 = way1_hit ? _GEN_1659 : ram_1_114; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1917 = way1_hit ? _GEN_1660 : ram_1_115; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1918 = way1_hit ? _GEN_1661 : ram_1_116; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1919 = way1_hit ? _GEN_1662 : ram_1_117; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1920 = way1_hit ? _GEN_1663 : ram_1_118; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1921 = way1_hit ? _GEN_1664 : ram_1_119; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1922 = way1_hit ? _GEN_1665 : ram_1_120; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1923 = way1_hit ? _GEN_1666 : ram_1_121; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1924 = way1_hit ? _GEN_1667 : ram_1_122; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1925 = way1_hit ? _GEN_1668 : ram_1_123; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1926 = way1_hit ? _GEN_1669 : ram_1_124; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1927 = way1_hit ? _GEN_1670 : ram_1_125; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1928 = way1_hit ? _GEN_1671 : ram_1_126; // @[d_cache.scala 111:33 19:24]
  wire [63:0] _GEN_1929 = way1_hit ? _GEN_1672 : ram_1_127; // @[d_cache.scala 111:33 19:24]
  wire  _GEN_1930 = way1_hit ? _GEN_1673 : dirty_1_0; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1931 = way1_hit ? _GEN_1674 : dirty_1_1; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1932 = way1_hit ? _GEN_1675 : dirty_1_2; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1933 = way1_hit ? _GEN_1676 : dirty_1_3; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1934 = way1_hit ? _GEN_1677 : dirty_1_4; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1935 = way1_hit ? _GEN_1678 : dirty_1_5; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1936 = way1_hit ? _GEN_1679 : dirty_1_6; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1937 = way1_hit ? _GEN_1680 : dirty_1_7; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1938 = way1_hit ? _GEN_1681 : dirty_1_8; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1939 = way1_hit ? _GEN_1682 : dirty_1_9; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1940 = way1_hit ? _GEN_1683 : dirty_1_10; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1941 = way1_hit ? _GEN_1684 : dirty_1_11; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1942 = way1_hit ? _GEN_1685 : dirty_1_12; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1943 = way1_hit ? _GEN_1686 : dirty_1_13; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1944 = way1_hit ? _GEN_1687 : dirty_1_14; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1945 = way1_hit ? _GEN_1688 : dirty_1_15; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1946 = way1_hit ? _GEN_1689 : dirty_1_16; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1947 = way1_hit ? _GEN_1690 : dirty_1_17; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1948 = way1_hit ? _GEN_1691 : dirty_1_18; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1949 = way1_hit ? _GEN_1692 : dirty_1_19; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1950 = way1_hit ? _GEN_1693 : dirty_1_20; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1951 = way1_hit ? _GEN_1694 : dirty_1_21; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1952 = way1_hit ? _GEN_1695 : dirty_1_22; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1953 = way1_hit ? _GEN_1696 : dirty_1_23; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1954 = way1_hit ? _GEN_1697 : dirty_1_24; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1955 = way1_hit ? _GEN_1698 : dirty_1_25; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1956 = way1_hit ? _GEN_1699 : dirty_1_26; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1957 = way1_hit ? _GEN_1700 : dirty_1_27; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1958 = way1_hit ? _GEN_1701 : dirty_1_28; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1959 = way1_hit ? _GEN_1702 : dirty_1_29; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1960 = way1_hit ? _GEN_1703 : dirty_1_30; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1961 = way1_hit ? _GEN_1704 : dirty_1_31; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1962 = way1_hit ? _GEN_1705 : dirty_1_32; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1963 = way1_hit ? _GEN_1706 : dirty_1_33; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1964 = way1_hit ? _GEN_1707 : dirty_1_34; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1965 = way1_hit ? _GEN_1708 : dirty_1_35; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1966 = way1_hit ? _GEN_1709 : dirty_1_36; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1967 = way1_hit ? _GEN_1710 : dirty_1_37; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1968 = way1_hit ? _GEN_1711 : dirty_1_38; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1969 = way1_hit ? _GEN_1712 : dirty_1_39; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1970 = way1_hit ? _GEN_1713 : dirty_1_40; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1971 = way1_hit ? _GEN_1714 : dirty_1_41; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1972 = way1_hit ? _GEN_1715 : dirty_1_42; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1973 = way1_hit ? _GEN_1716 : dirty_1_43; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1974 = way1_hit ? _GEN_1717 : dirty_1_44; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1975 = way1_hit ? _GEN_1718 : dirty_1_45; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1976 = way1_hit ? _GEN_1719 : dirty_1_46; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1977 = way1_hit ? _GEN_1720 : dirty_1_47; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1978 = way1_hit ? _GEN_1721 : dirty_1_48; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1979 = way1_hit ? _GEN_1722 : dirty_1_49; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1980 = way1_hit ? _GEN_1723 : dirty_1_50; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1981 = way1_hit ? _GEN_1724 : dirty_1_51; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1982 = way1_hit ? _GEN_1725 : dirty_1_52; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1983 = way1_hit ? _GEN_1726 : dirty_1_53; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1984 = way1_hit ? _GEN_1727 : dirty_1_54; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1985 = way1_hit ? _GEN_1728 : dirty_1_55; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1986 = way1_hit ? _GEN_1729 : dirty_1_56; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1987 = way1_hit ? _GEN_1730 : dirty_1_57; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1988 = way1_hit ? _GEN_1731 : dirty_1_58; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1989 = way1_hit ? _GEN_1732 : dirty_1_59; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1990 = way1_hit ? _GEN_1733 : dirty_1_60; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1991 = way1_hit ? _GEN_1734 : dirty_1_61; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1992 = way1_hit ? _GEN_1735 : dirty_1_62; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1993 = way1_hit ? _GEN_1736 : dirty_1_63; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1994 = way1_hit ? _GEN_1737 : dirty_1_64; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1995 = way1_hit ? _GEN_1738 : dirty_1_65; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1996 = way1_hit ? _GEN_1739 : dirty_1_66; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1997 = way1_hit ? _GEN_1740 : dirty_1_67; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1998 = way1_hit ? _GEN_1741 : dirty_1_68; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_1999 = way1_hit ? _GEN_1742 : dirty_1_69; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2000 = way1_hit ? _GEN_1743 : dirty_1_70; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2001 = way1_hit ? _GEN_1744 : dirty_1_71; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2002 = way1_hit ? _GEN_1745 : dirty_1_72; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2003 = way1_hit ? _GEN_1746 : dirty_1_73; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2004 = way1_hit ? _GEN_1747 : dirty_1_74; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2005 = way1_hit ? _GEN_1748 : dirty_1_75; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2006 = way1_hit ? _GEN_1749 : dirty_1_76; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2007 = way1_hit ? _GEN_1750 : dirty_1_77; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2008 = way1_hit ? _GEN_1751 : dirty_1_78; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2009 = way1_hit ? _GEN_1752 : dirty_1_79; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2010 = way1_hit ? _GEN_1753 : dirty_1_80; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2011 = way1_hit ? _GEN_1754 : dirty_1_81; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2012 = way1_hit ? _GEN_1755 : dirty_1_82; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2013 = way1_hit ? _GEN_1756 : dirty_1_83; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2014 = way1_hit ? _GEN_1757 : dirty_1_84; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2015 = way1_hit ? _GEN_1758 : dirty_1_85; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2016 = way1_hit ? _GEN_1759 : dirty_1_86; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2017 = way1_hit ? _GEN_1760 : dirty_1_87; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2018 = way1_hit ? _GEN_1761 : dirty_1_88; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2019 = way1_hit ? _GEN_1762 : dirty_1_89; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2020 = way1_hit ? _GEN_1763 : dirty_1_90; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2021 = way1_hit ? _GEN_1764 : dirty_1_91; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2022 = way1_hit ? _GEN_1765 : dirty_1_92; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2023 = way1_hit ? _GEN_1766 : dirty_1_93; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2024 = way1_hit ? _GEN_1767 : dirty_1_94; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2025 = way1_hit ? _GEN_1768 : dirty_1_95; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2026 = way1_hit ? _GEN_1769 : dirty_1_96; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2027 = way1_hit ? _GEN_1770 : dirty_1_97; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2028 = way1_hit ? _GEN_1771 : dirty_1_98; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2029 = way1_hit ? _GEN_1772 : dirty_1_99; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2030 = way1_hit ? _GEN_1773 : dirty_1_100; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2031 = way1_hit ? _GEN_1774 : dirty_1_101; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2032 = way1_hit ? _GEN_1775 : dirty_1_102; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2033 = way1_hit ? _GEN_1776 : dirty_1_103; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2034 = way1_hit ? _GEN_1777 : dirty_1_104; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2035 = way1_hit ? _GEN_1778 : dirty_1_105; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2036 = way1_hit ? _GEN_1779 : dirty_1_106; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2037 = way1_hit ? _GEN_1780 : dirty_1_107; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2038 = way1_hit ? _GEN_1781 : dirty_1_108; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2039 = way1_hit ? _GEN_1782 : dirty_1_109; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2040 = way1_hit ? _GEN_1783 : dirty_1_110; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2041 = way1_hit ? _GEN_1784 : dirty_1_111; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2042 = way1_hit ? _GEN_1785 : dirty_1_112; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2043 = way1_hit ? _GEN_1786 : dirty_1_113; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2044 = way1_hit ? _GEN_1787 : dirty_1_114; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2045 = way1_hit ? _GEN_1788 : dirty_1_115; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2046 = way1_hit ? _GEN_1789 : dirty_1_116; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2047 = way1_hit ? _GEN_1790 : dirty_1_117; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2048 = way1_hit ? _GEN_1791 : dirty_1_118; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2049 = way1_hit ? _GEN_1792 : dirty_1_119; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2050 = way1_hit ? _GEN_1793 : dirty_1_120; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2051 = way1_hit ? _GEN_1794 : dirty_1_121; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2052 = way1_hit ? _GEN_1795 : dirty_1_122; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2053 = way1_hit ? _GEN_1796 : dirty_1_123; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2054 = way1_hit ? _GEN_1797 : dirty_1_124; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2055 = way1_hit ? _GEN_1798 : dirty_1_125; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2056 = way1_hit ? _GEN_1799 : dirty_1_126; // @[d_cache.scala 111:33 25:26]
  wire  _GEN_2057 = way1_hit ? _GEN_1800 : dirty_1_127; // @[d_cache.scala 111:33 25:26]
  wire [2:0] _GEN_2058 = way0_hit ? 3'h0 : _GEN_1801; // @[d_cache.scala 104:27 105:23]
  wire [63:0] _GEN_2059 = way0_hit ? _GEN_1161 : ram_0_0; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2060 = way0_hit ? _GEN_1162 : ram_0_1; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2061 = way0_hit ? _GEN_1163 : ram_0_2; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2062 = way0_hit ? _GEN_1164 : ram_0_3; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2063 = way0_hit ? _GEN_1165 : ram_0_4; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2064 = way0_hit ? _GEN_1166 : ram_0_5; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2065 = way0_hit ? _GEN_1167 : ram_0_6; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2066 = way0_hit ? _GEN_1168 : ram_0_7; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2067 = way0_hit ? _GEN_1169 : ram_0_8; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2068 = way0_hit ? _GEN_1170 : ram_0_9; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2069 = way0_hit ? _GEN_1171 : ram_0_10; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2070 = way0_hit ? _GEN_1172 : ram_0_11; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2071 = way0_hit ? _GEN_1173 : ram_0_12; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2072 = way0_hit ? _GEN_1174 : ram_0_13; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2073 = way0_hit ? _GEN_1175 : ram_0_14; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2074 = way0_hit ? _GEN_1176 : ram_0_15; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2075 = way0_hit ? _GEN_1177 : ram_0_16; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2076 = way0_hit ? _GEN_1178 : ram_0_17; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2077 = way0_hit ? _GEN_1179 : ram_0_18; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2078 = way0_hit ? _GEN_1180 : ram_0_19; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2079 = way0_hit ? _GEN_1181 : ram_0_20; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2080 = way0_hit ? _GEN_1182 : ram_0_21; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2081 = way0_hit ? _GEN_1183 : ram_0_22; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2082 = way0_hit ? _GEN_1184 : ram_0_23; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2083 = way0_hit ? _GEN_1185 : ram_0_24; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2084 = way0_hit ? _GEN_1186 : ram_0_25; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2085 = way0_hit ? _GEN_1187 : ram_0_26; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2086 = way0_hit ? _GEN_1188 : ram_0_27; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2087 = way0_hit ? _GEN_1189 : ram_0_28; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2088 = way0_hit ? _GEN_1190 : ram_0_29; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2089 = way0_hit ? _GEN_1191 : ram_0_30; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2090 = way0_hit ? _GEN_1192 : ram_0_31; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2091 = way0_hit ? _GEN_1193 : ram_0_32; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2092 = way0_hit ? _GEN_1194 : ram_0_33; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2093 = way0_hit ? _GEN_1195 : ram_0_34; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2094 = way0_hit ? _GEN_1196 : ram_0_35; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2095 = way0_hit ? _GEN_1197 : ram_0_36; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2096 = way0_hit ? _GEN_1198 : ram_0_37; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2097 = way0_hit ? _GEN_1199 : ram_0_38; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2098 = way0_hit ? _GEN_1200 : ram_0_39; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2099 = way0_hit ? _GEN_1201 : ram_0_40; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2100 = way0_hit ? _GEN_1202 : ram_0_41; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2101 = way0_hit ? _GEN_1203 : ram_0_42; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2102 = way0_hit ? _GEN_1204 : ram_0_43; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2103 = way0_hit ? _GEN_1205 : ram_0_44; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2104 = way0_hit ? _GEN_1206 : ram_0_45; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2105 = way0_hit ? _GEN_1207 : ram_0_46; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2106 = way0_hit ? _GEN_1208 : ram_0_47; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2107 = way0_hit ? _GEN_1209 : ram_0_48; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2108 = way0_hit ? _GEN_1210 : ram_0_49; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2109 = way0_hit ? _GEN_1211 : ram_0_50; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2110 = way0_hit ? _GEN_1212 : ram_0_51; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2111 = way0_hit ? _GEN_1213 : ram_0_52; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2112 = way0_hit ? _GEN_1214 : ram_0_53; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2113 = way0_hit ? _GEN_1215 : ram_0_54; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2114 = way0_hit ? _GEN_1216 : ram_0_55; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2115 = way0_hit ? _GEN_1217 : ram_0_56; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2116 = way0_hit ? _GEN_1218 : ram_0_57; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2117 = way0_hit ? _GEN_1219 : ram_0_58; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2118 = way0_hit ? _GEN_1220 : ram_0_59; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2119 = way0_hit ? _GEN_1221 : ram_0_60; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2120 = way0_hit ? _GEN_1222 : ram_0_61; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2121 = way0_hit ? _GEN_1223 : ram_0_62; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2122 = way0_hit ? _GEN_1224 : ram_0_63; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2123 = way0_hit ? _GEN_1225 : ram_0_64; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2124 = way0_hit ? _GEN_1226 : ram_0_65; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2125 = way0_hit ? _GEN_1227 : ram_0_66; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2126 = way0_hit ? _GEN_1228 : ram_0_67; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2127 = way0_hit ? _GEN_1229 : ram_0_68; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2128 = way0_hit ? _GEN_1230 : ram_0_69; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2129 = way0_hit ? _GEN_1231 : ram_0_70; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2130 = way0_hit ? _GEN_1232 : ram_0_71; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2131 = way0_hit ? _GEN_1233 : ram_0_72; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2132 = way0_hit ? _GEN_1234 : ram_0_73; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2133 = way0_hit ? _GEN_1235 : ram_0_74; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2134 = way0_hit ? _GEN_1236 : ram_0_75; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2135 = way0_hit ? _GEN_1237 : ram_0_76; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2136 = way0_hit ? _GEN_1238 : ram_0_77; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2137 = way0_hit ? _GEN_1239 : ram_0_78; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2138 = way0_hit ? _GEN_1240 : ram_0_79; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2139 = way0_hit ? _GEN_1241 : ram_0_80; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2140 = way0_hit ? _GEN_1242 : ram_0_81; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2141 = way0_hit ? _GEN_1243 : ram_0_82; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2142 = way0_hit ? _GEN_1244 : ram_0_83; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2143 = way0_hit ? _GEN_1245 : ram_0_84; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2144 = way0_hit ? _GEN_1246 : ram_0_85; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2145 = way0_hit ? _GEN_1247 : ram_0_86; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2146 = way0_hit ? _GEN_1248 : ram_0_87; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2147 = way0_hit ? _GEN_1249 : ram_0_88; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2148 = way0_hit ? _GEN_1250 : ram_0_89; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2149 = way0_hit ? _GEN_1251 : ram_0_90; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2150 = way0_hit ? _GEN_1252 : ram_0_91; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2151 = way0_hit ? _GEN_1253 : ram_0_92; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2152 = way0_hit ? _GEN_1254 : ram_0_93; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2153 = way0_hit ? _GEN_1255 : ram_0_94; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2154 = way0_hit ? _GEN_1256 : ram_0_95; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2155 = way0_hit ? _GEN_1257 : ram_0_96; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2156 = way0_hit ? _GEN_1258 : ram_0_97; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2157 = way0_hit ? _GEN_1259 : ram_0_98; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2158 = way0_hit ? _GEN_1260 : ram_0_99; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2159 = way0_hit ? _GEN_1261 : ram_0_100; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2160 = way0_hit ? _GEN_1262 : ram_0_101; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2161 = way0_hit ? _GEN_1263 : ram_0_102; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2162 = way0_hit ? _GEN_1264 : ram_0_103; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2163 = way0_hit ? _GEN_1265 : ram_0_104; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2164 = way0_hit ? _GEN_1266 : ram_0_105; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2165 = way0_hit ? _GEN_1267 : ram_0_106; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2166 = way0_hit ? _GEN_1268 : ram_0_107; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2167 = way0_hit ? _GEN_1269 : ram_0_108; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2168 = way0_hit ? _GEN_1270 : ram_0_109; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2169 = way0_hit ? _GEN_1271 : ram_0_110; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2170 = way0_hit ? _GEN_1272 : ram_0_111; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2171 = way0_hit ? _GEN_1273 : ram_0_112; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2172 = way0_hit ? _GEN_1274 : ram_0_113; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2173 = way0_hit ? _GEN_1275 : ram_0_114; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2174 = way0_hit ? _GEN_1276 : ram_0_115; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2175 = way0_hit ? _GEN_1277 : ram_0_116; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2176 = way0_hit ? _GEN_1278 : ram_0_117; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2177 = way0_hit ? _GEN_1279 : ram_0_118; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2178 = way0_hit ? _GEN_1280 : ram_0_119; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2179 = way0_hit ? _GEN_1281 : ram_0_120; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2180 = way0_hit ? _GEN_1282 : ram_0_121; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2181 = way0_hit ? _GEN_1283 : ram_0_122; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2182 = way0_hit ? _GEN_1284 : ram_0_123; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2183 = way0_hit ? _GEN_1285 : ram_0_124; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2184 = way0_hit ? _GEN_1286 : ram_0_125; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2185 = way0_hit ? _GEN_1287 : ram_0_126; // @[d_cache.scala 104:27 18:24]
  wire [63:0] _GEN_2186 = way0_hit ? _GEN_1288 : ram_0_127; // @[d_cache.scala 104:27 18:24]
  wire  _GEN_2187 = way0_hit ? _GEN_1289 : dirty_0_0; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2188 = way0_hit ? _GEN_1290 : dirty_0_1; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2189 = way0_hit ? _GEN_1291 : dirty_0_2; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2190 = way0_hit ? _GEN_1292 : dirty_0_3; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2191 = way0_hit ? _GEN_1293 : dirty_0_4; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2192 = way0_hit ? _GEN_1294 : dirty_0_5; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2193 = way0_hit ? _GEN_1295 : dirty_0_6; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2194 = way0_hit ? _GEN_1296 : dirty_0_7; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2195 = way0_hit ? _GEN_1297 : dirty_0_8; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2196 = way0_hit ? _GEN_1298 : dirty_0_9; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2197 = way0_hit ? _GEN_1299 : dirty_0_10; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2198 = way0_hit ? _GEN_1300 : dirty_0_11; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2199 = way0_hit ? _GEN_1301 : dirty_0_12; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2200 = way0_hit ? _GEN_1302 : dirty_0_13; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2201 = way0_hit ? _GEN_1303 : dirty_0_14; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2202 = way0_hit ? _GEN_1304 : dirty_0_15; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2203 = way0_hit ? _GEN_1305 : dirty_0_16; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2204 = way0_hit ? _GEN_1306 : dirty_0_17; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2205 = way0_hit ? _GEN_1307 : dirty_0_18; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2206 = way0_hit ? _GEN_1308 : dirty_0_19; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2207 = way0_hit ? _GEN_1309 : dirty_0_20; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2208 = way0_hit ? _GEN_1310 : dirty_0_21; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2209 = way0_hit ? _GEN_1311 : dirty_0_22; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2210 = way0_hit ? _GEN_1312 : dirty_0_23; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2211 = way0_hit ? _GEN_1313 : dirty_0_24; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2212 = way0_hit ? _GEN_1314 : dirty_0_25; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2213 = way0_hit ? _GEN_1315 : dirty_0_26; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2214 = way0_hit ? _GEN_1316 : dirty_0_27; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2215 = way0_hit ? _GEN_1317 : dirty_0_28; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2216 = way0_hit ? _GEN_1318 : dirty_0_29; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2217 = way0_hit ? _GEN_1319 : dirty_0_30; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2218 = way0_hit ? _GEN_1320 : dirty_0_31; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2219 = way0_hit ? _GEN_1321 : dirty_0_32; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2220 = way0_hit ? _GEN_1322 : dirty_0_33; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2221 = way0_hit ? _GEN_1323 : dirty_0_34; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2222 = way0_hit ? _GEN_1324 : dirty_0_35; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2223 = way0_hit ? _GEN_1325 : dirty_0_36; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2224 = way0_hit ? _GEN_1326 : dirty_0_37; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2225 = way0_hit ? _GEN_1327 : dirty_0_38; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2226 = way0_hit ? _GEN_1328 : dirty_0_39; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2227 = way0_hit ? _GEN_1329 : dirty_0_40; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2228 = way0_hit ? _GEN_1330 : dirty_0_41; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2229 = way0_hit ? _GEN_1331 : dirty_0_42; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2230 = way0_hit ? _GEN_1332 : dirty_0_43; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2231 = way0_hit ? _GEN_1333 : dirty_0_44; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2232 = way0_hit ? _GEN_1334 : dirty_0_45; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2233 = way0_hit ? _GEN_1335 : dirty_0_46; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2234 = way0_hit ? _GEN_1336 : dirty_0_47; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2235 = way0_hit ? _GEN_1337 : dirty_0_48; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2236 = way0_hit ? _GEN_1338 : dirty_0_49; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2237 = way0_hit ? _GEN_1339 : dirty_0_50; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2238 = way0_hit ? _GEN_1340 : dirty_0_51; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2239 = way0_hit ? _GEN_1341 : dirty_0_52; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2240 = way0_hit ? _GEN_1342 : dirty_0_53; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2241 = way0_hit ? _GEN_1343 : dirty_0_54; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2242 = way0_hit ? _GEN_1344 : dirty_0_55; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2243 = way0_hit ? _GEN_1345 : dirty_0_56; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2244 = way0_hit ? _GEN_1346 : dirty_0_57; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2245 = way0_hit ? _GEN_1347 : dirty_0_58; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2246 = way0_hit ? _GEN_1348 : dirty_0_59; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2247 = way0_hit ? _GEN_1349 : dirty_0_60; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2248 = way0_hit ? _GEN_1350 : dirty_0_61; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2249 = way0_hit ? _GEN_1351 : dirty_0_62; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2250 = way0_hit ? _GEN_1352 : dirty_0_63; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2251 = way0_hit ? _GEN_1353 : dirty_0_64; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2252 = way0_hit ? _GEN_1354 : dirty_0_65; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2253 = way0_hit ? _GEN_1355 : dirty_0_66; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2254 = way0_hit ? _GEN_1356 : dirty_0_67; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2255 = way0_hit ? _GEN_1357 : dirty_0_68; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2256 = way0_hit ? _GEN_1358 : dirty_0_69; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2257 = way0_hit ? _GEN_1359 : dirty_0_70; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2258 = way0_hit ? _GEN_1360 : dirty_0_71; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2259 = way0_hit ? _GEN_1361 : dirty_0_72; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2260 = way0_hit ? _GEN_1362 : dirty_0_73; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2261 = way0_hit ? _GEN_1363 : dirty_0_74; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2262 = way0_hit ? _GEN_1364 : dirty_0_75; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2263 = way0_hit ? _GEN_1365 : dirty_0_76; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2264 = way0_hit ? _GEN_1366 : dirty_0_77; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2265 = way0_hit ? _GEN_1367 : dirty_0_78; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2266 = way0_hit ? _GEN_1368 : dirty_0_79; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2267 = way0_hit ? _GEN_1369 : dirty_0_80; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2268 = way0_hit ? _GEN_1370 : dirty_0_81; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2269 = way0_hit ? _GEN_1371 : dirty_0_82; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2270 = way0_hit ? _GEN_1372 : dirty_0_83; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2271 = way0_hit ? _GEN_1373 : dirty_0_84; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2272 = way0_hit ? _GEN_1374 : dirty_0_85; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2273 = way0_hit ? _GEN_1375 : dirty_0_86; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2274 = way0_hit ? _GEN_1376 : dirty_0_87; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2275 = way0_hit ? _GEN_1377 : dirty_0_88; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2276 = way0_hit ? _GEN_1378 : dirty_0_89; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2277 = way0_hit ? _GEN_1379 : dirty_0_90; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2278 = way0_hit ? _GEN_1380 : dirty_0_91; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2279 = way0_hit ? _GEN_1381 : dirty_0_92; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2280 = way0_hit ? _GEN_1382 : dirty_0_93; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2281 = way0_hit ? _GEN_1383 : dirty_0_94; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2282 = way0_hit ? _GEN_1384 : dirty_0_95; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2283 = way0_hit ? _GEN_1385 : dirty_0_96; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2284 = way0_hit ? _GEN_1386 : dirty_0_97; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2285 = way0_hit ? _GEN_1387 : dirty_0_98; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2286 = way0_hit ? _GEN_1388 : dirty_0_99; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2287 = way0_hit ? _GEN_1389 : dirty_0_100; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2288 = way0_hit ? _GEN_1390 : dirty_0_101; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2289 = way0_hit ? _GEN_1391 : dirty_0_102; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2290 = way0_hit ? _GEN_1392 : dirty_0_103; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2291 = way0_hit ? _GEN_1393 : dirty_0_104; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2292 = way0_hit ? _GEN_1394 : dirty_0_105; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2293 = way0_hit ? _GEN_1395 : dirty_0_106; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2294 = way0_hit ? _GEN_1396 : dirty_0_107; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2295 = way0_hit ? _GEN_1397 : dirty_0_108; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2296 = way0_hit ? _GEN_1398 : dirty_0_109; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2297 = way0_hit ? _GEN_1399 : dirty_0_110; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2298 = way0_hit ? _GEN_1400 : dirty_0_111; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2299 = way0_hit ? _GEN_1401 : dirty_0_112; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2300 = way0_hit ? _GEN_1402 : dirty_0_113; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2301 = way0_hit ? _GEN_1403 : dirty_0_114; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2302 = way0_hit ? _GEN_1404 : dirty_0_115; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2303 = way0_hit ? _GEN_1405 : dirty_0_116; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2304 = way0_hit ? _GEN_1406 : dirty_0_117; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2305 = way0_hit ? _GEN_1407 : dirty_0_118; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2306 = way0_hit ? _GEN_1408 : dirty_0_119; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2307 = way0_hit ? _GEN_1409 : dirty_0_120; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2308 = way0_hit ? _GEN_1410 : dirty_0_121; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2309 = way0_hit ? _GEN_1411 : dirty_0_122; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2310 = way0_hit ? _GEN_1412 : dirty_0_123; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2311 = way0_hit ? _GEN_1413 : dirty_0_124; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2312 = way0_hit ? _GEN_1414 : dirty_0_125; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2313 = way0_hit ? _GEN_1415 : dirty_0_126; // @[d_cache.scala 104:27 24:26]
  wire  _GEN_2314 = way0_hit ? _GEN_1416 : dirty_0_127; // @[d_cache.scala 104:27 24:26]
  wire [63:0] _GEN_2315 = way0_hit ? ram_1_0 : _GEN_1802; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2316 = way0_hit ? ram_1_1 : _GEN_1803; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2317 = way0_hit ? ram_1_2 : _GEN_1804; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2318 = way0_hit ? ram_1_3 : _GEN_1805; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2319 = way0_hit ? ram_1_4 : _GEN_1806; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2320 = way0_hit ? ram_1_5 : _GEN_1807; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2321 = way0_hit ? ram_1_6 : _GEN_1808; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2322 = way0_hit ? ram_1_7 : _GEN_1809; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2323 = way0_hit ? ram_1_8 : _GEN_1810; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2324 = way0_hit ? ram_1_9 : _GEN_1811; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2325 = way0_hit ? ram_1_10 : _GEN_1812; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2326 = way0_hit ? ram_1_11 : _GEN_1813; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2327 = way0_hit ? ram_1_12 : _GEN_1814; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2328 = way0_hit ? ram_1_13 : _GEN_1815; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2329 = way0_hit ? ram_1_14 : _GEN_1816; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2330 = way0_hit ? ram_1_15 : _GEN_1817; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2331 = way0_hit ? ram_1_16 : _GEN_1818; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2332 = way0_hit ? ram_1_17 : _GEN_1819; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2333 = way0_hit ? ram_1_18 : _GEN_1820; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2334 = way0_hit ? ram_1_19 : _GEN_1821; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2335 = way0_hit ? ram_1_20 : _GEN_1822; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2336 = way0_hit ? ram_1_21 : _GEN_1823; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2337 = way0_hit ? ram_1_22 : _GEN_1824; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2338 = way0_hit ? ram_1_23 : _GEN_1825; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2339 = way0_hit ? ram_1_24 : _GEN_1826; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2340 = way0_hit ? ram_1_25 : _GEN_1827; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2341 = way0_hit ? ram_1_26 : _GEN_1828; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2342 = way0_hit ? ram_1_27 : _GEN_1829; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2343 = way0_hit ? ram_1_28 : _GEN_1830; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2344 = way0_hit ? ram_1_29 : _GEN_1831; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2345 = way0_hit ? ram_1_30 : _GEN_1832; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2346 = way0_hit ? ram_1_31 : _GEN_1833; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2347 = way0_hit ? ram_1_32 : _GEN_1834; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2348 = way0_hit ? ram_1_33 : _GEN_1835; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2349 = way0_hit ? ram_1_34 : _GEN_1836; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2350 = way0_hit ? ram_1_35 : _GEN_1837; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2351 = way0_hit ? ram_1_36 : _GEN_1838; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2352 = way0_hit ? ram_1_37 : _GEN_1839; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2353 = way0_hit ? ram_1_38 : _GEN_1840; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2354 = way0_hit ? ram_1_39 : _GEN_1841; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2355 = way0_hit ? ram_1_40 : _GEN_1842; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2356 = way0_hit ? ram_1_41 : _GEN_1843; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2357 = way0_hit ? ram_1_42 : _GEN_1844; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2358 = way0_hit ? ram_1_43 : _GEN_1845; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2359 = way0_hit ? ram_1_44 : _GEN_1846; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2360 = way0_hit ? ram_1_45 : _GEN_1847; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2361 = way0_hit ? ram_1_46 : _GEN_1848; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2362 = way0_hit ? ram_1_47 : _GEN_1849; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2363 = way0_hit ? ram_1_48 : _GEN_1850; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2364 = way0_hit ? ram_1_49 : _GEN_1851; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2365 = way0_hit ? ram_1_50 : _GEN_1852; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2366 = way0_hit ? ram_1_51 : _GEN_1853; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2367 = way0_hit ? ram_1_52 : _GEN_1854; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2368 = way0_hit ? ram_1_53 : _GEN_1855; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2369 = way0_hit ? ram_1_54 : _GEN_1856; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2370 = way0_hit ? ram_1_55 : _GEN_1857; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2371 = way0_hit ? ram_1_56 : _GEN_1858; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2372 = way0_hit ? ram_1_57 : _GEN_1859; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2373 = way0_hit ? ram_1_58 : _GEN_1860; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2374 = way0_hit ? ram_1_59 : _GEN_1861; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2375 = way0_hit ? ram_1_60 : _GEN_1862; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2376 = way0_hit ? ram_1_61 : _GEN_1863; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2377 = way0_hit ? ram_1_62 : _GEN_1864; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2378 = way0_hit ? ram_1_63 : _GEN_1865; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2379 = way0_hit ? ram_1_64 : _GEN_1866; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2380 = way0_hit ? ram_1_65 : _GEN_1867; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2381 = way0_hit ? ram_1_66 : _GEN_1868; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2382 = way0_hit ? ram_1_67 : _GEN_1869; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2383 = way0_hit ? ram_1_68 : _GEN_1870; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2384 = way0_hit ? ram_1_69 : _GEN_1871; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2385 = way0_hit ? ram_1_70 : _GEN_1872; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2386 = way0_hit ? ram_1_71 : _GEN_1873; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2387 = way0_hit ? ram_1_72 : _GEN_1874; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2388 = way0_hit ? ram_1_73 : _GEN_1875; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2389 = way0_hit ? ram_1_74 : _GEN_1876; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2390 = way0_hit ? ram_1_75 : _GEN_1877; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2391 = way0_hit ? ram_1_76 : _GEN_1878; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2392 = way0_hit ? ram_1_77 : _GEN_1879; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2393 = way0_hit ? ram_1_78 : _GEN_1880; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2394 = way0_hit ? ram_1_79 : _GEN_1881; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2395 = way0_hit ? ram_1_80 : _GEN_1882; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2396 = way0_hit ? ram_1_81 : _GEN_1883; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2397 = way0_hit ? ram_1_82 : _GEN_1884; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2398 = way0_hit ? ram_1_83 : _GEN_1885; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2399 = way0_hit ? ram_1_84 : _GEN_1886; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2400 = way0_hit ? ram_1_85 : _GEN_1887; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2401 = way0_hit ? ram_1_86 : _GEN_1888; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2402 = way0_hit ? ram_1_87 : _GEN_1889; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2403 = way0_hit ? ram_1_88 : _GEN_1890; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2404 = way0_hit ? ram_1_89 : _GEN_1891; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2405 = way0_hit ? ram_1_90 : _GEN_1892; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2406 = way0_hit ? ram_1_91 : _GEN_1893; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2407 = way0_hit ? ram_1_92 : _GEN_1894; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2408 = way0_hit ? ram_1_93 : _GEN_1895; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2409 = way0_hit ? ram_1_94 : _GEN_1896; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2410 = way0_hit ? ram_1_95 : _GEN_1897; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2411 = way0_hit ? ram_1_96 : _GEN_1898; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2412 = way0_hit ? ram_1_97 : _GEN_1899; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2413 = way0_hit ? ram_1_98 : _GEN_1900; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2414 = way0_hit ? ram_1_99 : _GEN_1901; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2415 = way0_hit ? ram_1_100 : _GEN_1902; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2416 = way0_hit ? ram_1_101 : _GEN_1903; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2417 = way0_hit ? ram_1_102 : _GEN_1904; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2418 = way0_hit ? ram_1_103 : _GEN_1905; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2419 = way0_hit ? ram_1_104 : _GEN_1906; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2420 = way0_hit ? ram_1_105 : _GEN_1907; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2421 = way0_hit ? ram_1_106 : _GEN_1908; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2422 = way0_hit ? ram_1_107 : _GEN_1909; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2423 = way0_hit ? ram_1_108 : _GEN_1910; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2424 = way0_hit ? ram_1_109 : _GEN_1911; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2425 = way0_hit ? ram_1_110 : _GEN_1912; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2426 = way0_hit ? ram_1_111 : _GEN_1913; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2427 = way0_hit ? ram_1_112 : _GEN_1914; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2428 = way0_hit ? ram_1_113 : _GEN_1915; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2429 = way0_hit ? ram_1_114 : _GEN_1916; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2430 = way0_hit ? ram_1_115 : _GEN_1917; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2431 = way0_hit ? ram_1_116 : _GEN_1918; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2432 = way0_hit ? ram_1_117 : _GEN_1919; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2433 = way0_hit ? ram_1_118 : _GEN_1920; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2434 = way0_hit ? ram_1_119 : _GEN_1921; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2435 = way0_hit ? ram_1_120 : _GEN_1922; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2436 = way0_hit ? ram_1_121 : _GEN_1923; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2437 = way0_hit ? ram_1_122 : _GEN_1924; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2438 = way0_hit ? ram_1_123 : _GEN_1925; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2439 = way0_hit ? ram_1_124 : _GEN_1926; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2440 = way0_hit ? ram_1_125 : _GEN_1927; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2441 = way0_hit ? ram_1_126 : _GEN_1928; // @[d_cache.scala 104:27 19:24]
  wire [63:0] _GEN_2442 = way0_hit ? ram_1_127 : _GEN_1929; // @[d_cache.scala 104:27 19:24]
  wire  _GEN_2443 = way0_hit ? dirty_1_0 : _GEN_1930; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2444 = way0_hit ? dirty_1_1 : _GEN_1931; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2445 = way0_hit ? dirty_1_2 : _GEN_1932; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2446 = way0_hit ? dirty_1_3 : _GEN_1933; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2447 = way0_hit ? dirty_1_4 : _GEN_1934; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2448 = way0_hit ? dirty_1_5 : _GEN_1935; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2449 = way0_hit ? dirty_1_6 : _GEN_1936; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2450 = way0_hit ? dirty_1_7 : _GEN_1937; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2451 = way0_hit ? dirty_1_8 : _GEN_1938; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2452 = way0_hit ? dirty_1_9 : _GEN_1939; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2453 = way0_hit ? dirty_1_10 : _GEN_1940; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2454 = way0_hit ? dirty_1_11 : _GEN_1941; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2455 = way0_hit ? dirty_1_12 : _GEN_1942; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2456 = way0_hit ? dirty_1_13 : _GEN_1943; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2457 = way0_hit ? dirty_1_14 : _GEN_1944; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2458 = way0_hit ? dirty_1_15 : _GEN_1945; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2459 = way0_hit ? dirty_1_16 : _GEN_1946; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2460 = way0_hit ? dirty_1_17 : _GEN_1947; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2461 = way0_hit ? dirty_1_18 : _GEN_1948; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2462 = way0_hit ? dirty_1_19 : _GEN_1949; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2463 = way0_hit ? dirty_1_20 : _GEN_1950; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2464 = way0_hit ? dirty_1_21 : _GEN_1951; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2465 = way0_hit ? dirty_1_22 : _GEN_1952; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2466 = way0_hit ? dirty_1_23 : _GEN_1953; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2467 = way0_hit ? dirty_1_24 : _GEN_1954; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2468 = way0_hit ? dirty_1_25 : _GEN_1955; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2469 = way0_hit ? dirty_1_26 : _GEN_1956; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2470 = way0_hit ? dirty_1_27 : _GEN_1957; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2471 = way0_hit ? dirty_1_28 : _GEN_1958; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2472 = way0_hit ? dirty_1_29 : _GEN_1959; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2473 = way0_hit ? dirty_1_30 : _GEN_1960; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2474 = way0_hit ? dirty_1_31 : _GEN_1961; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2475 = way0_hit ? dirty_1_32 : _GEN_1962; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2476 = way0_hit ? dirty_1_33 : _GEN_1963; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2477 = way0_hit ? dirty_1_34 : _GEN_1964; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2478 = way0_hit ? dirty_1_35 : _GEN_1965; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2479 = way0_hit ? dirty_1_36 : _GEN_1966; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2480 = way0_hit ? dirty_1_37 : _GEN_1967; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2481 = way0_hit ? dirty_1_38 : _GEN_1968; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2482 = way0_hit ? dirty_1_39 : _GEN_1969; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2483 = way0_hit ? dirty_1_40 : _GEN_1970; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2484 = way0_hit ? dirty_1_41 : _GEN_1971; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2485 = way0_hit ? dirty_1_42 : _GEN_1972; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2486 = way0_hit ? dirty_1_43 : _GEN_1973; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2487 = way0_hit ? dirty_1_44 : _GEN_1974; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2488 = way0_hit ? dirty_1_45 : _GEN_1975; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2489 = way0_hit ? dirty_1_46 : _GEN_1976; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2490 = way0_hit ? dirty_1_47 : _GEN_1977; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2491 = way0_hit ? dirty_1_48 : _GEN_1978; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2492 = way0_hit ? dirty_1_49 : _GEN_1979; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2493 = way0_hit ? dirty_1_50 : _GEN_1980; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2494 = way0_hit ? dirty_1_51 : _GEN_1981; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2495 = way0_hit ? dirty_1_52 : _GEN_1982; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2496 = way0_hit ? dirty_1_53 : _GEN_1983; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2497 = way0_hit ? dirty_1_54 : _GEN_1984; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2498 = way0_hit ? dirty_1_55 : _GEN_1985; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2499 = way0_hit ? dirty_1_56 : _GEN_1986; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2500 = way0_hit ? dirty_1_57 : _GEN_1987; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2501 = way0_hit ? dirty_1_58 : _GEN_1988; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2502 = way0_hit ? dirty_1_59 : _GEN_1989; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2503 = way0_hit ? dirty_1_60 : _GEN_1990; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2504 = way0_hit ? dirty_1_61 : _GEN_1991; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2505 = way0_hit ? dirty_1_62 : _GEN_1992; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2506 = way0_hit ? dirty_1_63 : _GEN_1993; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2507 = way0_hit ? dirty_1_64 : _GEN_1994; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2508 = way0_hit ? dirty_1_65 : _GEN_1995; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2509 = way0_hit ? dirty_1_66 : _GEN_1996; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2510 = way0_hit ? dirty_1_67 : _GEN_1997; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2511 = way0_hit ? dirty_1_68 : _GEN_1998; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2512 = way0_hit ? dirty_1_69 : _GEN_1999; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2513 = way0_hit ? dirty_1_70 : _GEN_2000; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2514 = way0_hit ? dirty_1_71 : _GEN_2001; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2515 = way0_hit ? dirty_1_72 : _GEN_2002; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2516 = way0_hit ? dirty_1_73 : _GEN_2003; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2517 = way0_hit ? dirty_1_74 : _GEN_2004; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2518 = way0_hit ? dirty_1_75 : _GEN_2005; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2519 = way0_hit ? dirty_1_76 : _GEN_2006; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2520 = way0_hit ? dirty_1_77 : _GEN_2007; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2521 = way0_hit ? dirty_1_78 : _GEN_2008; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2522 = way0_hit ? dirty_1_79 : _GEN_2009; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2523 = way0_hit ? dirty_1_80 : _GEN_2010; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2524 = way0_hit ? dirty_1_81 : _GEN_2011; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2525 = way0_hit ? dirty_1_82 : _GEN_2012; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2526 = way0_hit ? dirty_1_83 : _GEN_2013; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2527 = way0_hit ? dirty_1_84 : _GEN_2014; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2528 = way0_hit ? dirty_1_85 : _GEN_2015; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2529 = way0_hit ? dirty_1_86 : _GEN_2016; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2530 = way0_hit ? dirty_1_87 : _GEN_2017; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2531 = way0_hit ? dirty_1_88 : _GEN_2018; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2532 = way0_hit ? dirty_1_89 : _GEN_2019; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2533 = way0_hit ? dirty_1_90 : _GEN_2020; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2534 = way0_hit ? dirty_1_91 : _GEN_2021; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2535 = way0_hit ? dirty_1_92 : _GEN_2022; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2536 = way0_hit ? dirty_1_93 : _GEN_2023; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2537 = way0_hit ? dirty_1_94 : _GEN_2024; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2538 = way0_hit ? dirty_1_95 : _GEN_2025; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2539 = way0_hit ? dirty_1_96 : _GEN_2026; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2540 = way0_hit ? dirty_1_97 : _GEN_2027; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2541 = way0_hit ? dirty_1_98 : _GEN_2028; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2542 = way0_hit ? dirty_1_99 : _GEN_2029; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2543 = way0_hit ? dirty_1_100 : _GEN_2030; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2544 = way0_hit ? dirty_1_101 : _GEN_2031; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2545 = way0_hit ? dirty_1_102 : _GEN_2032; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2546 = way0_hit ? dirty_1_103 : _GEN_2033; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2547 = way0_hit ? dirty_1_104 : _GEN_2034; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2548 = way0_hit ? dirty_1_105 : _GEN_2035; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2549 = way0_hit ? dirty_1_106 : _GEN_2036; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2550 = way0_hit ? dirty_1_107 : _GEN_2037; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2551 = way0_hit ? dirty_1_108 : _GEN_2038; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2552 = way0_hit ? dirty_1_109 : _GEN_2039; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2553 = way0_hit ? dirty_1_110 : _GEN_2040; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2554 = way0_hit ? dirty_1_111 : _GEN_2041; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2555 = way0_hit ? dirty_1_112 : _GEN_2042; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2556 = way0_hit ? dirty_1_113 : _GEN_2043; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2557 = way0_hit ? dirty_1_114 : _GEN_2044; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2558 = way0_hit ? dirty_1_115 : _GEN_2045; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2559 = way0_hit ? dirty_1_116 : _GEN_2046; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2560 = way0_hit ? dirty_1_117 : _GEN_2047; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2561 = way0_hit ? dirty_1_118 : _GEN_2048; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2562 = way0_hit ? dirty_1_119 : _GEN_2049; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2563 = way0_hit ? dirty_1_120 : _GEN_2050; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2564 = way0_hit ? dirty_1_121 : _GEN_2051; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2565 = way0_hit ? dirty_1_122 : _GEN_2052; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2566 = way0_hit ? dirty_1_123 : _GEN_2053; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2567 = way0_hit ? dirty_1_124 : _GEN_2054; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2568 = way0_hit ? dirty_1_125 : _GEN_2055; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2569 = way0_hit ? dirty_1_126 : _GEN_2056; // @[d_cache.scala 104:27 25:26]
  wire  _GEN_2570 = way0_hit ? dirty_1_127 : _GEN_2057; // @[d_cache.scala 104:27 25:26]
  wire [2:0] _GEN_2571 = io_from_axi_rvalid ? 3'h5 : state; // @[d_cache.scala 121:37 122:23 73:24]
  wire [63:0] _GEN_2572 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[d_cache.scala 124:37 125:30 34:31]
  wire [2:0] _GEN_2573 = io_from_axi_bvalid ? 3'h0 : state; // @[d_cache.scala 129:37 130:23 73:24]
  wire [63:0] _GEN_2574 = 7'h0 == index[6:0] ? receive_data : ram_0_0; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2575 = 7'h1 == index[6:0] ? receive_data : ram_0_1; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2576 = 7'h2 == index[6:0] ? receive_data : ram_0_2; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2577 = 7'h3 == index[6:0] ? receive_data : ram_0_3; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2578 = 7'h4 == index[6:0] ? receive_data : ram_0_4; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2579 = 7'h5 == index[6:0] ? receive_data : ram_0_5; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2580 = 7'h6 == index[6:0] ? receive_data : ram_0_6; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2581 = 7'h7 == index[6:0] ? receive_data : ram_0_7; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2582 = 7'h8 == index[6:0] ? receive_data : ram_0_8; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2583 = 7'h9 == index[6:0] ? receive_data : ram_0_9; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2584 = 7'ha == index[6:0] ? receive_data : ram_0_10; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2585 = 7'hb == index[6:0] ? receive_data : ram_0_11; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2586 = 7'hc == index[6:0] ? receive_data : ram_0_12; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2587 = 7'hd == index[6:0] ? receive_data : ram_0_13; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2588 = 7'he == index[6:0] ? receive_data : ram_0_14; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2589 = 7'hf == index[6:0] ? receive_data : ram_0_15; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2590 = 7'h10 == index[6:0] ? receive_data : ram_0_16; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2591 = 7'h11 == index[6:0] ? receive_data : ram_0_17; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2592 = 7'h12 == index[6:0] ? receive_data : ram_0_18; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2593 = 7'h13 == index[6:0] ? receive_data : ram_0_19; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2594 = 7'h14 == index[6:0] ? receive_data : ram_0_20; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2595 = 7'h15 == index[6:0] ? receive_data : ram_0_21; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2596 = 7'h16 == index[6:0] ? receive_data : ram_0_22; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2597 = 7'h17 == index[6:0] ? receive_data : ram_0_23; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2598 = 7'h18 == index[6:0] ? receive_data : ram_0_24; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2599 = 7'h19 == index[6:0] ? receive_data : ram_0_25; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2600 = 7'h1a == index[6:0] ? receive_data : ram_0_26; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2601 = 7'h1b == index[6:0] ? receive_data : ram_0_27; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2602 = 7'h1c == index[6:0] ? receive_data : ram_0_28; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2603 = 7'h1d == index[6:0] ? receive_data : ram_0_29; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2604 = 7'h1e == index[6:0] ? receive_data : ram_0_30; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2605 = 7'h1f == index[6:0] ? receive_data : ram_0_31; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2606 = 7'h20 == index[6:0] ? receive_data : ram_0_32; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2607 = 7'h21 == index[6:0] ? receive_data : ram_0_33; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2608 = 7'h22 == index[6:0] ? receive_data : ram_0_34; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2609 = 7'h23 == index[6:0] ? receive_data : ram_0_35; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2610 = 7'h24 == index[6:0] ? receive_data : ram_0_36; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2611 = 7'h25 == index[6:0] ? receive_data : ram_0_37; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2612 = 7'h26 == index[6:0] ? receive_data : ram_0_38; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2613 = 7'h27 == index[6:0] ? receive_data : ram_0_39; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2614 = 7'h28 == index[6:0] ? receive_data : ram_0_40; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2615 = 7'h29 == index[6:0] ? receive_data : ram_0_41; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2616 = 7'h2a == index[6:0] ? receive_data : ram_0_42; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2617 = 7'h2b == index[6:0] ? receive_data : ram_0_43; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2618 = 7'h2c == index[6:0] ? receive_data : ram_0_44; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2619 = 7'h2d == index[6:0] ? receive_data : ram_0_45; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2620 = 7'h2e == index[6:0] ? receive_data : ram_0_46; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2621 = 7'h2f == index[6:0] ? receive_data : ram_0_47; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2622 = 7'h30 == index[6:0] ? receive_data : ram_0_48; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2623 = 7'h31 == index[6:0] ? receive_data : ram_0_49; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2624 = 7'h32 == index[6:0] ? receive_data : ram_0_50; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2625 = 7'h33 == index[6:0] ? receive_data : ram_0_51; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2626 = 7'h34 == index[6:0] ? receive_data : ram_0_52; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2627 = 7'h35 == index[6:0] ? receive_data : ram_0_53; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2628 = 7'h36 == index[6:0] ? receive_data : ram_0_54; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2629 = 7'h37 == index[6:0] ? receive_data : ram_0_55; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2630 = 7'h38 == index[6:0] ? receive_data : ram_0_56; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2631 = 7'h39 == index[6:0] ? receive_data : ram_0_57; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2632 = 7'h3a == index[6:0] ? receive_data : ram_0_58; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2633 = 7'h3b == index[6:0] ? receive_data : ram_0_59; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2634 = 7'h3c == index[6:0] ? receive_data : ram_0_60; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2635 = 7'h3d == index[6:0] ? receive_data : ram_0_61; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2636 = 7'h3e == index[6:0] ? receive_data : ram_0_62; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2637 = 7'h3f == index[6:0] ? receive_data : ram_0_63; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2638 = 7'h40 == index[6:0] ? receive_data : ram_0_64; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2639 = 7'h41 == index[6:0] ? receive_data : ram_0_65; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2640 = 7'h42 == index[6:0] ? receive_data : ram_0_66; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2641 = 7'h43 == index[6:0] ? receive_data : ram_0_67; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2642 = 7'h44 == index[6:0] ? receive_data : ram_0_68; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2643 = 7'h45 == index[6:0] ? receive_data : ram_0_69; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2644 = 7'h46 == index[6:0] ? receive_data : ram_0_70; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2645 = 7'h47 == index[6:0] ? receive_data : ram_0_71; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2646 = 7'h48 == index[6:0] ? receive_data : ram_0_72; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2647 = 7'h49 == index[6:0] ? receive_data : ram_0_73; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2648 = 7'h4a == index[6:0] ? receive_data : ram_0_74; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2649 = 7'h4b == index[6:0] ? receive_data : ram_0_75; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2650 = 7'h4c == index[6:0] ? receive_data : ram_0_76; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2651 = 7'h4d == index[6:0] ? receive_data : ram_0_77; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2652 = 7'h4e == index[6:0] ? receive_data : ram_0_78; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2653 = 7'h4f == index[6:0] ? receive_data : ram_0_79; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2654 = 7'h50 == index[6:0] ? receive_data : ram_0_80; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2655 = 7'h51 == index[6:0] ? receive_data : ram_0_81; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2656 = 7'h52 == index[6:0] ? receive_data : ram_0_82; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2657 = 7'h53 == index[6:0] ? receive_data : ram_0_83; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2658 = 7'h54 == index[6:0] ? receive_data : ram_0_84; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2659 = 7'h55 == index[6:0] ? receive_data : ram_0_85; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2660 = 7'h56 == index[6:0] ? receive_data : ram_0_86; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2661 = 7'h57 == index[6:0] ? receive_data : ram_0_87; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2662 = 7'h58 == index[6:0] ? receive_data : ram_0_88; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2663 = 7'h59 == index[6:0] ? receive_data : ram_0_89; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2664 = 7'h5a == index[6:0] ? receive_data : ram_0_90; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2665 = 7'h5b == index[6:0] ? receive_data : ram_0_91; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2666 = 7'h5c == index[6:0] ? receive_data : ram_0_92; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2667 = 7'h5d == index[6:0] ? receive_data : ram_0_93; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2668 = 7'h5e == index[6:0] ? receive_data : ram_0_94; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2669 = 7'h5f == index[6:0] ? receive_data : ram_0_95; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2670 = 7'h60 == index[6:0] ? receive_data : ram_0_96; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2671 = 7'h61 == index[6:0] ? receive_data : ram_0_97; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2672 = 7'h62 == index[6:0] ? receive_data : ram_0_98; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2673 = 7'h63 == index[6:0] ? receive_data : ram_0_99; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2674 = 7'h64 == index[6:0] ? receive_data : ram_0_100; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2675 = 7'h65 == index[6:0] ? receive_data : ram_0_101; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2676 = 7'h66 == index[6:0] ? receive_data : ram_0_102; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2677 = 7'h67 == index[6:0] ? receive_data : ram_0_103; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2678 = 7'h68 == index[6:0] ? receive_data : ram_0_104; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2679 = 7'h69 == index[6:0] ? receive_data : ram_0_105; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2680 = 7'h6a == index[6:0] ? receive_data : ram_0_106; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2681 = 7'h6b == index[6:0] ? receive_data : ram_0_107; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2682 = 7'h6c == index[6:0] ? receive_data : ram_0_108; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2683 = 7'h6d == index[6:0] ? receive_data : ram_0_109; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2684 = 7'h6e == index[6:0] ? receive_data : ram_0_110; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2685 = 7'h6f == index[6:0] ? receive_data : ram_0_111; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2686 = 7'h70 == index[6:0] ? receive_data : ram_0_112; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2687 = 7'h71 == index[6:0] ? receive_data : ram_0_113; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2688 = 7'h72 == index[6:0] ? receive_data : ram_0_114; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2689 = 7'h73 == index[6:0] ? receive_data : ram_0_115; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2690 = 7'h74 == index[6:0] ? receive_data : ram_0_116; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2691 = 7'h75 == index[6:0] ? receive_data : ram_0_117; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2692 = 7'h76 == index[6:0] ? receive_data : ram_0_118; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2693 = 7'h77 == index[6:0] ? receive_data : ram_0_119; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2694 = 7'h78 == index[6:0] ? receive_data : ram_0_120; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2695 = 7'h79 == index[6:0] ? receive_data : ram_0_121; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2696 = 7'h7a == index[6:0] ? receive_data : ram_0_122; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2697 = 7'h7b == index[6:0] ? receive_data : ram_0_123; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2698 = 7'h7c == index[6:0] ? receive_data : ram_0_124; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2699 = 7'h7d == index[6:0] ? receive_data : ram_0_125; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2700 = 7'h7e == index[6:0] ? receive_data : ram_0_126; // @[d_cache.scala 136:{30,30} 18:24]
  wire [63:0] _GEN_2701 = 7'h7f == index[6:0] ? receive_data : ram_0_127; // @[d_cache.scala 136:{30,30} 18:24]
  wire [31:0] _GEN_2702 = 7'h0 == index[6:0] ? _GEN_16801 : tag_0_0; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2703 = 7'h1 == index[6:0] ? _GEN_16801 : tag_0_1; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2704 = 7'h2 == index[6:0] ? _GEN_16801 : tag_0_2; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2705 = 7'h3 == index[6:0] ? _GEN_16801 : tag_0_3; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2706 = 7'h4 == index[6:0] ? _GEN_16801 : tag_0_4; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2707 = 7'h5 == index[6:0] ? _GEN_16801 : tag_0_5; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2708 = 7'h6 == index[6:0] ? _GEN_16801 : tag_0_6; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2709 = 7'h7 == index[6:0] ? _GEN_16801 : tag_0_7; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2710 = 7'h8 == index[6:0] ? _GEN_16801 : tag_0_8; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2711 = 7'h9 == index[6:0] ? _GEN_16801 : tag_0_9; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2712 = 7'ha == index[6:0] ? _GEN_16801 : tag_0_10; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2713 = 7'hb == index[6:0] ? _GEN_16801 : tag_0_11; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2714 = 7'hc == index[6:0] ? _GEN_16801 : tag_0_12; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2715 = 7'hd == index[6:0] ? _GEN_16801 : tag_0_13; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2716 = 7'he == index[6:0] ? _GEN_16801 : tag_0_14; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2717 = 7'hf == index[6:0] ? _GEN_16801 : tag_0_15; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2718 = 7'h10 == index[6:0] ? _GEN_16801 : tag_0_16; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2719 = 7'h11 == index[6:0] ? _GEN_16801 : tag_0_17; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2720 = 7'h12 == index[6:0] ? _GEN_16801 : tag_0_18; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2721 = 7'h13 == index[6:0] ? _GEN_16801 : tag_0_19; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2722 = 7'h14 == index[6:0] ? _GEN_16801 : tag_0_20; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2723 = 7'h15 == index[6:0] ? _GEN_16801 : tag_0_21; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2724 = 7'h16 == index[6:0] ? _GEN_16801 : tag_0_22; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2725 = 7'h17 == index[6:0] ? _GEN_16801 : tag_0_23; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2726 = 7'h18 == index[6:0] ? _GEN_16801 : tag_0_24; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2727 = 7'h19 == index[6:0] ? _GEN_16801 : tag_0_25; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2728 = 7'h1a == index[6:0] ? _GEN_16801 : tag_0_26; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2729 = 7'h1b == index[6:0] ? _GEN_16801 : tag_0_27; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2730 = 7'h1c == index[6:0] ? _GEN_16801 : tag_0_28; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2731 = 7'h1d == index[6:0] ? _GEN_16801 : tag_0_29; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2732 = 7'h1e == index[6:0] ? _GEN_16801 : tag_0_30; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2733 = 7'h1f == index[6:0] ? _GEN_16801 : tag_0_31; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2734 = 7'h20 == index[6:0] ? _GEN_16801 : tag_0_32; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2735 = 7'h21 == index[6:0] ? _GEN_16801 : tag_0_33; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2736 = 7'h22 == index[6:0] ? _GEN_16801 : tag_0_34; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2737 = 7'h23 == index[6:0] ? _GEN_16801 : tag_0_35; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2738 = 7'h24 == index[6:0] ? _GEN_16801 : tag_0_36; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2739 = 7'h25 == index[6:0] ? _GEN_16801 : tag_0_37; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2740 = 7'h26 == index[6:0] ? _GEN_16801 : tag_0_38; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2741 = 7'h27 == index[6:0] ? _GEN_16801 : tag_0_39; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2742 = 7'h28 == index[6:0] ? _GEN_16801 : tag_0_40; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2743 = 7'h29 == index[6:0] ? _GEN_16801 : tag_0_41; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2744 = 7'h2a == index[6:0] ? _GEN_16801 : tag_0_42; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2745 = 7'h2b == index[6:0] ? _GEN_16801 : tag_0_43; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2746 = 7'h2c == index[6:0] ? _GEN_16801 : tag_0_44; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2747 = 7'h2d == index[6:0] ? _GEN_16801 : tag_0_45; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2748 = 7'h2e == index[6:0] ? _GEN_16801 : tag_0_46; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2749 = 7'h2f == index[6:0] ? _GEN_16801 : tag_0_47; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2750 = 7'h30 == index[6:0] ? _GEN_16801 : tag_0_48; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2751 = 7'h31 == index[6:0] ? _GEN_16801 : tag_0_49; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2752 = 7'h32 == index[6:0] ? _GEN_16801 : tag_0_50; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2753 = 7'h33 == index[6:0] ? _GEN_16801 : tag_0_51; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2754 = 7'h34 == index[6:0] ? _GEN_16801 : tag_0_52; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2755 = 7'h35 == index[6:0] ? _GEN_16801 : tag_0_53; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2756 = 7'h36 == index[6:0] ? _GEN_16801 : tag_0_54; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2757 = 7'h37 == index[6:0] ? _GEN_16801 : tag_0_55; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2758 = 7'h38 == index[6:0] ? _GEN_16801 : tag_0_56; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2759 = 7'h39 == index[6:0] ? _GEN_16801 : tag_0_57; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2760 = 7'h3a == index[6:0] ? _GEN_16801 : tag_0_58; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2761 = 7'h3b == index[6:0] ? _GEN_16801 : tag_0_59; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2762 = 7'h3c == index[6:0] ? _GEN_16801 : tag_0_60; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2763 = 7'h3d == index[6:0] ? _GEN_16801 : tag_0_61; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2764 = 7'h3e == index[6:0] ? _GEN_16801 : tag_0_62; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2765 = 7'h3f == index[6:0] ? _GEN_16801 : tag_0_63; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2766 = 7'h40 == index[6:0] ? _GEN_16801 : tag_0_64; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2767 = 7'h41 == index[6:0] ? _GEN_16801 : tag_0_65; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2768 = 7'h42 == index[6:0] ? _GEN_16801 : tag_0_66; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2769 = 7'h43 == index[6:0] ? _GEN_16801 : tag_0_67; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2770 = 7'h44 == index[6:0] ? _GEN_16801 : tag_0_68; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2771 = 7'h45 == index[6:0] ? _GEN_16801 : tag_0_69; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2772 = 7'h46 == index[6:0] ? _GEN_16801 : tag_0_70; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2773 = 7'h47 == index[6:0] ? _GEN_16801 : tag_0_71; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2774 = 7'h48 == index[6:0] ? _GEN_16801 : tag_0_72; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2775 = 7'h49 == index[6:0] ? _GEN_16801 : tag_0_73; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2776 = 7'h4a == index[6:0] ? _GEN_16801 : tag_0_74; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2777 = 7'h4b == index[6:0] ? _GEN_16801 : tag_0_75; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2778 = 7'h4c == index[6:0] ? _GEN_16801 : tag_0_76; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2779 = 7'h4d == index[6:0] ? _GEN_16801 : tag_0_77; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2780 = 7'h4e == index[6:0] ? _GEN_16801 : tag_0_78; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2781 = 7'h4f == index[6:0] ? _GEN_16801 : tag_0_79; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2782 = 7'h50 == index[6:0] ? _GEN_16801 : tag_0_80; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2783 = 7'h51 == index[6:0] ? _GEN_16801 : tag_0_81; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2784 = 7'h52 == index[6:0] ? _GEN_16801 : tag_0_82; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2785 = 7'h53 == index[6:0] ? _GEN_16801 : tag_0_83; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2786 = 7'h54 == index[6:0] ? _GEN_16801 : tag_0_84; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2787 = 7'h55 == index[6:0] ? _GEN_16801 : tag_0_85; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2788 = 7'h56 == index[6:0] ? _GEN_16801 : tag_0_86; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2789 = 7'h57 == index[6:0] ? _GEN_16801 : tag_0_87; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2790 = 7'h58 == index[6:0] ? _GEN_16801 : tag_0_88; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2791 = 7'h59 == index[6:0] ? _GEN_16801 : tag_0_89; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2792 = 7'h5a == index[6:0] ? _GEN_16801 : tag_0_90; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2793 = 7'h5b == index[6:0] ? _GEN_16801 : tag_0_91; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2794 = 7'h5c == index[6:0] ? _GEN_16801 : tag_0_92; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2795 = 7'h5d == index[6:0] ? _GEN_16801 : tag_0_93; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2796 = 7'h5e == index[6:0] ? _GEN_16801 : tag_0_94; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2797 = 7'h5f == index[6:0] ? _GEN_16801 : tag_0_95; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2798 = 7'h60 == index[6:0] ? _GEN_16801 : tag_0_96; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2799 = 7'h61 == index[6:0] ? _GEN_16801 : tag_0_97; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2800 = 7'h62 == index[6:0] ? _GEN_16801 : tag_0_98; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2801 = 7'h63 == index[6:0] ? _GEN_16801 : tag_0_99; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2802 = 7'h64 == index[6:0] ? _GEN_16801 : tag_0_100; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2803 = 7'h65 == index[6:0] ? _GEN_16801 : tag_0_101; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2804 = 7'h66 == index[6:0] ? _GEN_16801 : tag_0_102; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2805 = 7'h67 == index[6:0] ? _GEN_16801 : tag_0_103; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2806 = 7'h68 == index[6:0] ? _GEN_16801 : tag_0_104; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2807 = 7'h69 == index[6:0] ? _GEN_16801 : tag_0_105; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2808 = 7'h6a == index[6:0] ? _GEN_16801 : tag_0_106; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2809 = 7'h6b == index[6:0] ? _GEN_16801 : tag_0_107; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2810 = 7'h6c == index[6:0] ? _GEN_16801 : tag_0_108; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2811 = 7'h6d == index[6:0] ? _GEN_16801 : tag_0_109; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2812 = 7'h6e == index[6:0] ? _GEN_16801 : tag_0_110; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2813 = 7'h6f == index[6:0] ? _GEN_16801 : tag_0_111; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2814 = 7'h70 == index[6:0] ? _GEN_16801 : tag_0_112; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2815 = 7'h71 == index[6:0] ? _GEN_16801 : tag_0_113; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2816 = 7'h72 == index[6:0] ? _GEN_16801 : tag_0_114; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2817 = 7'h73 == index[6:0] ? _GEN_16801 : tag_0_115; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2818 = 7'h74 == index[6:0] ? _GEN_16801 : tag_0_116; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2819 = 7'h75 == index[6:0] ? _GEN_16801 : tag_0_117; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2820 = 7'h76 == index[6:0] ? _GEN_16801 : tag_0_118; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2821 = 7'h77 == index[6:0] ? _GEN_16801 : tag_0_119; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2822 = 7'h78 == index[6:0] ? _GEN_16801 : tag_0_120; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2823 = 7'h79 == index[6:0] ? _GEN_16801 : tag_0_121; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2824 = 7'h7a == index[6:0] ? _GEN_16801 : tag_0_122; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2825 = 7'h7b == index[6:0] ? _GEN_16801 : tag_0_123; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2826 = 7'h7c == index[6:0] ? _GEN_16801 : tag_0_124; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2827 = 7'h7d == index[6:0] ? _GEN_16801 : tag_0_125; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2828 = 7'h7e == index[6:0] ? _GEN_16801 : tag_0_126; // @[d_cache.scala 137:{30,30} 20:24]
  wire [31:0] _GEN_2829 = 7'h7f == index[6:0] ? _GEN_16801 : tag_0_127; // @[d_cache.scala 137:{30,30} 20:24]
  wire  _GEN_2830 = _GEN_16805 | valid_0_0; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2831 = _GEN_16806 | valid_0_1; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2832 = _GEN_16807 | valid_0_2; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2833 = _GEN_16808 | valid_0_3; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2834 = _GEN_16809 | valid_0_4; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2835 = _GEN_16810 | valid_0_5; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2836 = _GEN_16811 | valid_0_6; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2837 = _GEN_16812 | valid_0_7; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2838 = _GEN_16813 | valid_0_8; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2839 = _GEN_16814 | valid_0_9; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2840 = _GEN_16815 | valid_0_10; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2841 = _GEN_16816 | valid_0_11; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2842 = _GEN_16817 | valid_0_12; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2843 = _GEN_16818 | valid_0_13; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2844 = _GEN_16819 | valid_0_14; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2845 = _GEN_16820 | valid_0_15; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2846 = _GEN_16821 | valid_0_16; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2847 = _GEN_16822 | valid_0_17; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2848 = _GEN_16823 | valid_0_18; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2849 = _GEN_16824 | valid_0_19; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2850 = _GEN_16825 | valid_0_20; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2851 = _GEN_16826 | valid_0_21; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2852 = _GEN_16827 | valid_0_22; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2853 = _GEN_16828 | valid_0_23; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2854 = _GEN_16829 | valid_0_24; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2855 = _GEN_16830 | valid_0_25; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2856 = _GEN_16831 | valid_0_26; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2857 = _GEN_16832 | valid_0_27; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2858 = _GEN_16833 | valid_0_28; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2859 = _GEN_16834 | valid_0_29; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2860 = _GEN_16835 | valid_0_30; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2861 = _GEN_16836 | valid_0_31; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2862 = _GEN_16837 | valid_0_32; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2863 = _GEN_16838 | valid_0_33; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2864 = _GEN_16839 | valid_0_34; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2865 = _GEN_16840 | valid_0_35; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2866 = _GEN_16841 | valid_0_36; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2867 = _GEN_16842 | valid_0_37; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2868 = _GEN_16843 | valid_0_38; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2869 = _GEN_16844 | valid_0_39; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2870 = _GEN_16845 | valid_0_40; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2871 = _GEN_16846 | valid_0_41; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2872 = _GEN_16847 | valid_0_42; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2873 = _GEN_16848 | valid_0_43; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2874 = _GEN_16849 | valid_0_44; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2875 = _GEN_16850 | valid_0_45; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2876 = _GEN_16851 | valid_0_46; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2877 = _GEN_16852 | valid_0_47; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2878 = _GEN_16853 | valid_0_48; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2879 = _GEN_16854 | valid_0_49; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2880 = _GEN_16855 | valid_0_50; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2881 = _GEN_16856 | valid_0_51; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2882 = _GEN_16857 | valid_0_52; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2883 = _GEN_16858 | valid_0_53; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2884 = _GEN_16859 | valid_0_54; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2885 = _GEN_16860 | valid_0_55; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2886 = _GEN_16861 | valid_0_56; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2887 = _GEN_16862 | valid_0_57; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2888 = _GEN_16863 | valid_0_58; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2889 = _GEN_16864 | valid_0_59; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2890 = _GEN_16865 | valid_0_60; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2891 = _GEN_16866 | valid_0_61; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2892 = _GEN_16867 | valid_0_62; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2893 = _GEN_16868 | valid_0_63; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2894 = _GEN_16869 | valid_0_64; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2895 = _GEN_16870 | valid_0_65; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2896 = _GEN_16871 | valid_0_66; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2897 = _GEN_16872 | valid_0_67; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2898 = _GEN_16873 | valid_0_68; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2899 = _GEN_16874 | valid_0_69; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2900 = _GEN_16875 | valid_0_70; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2901 = _GEN_16876 | valid_0_71; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2902 = _GEN_16877 | valid_0_72; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2903 = _GEN_16878 | valid_0_73; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2904 = _GEN_16879 | valid_0_74; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2905 = _GEN_16880 | valid_0_75; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2906 = _GEN_16881 | valid_0_76; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2907 = _GEN_16882 | valid_0_77; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2908 = _GEN_16883 | valid_0_78; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2909 = _GEN_16884 | valid_0_79; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2910 = _GEN_16885 | valid_0_80; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2911 = _GEN_16886 | valid_0_81; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2912 = _GEN_16887 | valid_0_82; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2913 = _GEN_16888 | valid_0_83; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2914 = _GEN_16889 | valid_0_84; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2915 = _GEN_16890 | valid_0_85; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2916 = _GEN_16891 | valid_0_86; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2917 = _GEN_16892 | valid_0_87; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2918 = _GEN_16893 | valid_0_88; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2919 = _GEN_16894 | valid_0_89; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2920 = _GEN_16895 | valid_0_90; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2921 = _GEN_16896 | valid_0_91; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2922 = _GEN_16897 | valid_0_92; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2923 = _GEN_16898 | valid_0_93; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2924 = _GEN_16899 | valid_0_94; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2925 = _GEN_16900 | valid_0_95; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2926 = _GEN_16901 | valid_0_96; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2927 = _GEN_16902 | valid_0_97; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2928 = _GEN_16903 | valid_0_98; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2929 = _GEN_16904 | valid_0_99; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2930 = _GEN_16905 | valid_0_100; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2931 = _GEN_16906 | valid_0_101; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2932 = _GEN_16907 | valid_0_102; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2933 = _GEN_16908 | valid_0_103; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2934 = _GEN_16909 | valid_0_104; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2935 = _GEN_16910 | valid_0_105; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2936 = _GEN_16911 | valid_0_106; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2937 = _GEN_16912 | valid_0_107; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2938 = _GEN_16913 | valid_0_108; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2939 = _GEN_16914 | valid_0_109; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2940 = _GEN_16915 | valid_0_110; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2941 = _GEN_16916 | valid_0_111; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2942 = _GEN_16917 | valid_0_112; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2943 = _GEN_16918 | valid_0_113; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2944 = _GEN_16919 | valid_0_114; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2945 = _GEN_16920 | valid_0_115; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2946 = _GEN_16921 | valid_0_116; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2947 = _GEN_16922 | valid_0_117; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2948 = _GEN_16923 | valid_0_118; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2949 = _GEN_16924 | valid_0_119; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2950 = _GEN_16925 | valid_0_120; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2951 = _GEN_16926 | valid_0_121; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2952 = _GEN_16927 | valid_0_122; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2953 = _GEN_16928 | valid_0_123; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2954 = _GEN_16929 | valid_0_124; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2955 = _GEN_16930 | valid_0_125; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2956 = _GEN_16931 | valid_0_126; // @[d_cache.scala 138:{32,32} 22:26]
  wire  _GEN_2957 = _GEN_16932 | valid_0_127; // @[d_cache.scala 138:{32,32} 22:26]
  wire [63:0] _GEN_2958 = 7'h0 == index[6:0] ? receive_data : ram_1_0; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2959 = 7'h1 == index[6:0] ? receive_data : ram_1_1; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2960 = 7'h2 == index[6:0] ? receive_data : ram_1_2; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2961 = 7'h3 == index[6:0] ? receive_data : ram_1_3; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2962 = 7'h4 == index[6:0] ? receive_data : ram_1_4; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2963 = 7'h5 == index[6:0] ? receive_data : ram_1_5; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2964 = 7'h6 == index[6:0] ? receive_data : ram_1_6; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2965 = 7'h7 == index[6:0] ? receive_data : ram_1_7; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2966 = 7'h8 == index[6:0] ? receive_data : ram_1_8; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2967 = 7'h9 == index[6:0] ? receive_data : ram_1_9; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2968 = 7'ha == index[6:0] ? receive_data : ram_1_10; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2969 = 7'hb == index[6:0] ? receive_data : ram_1_11; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2970 = 7'hc == index[6:0] ? receive_data : ram_1_12; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2971 = 7'hd == index[6:0] ? receive_data : ram_1_13; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2972 = 7'he == index[6:0] ? receive_data : ram_1_14; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2973 = 7'hf == index[6:0] ? receive_data : ram_1_15; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2974 = 7'h10 == index[6:0] ? receive_data : ram_1_16; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2975 = 7'h11 == index[6:0] ? receive_data : ram_1_17; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2976 = 7'h12 == index[6:0] ? receive_data : ram_1_18; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2977 = 7'h13 == index[6:0] ? receive_data : ram_1_19; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2978 = 7'h14 == index[6:0] ? receive_data : ram_1_20; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2979 = 7'h15 == index[6:0] ? receive_data : ram_1_21; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2980 = 7'h16 == index[6:0] ? receive_data : ram_1_22; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2981 = 7'h17 == index[6:0] ? receive_data : ram_1_23; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2982 = 7'h18 == index[6:0] ? receive_data : ram_1_24; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2983 = 7'h19 == index[6:0] ? receive_data : ram_1_25; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2984 = 7'h1a == index[6:0] ? receive_data : ram_1_26; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2985 = 7'h1b == index[6:0] ? receive_data : ram_1_27; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2986 = 7'h1c == index[6:0] ? receive_data : ram_1_28; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2987 = 7'h1d == index[6:0] ? receive_data : ram_1_29; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2988 = 7'h1e == index[6:0] ? receive_data : ram_1_30; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2989 = 7'h1f == index[6:0] ? receive_data : ram_1_31; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2990 = 7'h20 == index[6:0] ? receive_data : ram_1_32; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2991 = 7'h21 == index[6:0] ? receive_data : ram_1_33; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2992 = 7'h22 == index[6:0] ? receive_data : ram_1_34; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2993 = 7'h23 == index[6:0] ? receive_data : ram_1_35; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2994 = 7'h24 == index[6:0] ? receive_data : ram_1_36; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2995 = 7'h25 == index[6:0] ? receive_data : ram_1_37; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2996 = 7'h26 == index[6:0] ? receive_data : ram_1_38; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2997 = 7'h27 == index[6:0] ? receive_data : ram_1_39; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2998 = 7'h28 == index[6:0] ? receive_data : ram_1_40; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_2999 = 7'h29 == index[6:0] ? receive_data : ram_1_41; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3000 = 7'h2a == index[6:0] ? receive_data : ram_1_42; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3001 = 7'h2b == index[6:0] ? receive_data : ram_1_43; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3002 = 7'h2c == index[6:0] ? receive_data : ram_1_44; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3003 = 7'h2d == index[6:0] ? receive_data : ram_1_45; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3004 = 7'h2e == index[6:0] ? receive_data : ram_1_46; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3005 = 7'h2f == index[6:0] ? receive_data : ram_1_47; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3006 = 7'h30 == index[6:0] ? receive_data : ram_1_48; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3007 = 7'h31 == index[6:0] ? receive_data : ram_1_49; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3008 = 7'h32 == index[6:0] ? receive_data : ram_1_50; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3009 = 7'h33 == index[6:0] ? receive_data : ram_1_51; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3010 = 7'h34 == index[6:0] ? receive_data : ram_1_52; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3011 = 7'h35 == index[6:0] ? receive_data : ram_1_53; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3012 = 7'h36 == index[6:0] ? receive_data : ram_1_54; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3013 = 7'h37 == index[6:0] ? receive_data : ram_1_55; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3014 = 7'h38 == index[6:0] ? receive_data : ram_1_56; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3015 = 7'h39 == index[6:0] ? receive_data : ram_1_57; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3016 = 7'h3a == index[6:0] ? receive_data : ram_1_58; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3017 = 7'h3b == index[6:0] ? receive_data : ram_1_59; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3018 = 7'h3c == index[6:0] ? receive_data : ram_1_60; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3019 = 7'h3d == index[6:0] ? receive_data : ram_1_61; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3020 = 7'h3e == index[6:0] ? receive_data : ram_1_62; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3021 = 7'h3f == index[6:0] ? receive_data : ram_1_63; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3022 = 7'h40 == index[6:0] ? receive_data : ram_1_64; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3023 = 7'h41 == index[6:0] ? receive_data : ram_1_65; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3024 = 7'h42 == index[6:0] ? receive_data : ram_1_66; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3025 = 7'h43 == index[6:0] ? receive_data : ram_1_67; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3026 = 7'h44 == index[6:0] ? receive_data : ram_1_68; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3027 = 7'h45 == index[6:0] ? receive_data : ram_1_69; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3028 = 7'h46 == index[6:0] ? receive_data : ram_1_70; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3029 = 7'h47 == index[6:0] ? receive_data : ram_1_71; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3030 = 7'h48 == index[6:0] ? receive_data : ram_1_72; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3031 = 7'h49 == index[6:0] ? receive_data : ram_1_73; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3032 = 7'h4a == index[6:0] ? receive_data : ram_1_74; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3033 = 7'h4b == index[6:0] ? receive_data : ram_1_75; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3034 = 7'h4c == index[6:0] ? receive_data : ram_1_76; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3035 = 7'h4d == index[6:0] ? receive_data : ram_1_77; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3036 = 7'h4e == index[6:0] ? receive_data : ram_1_78; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3037 = 7'h4f == index[6:0] ? receive_data : ram_1_79; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3038 = 7'h50 == index[6:0] ? receive_data : ram_1_80; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3039 = 7'h51 == index[6:0] ? receive_data : ram_1_81; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3040 = 7'h52 == index[6:0] ? receive_data : ram_1_82; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3041 = 7'h53 == index[6:0] ? receive_data : ram_1_83; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3042 = 7'h54 == index[6:0] ? receive_data : ram_1_84; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3043 = 7'h55 == index[6:0] ? receive_data : ram_1_85; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3044 = 7'h56 == index[6:0] ? receive_data : ram_1_86; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3045 = 7'h57 == index[6:0] ? receive_data : ram_1_87; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3046 = 7'h58 == index[6:0] ? receive_data : ram_1_88; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3047 = 7'h59 == index[6:0] ? receive_data : ram_1_89; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3048 = 7'h5a == index[6:0] ? receive_data : ram_1_90; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3049 = 7'h5b == index[6:0] ? receive_data : ram_1_91; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3050 = 7'h5c == index[6:0] ? receive_data : ram_1_92; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3051 = 7'h5d == index[6:0] ? receive_data : ram_1_93; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3052 = 7'h5e == index[6:0] ? receive_data : ram_1_94; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3053 = 7'h5f == index[6:0] ? receive_data : ram_1_95; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3054 = 7'h60 == index[6:0] ? receive_data : ram_1_96; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3055 = 7'h61 == index[6:0] ? receive_data : ram_1_97; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3056 = 7'h62 == index[6:0] ? receive_data : ram_1_98; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3057 = 7'h63 == index[6:0] ? receive_data : ram_1_99; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3058 = 7'h64 == index[6:0] ? receive_data : ram_1_100; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3059 = 7'h65 == index[6:0] ? receive_data : ram_1_101; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3060 = 7'h66 == index[6:0] ? receive_data : ram_1_102; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3061 = 7'h67 == index[6:0] ? receive_data : ram_1_103; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3062 = 7'h68 == index[6:0] ? receive_data : ram_1_104; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3063 = 7'h69 == index[6:0] ? receive_data : ram_1_105; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3064 = 7'h6a == index[6:0] ? receive_data : ram_1_106; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3065 = 7'h6b == index[6:0] ? receive_data : ram_1_107; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3066 = 7'h6c == index[6:0] ? receive_data : ram_1_108; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3067 = 7'h6d == index[6:0] ? receive_data : ram_1_109; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3068 = 7'h6e == index[6:0] ? receive_data : ram_1_110; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3069 = 7'h6f == index[6:0] ? receive_data : ram_1_111; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3070 = 7'h70 == index[6:0] ? receive_data : ram_1_112; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3071 = 7'h71 == index[6:0] ? receive_data : ram_1_113; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3072 = 7'h72 == index[6:0] ? receive_data : ram_1_114; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3073 = 7'h73 == index[6:0] ? receive_data : ram_1_115; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3074 = 7'h74 == index[6:0] ? receive_data : ram_1_116; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3075 = 7'h75 == index[6:0] ? receive_data : ram_1_117; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3076 = 7'h76 == index[6:0] ? receive_data : ram_1_118; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3077 = 7'h77 == index[6:0] ? receive_data : ram_1_119; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3078 = 7'h78 == index[6:0] ? receive_data : ram_1_120; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3079 = 7'h79 == index[6:0] ? receive_data : ram_1_121; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3080 = 7'h7a == index[6:0] ? receive_data : ram_1_122; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3081 = 7'h7b == index[6:0] ? receive_data : ram_1_123; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3082 = 7'h7c == index[6:0] ? receive_data : ram_1_124; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3083 = 7'h7d == index[6:0] ? receive_data : ram_1_125; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3084 = 7'h7e == index[6:0] ? receive_data : ram_1_126; // @[d_cache.scala 142:{30,30} 19:24]
  wire [63:0] _GEN_3085 = 7'h7f == index[6:0] ? receive_data : ram_1_127; // @[d_cache.scala 142:{30,30} 19:24]
  wire [31:0] _GEN_3086 = 7'h0 == index[6:0] ? _GEN_16801 : tag_1_0; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3087 = 7'h1 == index[6:0] ? _GEN_16801 : tag_1_1; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3088 = 7'h2 == index[6:0] ? _GEN_16801 : tag_1_2; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3089 = 7'h3 == index[6:0] ? _GEN_16801 : tag_1_3; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3090 = 7'h4 == index[6:0] ? _GEN_16801 : tag_1_4; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3091 = 7'h5 == index[6:0] ? _GEN_16801 : tag_1_5; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3092 = 7'h6 == index[6:0] ? _GEN_16801 : tag_1_6; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3093 = 7'h7 == index[6:0] ? _GEN_16801 : tag_1_7; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3094 = 7'h8 == index[6:0] ? _GEN_16801 : tag_1_8; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3095 = 7'h9 == index[6:0] ? _GEN_16801 : tag_1_9; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3096 = 7'ha == index[6:0] ? _GEN_16801 : tag_1_10; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3097 = 7'hb == index[6:0] ? _GEN_16801 : tag_1_11; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3098 = 7'hc == index[6:0] ? _GEN_16801 : tag_1_12; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3099 = 7'hd == index[6:0] ? _GEN_16801 : tag_1_13; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3100 = 7'he == index[6:0] ? _GEN_16801 : tag_1_14; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3101 = 7'hf == index[6:0] ? _GEN_16801 : tag_1_15; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3102 = 7'h10 == index[6:0] ? _GEN_16801 : tag_1_16; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3103 = 7'h11 == index[6:0] ? _GEN_16801 : tag_1_17; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3104 = 7'h12 == index[6:0] ? _GEN_16801 : tag_1_18; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3105 = 7'h13 == index[6:0] ? _GEN_16801 : tag_1_19; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3106 = 7'h14 == index[6:0] ? _GEN_16801 : tag_1_20; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3107 = 7'h15 == index[6:0] ? _GEN_16801 : tag_1_21; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3108 = 7'h16 == index[6:0] ? _GEN_16801 : tag_1_22; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3109 = 7'h17 == index[6:0] ? _GEN_16801 : tag_1_23; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3110 = 7'h18 == index[6:0] ? _GEN_16801 : tag_1_24; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3111 = 7'h19 == index[6:0] ? _GEN_16801 : tag_1_25; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3112 = 7'h1a == index[6:0] ? _GEN_16801 : tag_1_26; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3113 = 7'h1b == index[6:0] ? _GEN_16801 : tag_1_27; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3114 = 7'h1c == index[6:0] ? _GEN_16801 : tag_1_28; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3115 = 7'h1d == index[6:0] ? _GEN_16801 : tag_1_29; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3116 = 7'h1e == index[6:0] ? _GEN_16801 : tag_1_30; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3117 = 7'h1f == index[6:0] ? _GEN_16801 : tag_1_31; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3118 = 7'h20 == index[6:0] ? _GEN_16801 : tag_1_32; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3119 = 7'h21 == index[6:0] ? _GEN_16801 : tag_1_33; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3120 = 7'h22 == index[6:0] ? _GEN_16801 : tag_1_34; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3121 = 7'h23 == index[6:0] ? _GEN_16801 : tag_1_35; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3122 = 7'h24 == index[6:0] ? _GEN_16801 : tag_1_36; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3123 = 7'h25 == index[6:0] ? _GEN_16801 : tag_1_37; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3124 = 7'h26 == index[6:0] ? _GEN_16801 : tag_1_38; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3125 = 7'h27 == index[6:0] ? _GEN_16801 : tag_1_39; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3126 = 7'h28 == index[6:0] ? _GEN_16801 : tag_1_40; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3127 = 7'h29 == index[6:0] ? _GEN_16801 : tag_1_41; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3128 = 7'h2a == index[6:0] ? _GEN_16801 : tag_1_42; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3129 = 7'h2b == index[6:0] ? _GEN_16801 : tag_1_43; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3130 = 7'h2c == index[6:0] ? _GEN_16801 : tag_1_44; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3131 = 7'h2d == index[6:0] ? _GEN_16801 : tag_1_45; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3132 = 7'h2e == index[6:0] ? _GEN_16801 : tag_1_46; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3133 = 7'h2f == index[6:0] ? _GEN_16801 : tag_1_47; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3134 = 7'h30 == index[6:0] ? _GEN_16801 : tag_1_48; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3135 = 7'h31 == index[6:0] ? _GEN_16801 : tag_1_49; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3136 = 7'h32 == index[6:0] ? _GEN_16801 : tag_1_50; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3137 = 7'h33 == index[6:0] ? _GEN_16801 : tag_1_51; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3138 = 7'h34 == index[6:0] ? _GEN_16801 : tag_1_52; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3139 = 7'h35 == index[6:0] ? _GEN_16801 : tag_1_53; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3140 = 7'h36 == index[6:0] ? _GEN_16801 : tag_1_54; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3141 = 7'h37 == index[6:0] ? _GEN_16801 : tag_1_55; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3142 = 7'h38 == index[6:0] ? _GEN_16801 : tag_1_56; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3143 = 7'h39 == index[6:0] ? _GEN_16801 : tag_1_57; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3144 = 7'h3a == index[6:0] ? _GEN_16801 : tag_1_58; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3145 = 7'h3b == index[6:0] ? _GEN_16801 : tag_1_59; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3146 = 7'h3c == index[6:0] ? _GEN_16801 : tag_1_60; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3147 = 7'h3d == index[6:0] ? _GEN_16801 : tag_1_61; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3148 = 7'h3e == index[6:0] ? _GEN_16801 : tag_1_62; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3149 = 7'h3f == index[6:0] ? _GEN_16801 : tag_1_63; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3150 = 7'h40 == index[6:0] ? _GEN_16801 : tag_1_64; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3151 = 7'h41 == index[6:0] ? _GEN_16801 : tag_1_65; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3152 = 7'h42 == index[6:0] ? _GEN_16801 : tag_1_66; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3153 = 7'h43 == index[6:0] ? _GEN_16801 : tag_1_67; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3154 = 7'h44 == index[6:0] ? _GEN_16801 : tag_1_68; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3155 = 7'h45 == index[6:0] ? _GEN_16801 : tag_1_69; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3156 = 7'h46 == index[6:0] ? _GEN_16801 : tag_1_70; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3157 = 7'h47 == index[6:0] ? _GEN_16801 : tag_1_71; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3158 = 7'h48 == index[6:0] ? _GEN_16801 : tag_1_72; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3159 = 7'h49 == index[6:0] ? _GEN_16801 : tag_1_73; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3160 = 7'h4a == index[6:0] ? _GEN_16801 : tag_1_74; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3161 = 7'h4b == index[6:0] ? _GEN_16801 : tag_1_75; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3162 = 7'h4c == index[6:0] ? _GEN_16801 : tag_1_76; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3163 = 7'h4d == index[6:0] ? _GEN_16801 : tag_1_77; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3164 = 7'h4e == index[6:0] ? _GEN_16801 : tag_1_78; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3165 = 7'h4f == index[6:0] ? _GEN_16801 : tag_1_79; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3166 = 7'h50 == index[6:0] ? _GEN_16801 : tag_1_80; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3167 = 7'h51 == index[6:0] ? _GEN_16801 : tag_1_81; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3168 = 7'h52 == index[6:0] ? _GEN_16801 : tag_1_82; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3169 = 7'h53 == index[6:0] ? _GEN_16801 : tag_1_83; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3170 = 7'h54 == index[6:0] ? _GEN_16801 : tag_1_84; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3171 = 7'h55 == index[6:0] ? _GEN_16801 : tag_1_85; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3172 = 7'h56 == index[6:0] ? _GEN_16801 : tag_1_86; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3173 = 7'h57 == index[6:0] ? _GEN_16801 : tag_1_87; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3174 = 7'h58 == index[6:0] ? _GEN_16801 : tag_1_88; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3175 = 7'h59 == index[6:0] ? _GEN_16801 : tag_1_89; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3176 = 7'h5a == index[6:0] ? _GEN_16801 : tag_1_90; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3177 = 7'h5b == index[6:0] ? _GEN_16801 : tag_1_91; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3178 = 7'h5c == index[6:0] ? _GEN_16801 : tag_1_92; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3179 = 7'h5d == index[6:0] ? _GEN_16801 : tag_1_93; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3180 = 7'h5e == index[6:0] ? _GEN_16801 : tag_1_94; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3181 = 7'h5f == index[6:0] ? _GEN_16801 : tag_1_95; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3182 = 7'h60 == index[6:0] ? _GEN_16801 : tag_1_96; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3183 = 7'h61 == index[6:0] ? _GEN_16801 : tag_1_97; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3184 = 7'h62 == index[6:0] ? _GEN_16801 : tag_1_98; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3185 = 7'h63 == index[6:0] ? _GEN_16801 : tag_1_99; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3186 = 7'h64 == index[6:0] ? _GEN_16801 : tag_1_100; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3187 = 7'h65 == index[6:0] ? _GEN_16801 : tag_1_101; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3188 = 7'h66 == index[6:0] ? _GEN_16801 : tag_1_102; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3189 = 7'h67 == index[6:0] ? _GEN_16801 : tag_1_103; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3190 = 7'h68 == index[6:0] ? _GEN_16801 : tag_1_104; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3191 = 7'h69 == index[6:0] ? _GEN_16801 : tag_1_105; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3192 = 7'h6a == index[6:0] ? _GEN_16801 : tag_1_106; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3193 = 7'h6b == index[6:0] ? _GEN_16801 : tag_1_107; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3194 = 7'h6c == index[6:0] ? _GEN_16801 : tag_1_108; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3195 = 7'h6d == index[6:0] ? _GEN_16801 : tag_1_109; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3196 = 7'h6e == index[6:0] ? _GEN_16801 : tag_1_110; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3197 = 7'h6f == index[6:0] ? _GEN_16801 : tag_1_111; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3198 = 7'h70 == index[6:0] ? _GEN_16801 : tag_1_112; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3199 = 7'h71 == index[6:0] ? _GEN_16801 : tag_1_113; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3200 = 7'h72 == index[6:0] ? _GEN_16801 : tag_1_114; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3201 = 7'h73 == index[6:0] ? _GEN_16801 : tag_1_115; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3202 = 7'h74 == index[6:0] ? _GEN_16801 : tag_1_116; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3203 = 7'h75 == index[6:0] ? _GEN_16801 : tag_1_117; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3204 = 7'h76 == index[6:0] ? _GEN_16801 : tag_1_118; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3205 = 7'h77 == index[6:0] ? _GEN_16801 : tag_1_119; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3206 = 7'h78 == index[6:0] ? _GEN_16801 : tag_1_120; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3207 = 7'h79 == index[6:0] ? _GEN_16801 : tag_1_121; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3208 = 7'h7a == index[6:0] ? _GEN_16801 : tag_1_122; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3209 = 7'h7b == index[6:0] ? _GEN_16801 : tag_1_123; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3210 = 7'h7c == index[6:0] ? _GEN_16801 : tag_1_124; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3211 = 7'h7d == index[6:0] ? _GEN_16801 : tag_1_125; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3212 = 7'h7e == index[6:0] ? _GEN_16801 : tag_1_126; // @[d_cache.scala 143:{30,30} 21:24]
  wire [31:0] _GEN_3213 = 7'h7f == index[6:0] ? _GEN_16801 : tag_1_127; // @[d_cache.scala 143:{30,30} 21:24]
  wire  _GEN_3214 = _GEN_16805 | valid_1_0; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3215 = _GEN_16806 | valid_1_1; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3216 = _GEN_16807 | valid_1_2; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3217 = _GEN_16808 | valid_1_3; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3218 = _GEN_16809 | valid_1_4; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3219 = _GEN_16810 | valid_1_5; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3220 = _GEN_16811 | valid_1_6; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3221 = _GEN_16812 | valid_1_7; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3222 = _GEN_16813 | valid_1_8; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3223 = _GEN_16814 | valid_1_9; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3224 = _GEN_16815 | valid_1_10; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3225 = _GEN_16816 | valid_1_11; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3226 = _GEN_16817 | valid_1_12; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3227 = _GEN_16818 | valid_1_13; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3228 = _GEN_16819 | valid_1_14; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3229 = _GEN_16820 | valid_1_15; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3230 = _GEN_16821 | valid_1_16; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3231 = _GEN_16822 | valid_1_17; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3232 = _GEN_16823 | valid_1_18; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3233 = _GEN_16824 | valid_1_19; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3234 = _GEN_16825 | valid_1_20; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3235 = _GEN_16826 | valid_1_21; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3236 = _GEN_16827 | valid_1_22; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3237 = _GEN_16828 | valid_1_23; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3238 = _GEN_16829 | valid_1_24; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3239 = _GEN_16830 | valid_1_25; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3240 = _GEN_16831 | valid_1_26; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3241 = _GEN_16832 | valid_1_27; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3242 = _GEN_16833 | valid_1_28; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3243 = _GEN_16834 | valid_1_29; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3244 = _GEN_16835 | valid_1_30; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3245 = _GEN_16836 | valid_1_31; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3246 = _GEN_16837 | valid_1_32; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3247 = _GEN_16838 | valid_1_33; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3248 = _GEN_16839 | valid_1_34; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3249 = _GEN_16840 | valid_1_35; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3250 = _GEN_16841 | valid_1_36; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3251 = _GEN_16842 | valid_1_37; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3252 = _GEN_16843 | valid_1_38; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3253 = _GEN_16844 | valid_1_39; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3254 = _GEN_16845 | valid_1_40; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3255 = _GEN_16846 | valid_1_41; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3256 = _GEN_16847 | valid_1_42; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3257 = _GEN_16848 | valid_1_43; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3258 = _GEN_16849 | valid_1_44; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3259 = _GEN_16850 | valid_1_45; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3260 = _GEN_16851 | valid_1_46; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3261 = _GEN_16852 | valid_1_47; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3262 = _GEN_16853 | valid_1_48; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3263 = _GEN_16854 | valid_1_49; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3264 = _GEN_16855 | valid_1_50; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3265 = _GEN_16856 | valid_1_51; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3266 = _GEN_16857 | valid_1_52; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3267 = _GEN_16858 | valid_1_53; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3268 = _GEN_16859 | valid_1_54; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3269 = _GEN_16860 | valid_1_55; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3270 = _GEN_16861 | valid_1_56; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3271 = _GEN_16862 | valid_1_57; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3272 = _GEN_16863 | valid_1_58; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3273 = _GEN_16864 | valid_1_59; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3274 = _GEN_16865 | valid_1_60; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3275 = _GEN_16866 | valid_1_61; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3276 = _GEN_16867 | valid_1_62; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3277 = _GEN_16868 | valid_1_63; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3278 = _GEN_16869 | valid_1_64; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3279 = _GEN_16870 | valid_1_65; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3280 = _GEN_16871 | valid_1_66; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3281 = _GEN_16872 | valid_1_67; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3282 = _GEN_16873 | valid_1_68; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3283 = _GEN_16874 | valid_1_69; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3284 = _GEN_16875 | valid_1_70; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3285 = _GEN_16876 | valid_1_71; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3286 = _GEN_16877 | valid_1_72; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3287 = _GEN_16878 | valid_1_73; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3288 = _GEN_16879 | valid_1_74; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3289 = _GEN_16880 | valid_1_75; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3290 = _GEN_16881 | valid_1_76; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3291 = _GEN_16882 | valid_1_77; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3292 = _GEN_16883 | valid_1_78; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3293 = _GEN_16884 | valid_1_79; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3294 = _GEN_16885 | valid_1_80; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3295 = _GEN_16886 | valid_1_81; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3296 = _GEN_16887 | valid_1_82; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3297 = _GEN_16888 | valid_1_83; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3298 = _GEN_16889 | valid_1_84; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3299 = _GEN_16890 | valid_1_85; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3300 = _GEN_16891 | valid_1_86; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3301 = _GEN_16892 | valid_1_87; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3302 = _GEN_16893 | valid_1_88; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3303 = _GEN_16894 | valid_1_89; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3304 = _GEN_16895 | valid_1_90; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3305 = _GEN_16896 | valid_1_91; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3306 = _GEN_16897 | valid_1_92; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3307 = _GEN_16898 | valid_1_93; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3308 = _GEN_16899 | valid_1_94; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3309 = _GEN_16900 | valid_1_95; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3310 = _GEN_16901 | valid_1_96; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3311 = _GEN_16902 | valid_1_97; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3312 = _GEN_16903 | valid_1_98; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3313 = _GEN_16904 | valid_1_99; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3314 = _GEN_16905 | valid_1_100; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3315 = _GEN_16906 | valid_1_101; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3316 = _GEN_16907 | valid_1_102; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3317 = _GEN_16908 | valid_1_103; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3318 = _GEN_16909 | valid_1_104; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3319 = _GEN_16910 | valid_1_105; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3320 = _GEN_16911 | valid_1_106; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3321 = _GEN_16912 | valid_1_107; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3322 = _GEN_16913 | valid_1_108; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3323 = _GEN_16914 | valid_1_109; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3324 = _GEN_16915 | valid_1_110; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3325 = _GEN_16916 | valid_1_111; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3326 = _GEN_16917 | valid_1_112; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3327 = _GEN_16918 | valid_1_113; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3328 = _GEN_16919 | valid_1_114; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3329 = _GEN_16920 | valid_1_115; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3330 = _GEN_16921 | valid_1_116; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3331 = _GEN_16922 | valid_1_117; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3332 = _GEN_16923 | valid_1_118; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3333 = _GEN_16924 | valid_1_119; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3334 = _GEN_16925 | valid_1_120; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3335 = _GEN_16926 | valid_1_121; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3336 = _GEN_16927 | valid_1_122; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3337 = _GEN_16928 | valid_1_123; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3338 = _GEN_16929 | valid_1_124; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3339 = _GEN_16930 | valid_1_125; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3340 = _GEN_16931 | valid_1_126; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _GEN_3341 = _GEN_16932 | valid_1_127; // @[d_cache.scala 144:{32,32} 23:26]
  wire  _T_48 = ~quene; // @[d_cache.scala 147:27]
  wire [41:0] _write_back_addr_T_1 = {_GEN_127, 10'h0}; // @[d_cache.scala 151:58]
  wire [34:0] _write_back_addr_T_2 = {index, 3'h0}; // @[d_cache.scala 151:74]
  wire [41:0] _GEN_17319 = {{7'd0}, _write_back_addr_T_2}; // @[d_cache.scala 151:65]
  wire [41:0] _write_back_addr_T_3 = _write_back_addr_T_1 | _GEN_17319; // @[d_cache.scala 151:65]
  wire  _GEN_3982 = 7'h0 == index[6:0] ? 1'h0 : dirty_0_0; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3983 = 7'h1 == index[6:0] ? 1'h0 : dirty_0_1; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3984 = 7'h2 == index[6:0] ? 1'h0 : dirty_0_2; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3985 = 7'h3 == index[6:0] ? 1'h0 : dirty_0_3; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3986 = 7'h4 == index[6:0] ? 1'h0 : dirty_0_4; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3987 = 7'h5 == index[6:0] ? 1'h0 : dirty_0_5; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3988 = 7'h6 == index[6:0] ? 1'h0 : dirty_0_6; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3989 = 7'h7 == index[6:0] ? 1'h0 : dirty_0_7; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3990 = 7'h8 == index[6:0] ? 1'h0 : dirty_0_8; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3991 = 7'h9 == index[6:0] ? 1'h0 : dirty_0_9; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3992 = 7'ha == index[6:0] ? 1'h0 : dirty_0_10; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3993 = 7'hb == index[6:0] ? 1'h0 : dirty_0_11; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3994 = 7'hc == index[6:0] ? 1'h0 : dirty_0_12; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3995 = 7'hd == index[6:0] ? 1'h0 : dirty_0_13; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3996 = 7'he == index[6:0] ? 1'h0 : dirty_0_14; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3997 = 7'hf == index[6:0] ? 1'h0 : dirty_0_15; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3998 = 7'h10 == index[6:0] ? 1'h0 : dirty_0_16; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_3999 = 7'h11 == index[6:0] ? 1'h0 : dirty_0_17; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4000 = 7'h12 == index[6:0] ? 1'h0 : dirty_0_18; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4001 = 7'h13 == index[6:0] ? 1'h0 : dirty_0_19; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4002 = 7'h14 == index[6:0] ? 1'h0 : dirty_0_20; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4003 = 7'h15 == index[6:0] ? 1'h0 : dirty_0_21; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4004 = 7'h16 == index[6:0] ? 1'h0 : dirty_0_22; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4005 = 7'h17 == index[6:0] ? 1'h0 : dirty_0_23; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4006 = 7'h18 == index[6:0] ? 1'h0 : dirty_0_24; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4007 = 7'h19 == index[6:0] ? 1'h0 : dirty_0_25; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4008 = 7'h1a == index[6:0] ? 1'h0 : dirty_0_26; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4009 = 7'h1b == index[6:0] ? 1'h0 : dirty_0_27; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4010 = 7'h1c == index[6:0] ? 1'h0 : dirty_0_28; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4011 = 7'h1d == index[6:0] ? 1'h0 : dirty_0_29; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4012 = 7'h1e == index[6:0] ? 1'h0 : dirty_0_30; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4013 = 7'h1f == index[6:0] ? 1'h0 : dirty_0_31; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4014 = 7'h20 == index[6:0] ? 1'h0 : dirty_0_32; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4015 = 7'h21 == index[6:0] ? 1'h0 : dirty_0_33; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4016 = 7'h22 == index[6:0] ? 1'h0 : dirty_0_34; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4017 = 7'h23 == index[6:0] ? 1'h0 : dirty_0_35; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4018 = 7'h24 == index[6:0] ? 1'h0 : dirty_0_36; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4019 = 7'h25 == index[6:0] ? 1'h0 : dirty_0_37; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4020 = 7'h26 == index[6:0] ? 1'h0 : dirty_0_38; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4021 = 7'h27 == index[6:0] ? 1'h0 : dirty_0_39; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4022 = 7'h28 == index[6:0] ? 1'h0 : dirty_0_40; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4023 = 7'h29 == index[6:0] ? 1'h0 : dirty_0_41; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4024 = 7'h2a == index[6:0] ? 1'h0 : dirty_0_42; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4025 = 7'h2b == index[6:0] ? 1'h0 : dirty_0_43; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4026 = 7'h2c == index[6:0] ? 1'h0 : dirty_0_44; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4027 = 7'h2d == index[6:0] ? 1'h0 : dirty_0_45; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4028 = 7'h2e == index[6:0] ? 1'h0 : dirty_0_46; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4029 = 7'h2f == index[6:0] ? 1'h0 : dirty_0_47; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4030 = 7'h30 == index[6:0] ? 1'h0 : dirty_0_48; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4031 = 7'h31 == index[6:0] ? 1'h0 : dirty_0_49; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4032 = 7'h32 == index[6:0] ? 1'h0 : dirty_0_50; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4033 = 7'h33 == index[6:0] ? 1'h0 : dirty_0_51; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4034 = 7'h34 == index[6:0] ? 1'h0 : dirty_0_52; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4035 = 7'h35 == index[6:0] ? 1'h0 : dirty_0_53; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4036 = 7'h36 == index[6:0] ? 1'h0 : dirty_0_54; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4037 = 7'h37 == index[6:0] ? 1'h0 : dirty_0_55; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4038 = 7'h38 == index[6:0] ? 1'h0 : dirty_0_56; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4039 = 7'h39 == index[6:0] ? 1'h0 : dirty_0_57; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4040 = 7'h3a == index[6:0] ? 1'h0 : dirty_0_58; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4041 = 7'h3b == index[6:0] ? 1'h0 : dirty_0_59; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4042 = 7'h3c == index[6:0] ? 1'h0 : dirty_0_60; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4043 = 7'h3d == index[6:0] ? 1'h0 : dirty_0_61; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4044 = 7'h3e == index[6:0] ? 1'h0 : dirty_0_62; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4045 = 7'h3f == index[6:0] ? 1'h0 : dirty_0_63; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4046 = 7'h40 == index[6:0] ? 1'h0 : dirty_0_64; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4047 = 7'h41 == index[6:0] ? 1'h0 : dirty_0_65; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4048 = 7'h42 == index[6:0] ? 1'h0 : dirty_0_66; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4049 = 7'h43 == index[6:0] ? 1'h0 : dirty_0_67; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4050 = 7'h44 == index[6:0] ? 1'h0 : dirty_0_68; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4051 = 7'h45 == index[6:0] ? 1'h0 : dirty_0_69; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4052 = 7'h46 == index[6:0] ? 1'h0 : dirty_0_70; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4053 = 7'h47 == index[6:0] ? 1'h0 : dirty_0_71; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4054 = 7'h48 == index[6:0] ? 1'h0 : dirty_0_72; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4055 = 7'h49 == index[6:0] ? 1'h0 : dirty_0_73; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4056 = 7'h4a == index[6:0] ? 1'h0 : dirty_0_74; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4057 = 7'h4b == index[6:0] ? 1'h0 : dirty_0_75; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4058 = 7'h4c == index[6:0] ? 1'h0 : dirty_0_76; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4059 = 7'h4d == index[6:0] ? 1'h0 : dirty_0_77; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4060 = 7'h4e == index[6:0] ? 1'h0 : dirty_0_78; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4061 = 7'h4f == index[6:0] ? 1'h0 : dirty_0_79; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4062 = 7'h50 == index[6:0] ? 1'h0 : dirty_0_80; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4063 = 7'h51 == index[6:0] ? 1'h0 : dirty_0_81; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4064 = 7'h52 == index[6:0] ? 1'h0 : dirty_0_82; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4065 = 7'h53 == index[6:0] ? 1'h0 : dirty_0_83; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4066 = 7'h54 == index[6:0] ? 1'h0 : dirty_0_84; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4067 = 7'h55 == index[6:0] ? 1'h0 : dirty_0_85; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4068 = 7'h56 == index[6:0] ? 1'h0 : dirty_0_86; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4069 = 7'h57 == index[6:0] ? 1'h0 : dirty_0_87; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4070 = 7'h58 == index[6:0] ? 1'h0 : dirty_0_88; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4071 = 7'h59 == index[6:0] ? 1'h0 : dirty_0_89; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4072 = 7'h5a == index[6:0] ? 1'h0 : dirty_0_90; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4073 = 7'h5b == index[6:0] ? 1'h0 : dirty_0_91; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4074 = 7'h5c == index[6:0] ? 1'h0 : dirty_0_92; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4075 = 7'h5d == index[6:0] ? 1'h0 : dirty_0_93; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4076 = 7'h5e == index[6:0] ? 1'h0 : dirty_0_94; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4077 = 7'h5f == index[6:0] ? 1'h0 : dirty_0_95; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4078 = 7'h60 == index[6:0] ? 1'h0 : dirty_0_96; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4079 = 7'h61 == index[6:0] ? 1'h0 : dirty_0_97; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4080 = 7'h62 == index[6:0] ? 1'h0 : dirty_0_98; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4081 = 7'h63 == index[6:0] ? 1'h0 : dirty_0_99; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4082 = 7'h64 == index[6:0] ? 1'h0 : dirty_0_100; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4083 = 7'h65 == index[6:0] ? 1'h0 : dirty_0_101; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4084 = 7'h66 == index[6:0] ? 1'h0 : dirty_0_102; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4085 = 7'h67 == index[6:0] ? 1'h0 : dirty_0_103; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4086 = 7'h68 == index[6:0] ? 1'h0 : dirty_0_104; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4087 = 7'h69 == index[6:0] ? 1'h0 : dirty_0_105; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4088 = 7'h6a == index[6:0] ? 1'h0 : dirty_0_106; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4089 = 7'h6b == index[6:0] ? 1'h0 : dirty_0_107; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4090 = 7'h6c == index[6:0] ? 1'h0 : dirty_0_108; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4091 = 7'h6d == index[6:0] ? 1'h0 : dirty_0_109; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4092 = 7'h6e == index[6:0] ? 1'h0 : dirty_0_110; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4093 = 7'h6f == index[6:0] ? 1'h0 : dirty_0_111; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4094 = 7'h70 == index[6:0] ? 1'h0 : dirty_0_112; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4095 = 7'h71 == index[6:0] ? 1'h0 : dirty_0_113; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4096 = 7'h72 == index[6:0] ? 1'h0 : dirty_0_114; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4097 = 7'h73 == index[6:0] ? 1'h0 : dirty_0_115; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4098 = 7'h74 == index[6:0] ? 1'h0 : dirty_0_116; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4099 = 7'h75 == index[6:0] ? 1'h0 : dirty_0_117; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4100 = 7'h76 == index[6:0] ? 1'h0 : dirty_0_118; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4101 = 7'h77 == index[6:0] ? 1'h0 : dirty_0_119; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4102 = 7'h78 == index[6:0] ? 1'h0 : dirty_0_120; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4103 = 7'h79 == index[6:0] ? 1'h0 : dirty_0_121; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4104 = 7'h7a == index[6:0] ? 1'h0 : dirty_0_122; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4105 = 7'h7b == index[6:0] ? 1'h0 : dirty_0_123; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4106 = 7'h7c == index[6:0] ? 1'h0 : dirty_0_124; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4107 = 7'h7d == index[6:0] ? 1'h0 : dirty_0_125; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4108 = 7'h7e == index[6:0] ? 1'h0 : dirty_0_126; // @[d_cache.scala 154:{40,40} 24:26]
  wire  _GEN_4109 = 7'h7f == index[6:0] ? 1'h0 : dirty_0_127; // @[d_cache.scala 154:{40,40} 24:26]
  wire [63:0] _GEN_4622 = _GEN_901 ? _GEN_1160 : write_back_data; // @[d_cache.scala 149:47 150:41 29:34]
  wire [41:0] _GEN_4623 = _GEN_901 ? _write_back_addr_T_3 : {{10'd0}, write_back_addr}; // @[d_cache.scala 149:47 151:41 30:34]
  wire [63:0] _GEN_4624 = _GEN_901 ? _GEN_2574 : _GEN_2574; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4625 = _GEN_901 ? _GEN_2575 : _GEN_2575; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4626 = _GEN_901 ? _GEN_2576 : _GEN_2576; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4627 = _GEN_901 ? _GEN_2577 : _GEN_2577; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4628 = _GEN_901 ? _GEN_2578 : _GEN_2578; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4629 = _GEN_901 ? _GEN_2579 : _GEN_2579; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4630 = _GEN_901 ? _GEN_2580 : _GEN_2580; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4631 = _GEN_901 ? _GEN_2581 : _GEN_2581; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4632 = _GEN_901 ? _GEN_2582 : _GEN_2582; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4633 = _GEN_901 ? _GEN_2583 : _GEN_2583; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4634 = _GEN_901 ? _GEN_2584 : _GEN_2584; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4635 = _GEN_901 ? _GEN_2585 : _GEN_2585; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4636 = _GEN_901 ? _GEN_2586 : _GEN_2586; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4637 = _GEN_901 ? _GEN_2587 : _GEN_2587; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4638 = _GEN_901 ? _GEN_2588 : _GEN_2588; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4639 = _GEN_901 ? _GEN_2589 : _GEN_2589; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4640 = _GEN_901 ? _GEN_2590 : _GEN_2590; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4641 = _GEN_901 ? _GEN_2591 : _GEN_2591; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4642 = _GEN_901 ? _GEN_2592 : _GEN_2592; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4643 = _GEN_901 ? _GEN_2593 : _GEN_2593; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4644 = _GEN_901 ? _GEN_2594 : _GEN_2594; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4645 = _GEN_901 ? _GEN_2595 : _GEN_2595; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4646 = _GEN_901 ? _GEN_2596 : _GEN_2596; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4647 = _GEN_901 ? _GEN_2597 : _GEN_2597; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4648 = _GEN_901 ? _GEN_2598 : _GEN_2598; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4649 = _GEN_901 ? _GEN_2599 : _GEN_2599; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4650 = _GEN_901 ? _GEN_2600 : _GEN_2600; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4651 = _GEN_901 ? _GEN_2601 : _GEN_2601; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4652 = _GEN_901 ? _GEN_2602 : _GEN_2602; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4653 = _GEN_901 ? _GEN_2603 : _GEN_2603; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4654 = _GEN_901 ? _GEN_2604 : _GEN_2604; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4655 = _GEN_901 ? _GEN_2605 : _GEN_2605; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4656 = _GEN_901 ? _GEN_2606 : _GEN_2606; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4657 = _GEN_901 ? _GEN_2607 : _GEN_2607; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4658 = _GEN_901 ? _GEN_2608 : _GEN_2608; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4659 = _GEN_901 ? _GEN_2609 : _GEN_2609; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4660 = _GEN_901 ? _GEN_2610 : _GEN_2610; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4661 = _GEN_901 ? _GEN_2611 : _GEN_2611; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4662 = _GEN_901 ? _GEN_2612 : _GEN_2612; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4663 = _GEN_901 ? _GEN_2613 : _GEN_2613; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4664 = _GEN_901 ? _GEN_2614 : _GEN_2614; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4665 = _GEN_901 ? _GEN_2615 : _GEN_2615; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4666 = _GEN_901 ? _GEN_2616 : _GEN_2616; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4667 = _GEN_901 ? _GEN_2617 : _GEN_2617; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4668 = _GEN_901 ? _GEN_2618 : _GEN_2618; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4669 = _GEN_901 ? _GEN_2619 : _GEN_2619; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4670 = _GEN_901 ? _GEN_2620 : _GEN_2620; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4671 = _GEN_901 ? _GEN_2621 : _GEN_2621; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4672 = _GEN_901 ? _GEN_2622 : _GEN_2622; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4673 = _GEN_901 ? _GEN_2623 : _GEN_2623; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4674 = _GEN_901 ? _GEN_2624 : _GEN_2624; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4675 = _GEN_901 ? _GEN_2625 : _GEN_2625; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4676 = _GEN_901 ? _GEN_2626 : _GEN_2626; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4677 = _GEN_901 ? _GEN_2627 : _GEN_2627; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4678 = _GEN_901 ? _GEN_2628 : _GEN_2628; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4679 = _GEN_901 ? _GEN_2629 : _GEN_2629; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4680 = _GEN_901 ? _GEN_2630 : _GEN_2630; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4681 = _GEN_901 ? _GEN_2631 : _GEN_2631; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4682 = _GEN_901 ? _GEN_2632 : _GEN_2632; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4683 = _GEN_901 ? _GEN_2633 : _GEN_2633; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4684 = _GEN_901 ? _GEN_2634 : _GEN_2634; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4685 = _GEN_901 ? _GEN_2635 : _GEN_2635; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4686 = _GEN_901 ? _GEN_2636 : _GEN_2636; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4687 = _GEN_901 ? _GEN_2637 : _GEN_2637; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4688 = _GEN_901 ? _GEN_2638 : _GEN_2638; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4689 = _GEN_901 ? _GEN_2639 : _GEN_2639; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4690 = _GEN_901 ? _GEN_2640 : _GEN_2640; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4691 = _GEN_901 ? _GEN_2641 : _GEN_2641; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4692 = _GEN_901 ? _GEN_2642 : _GEN_2642; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4693 = _GEN_901 ? _GEN_2643 : _GEN_2643; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4694 = _GEN_901 ? _GEN_2644 : _GEN_2644; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4695 = _GEN_901 ? _GEN_2645 : _GEN_2645; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4696 = _GEN_901 ? _GEN_2646 : _GEN_2646; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4697 = _GEN_901 ? _GEN_2647 : _GEN_2647; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4698 = _GEN_901 ? _GEN_2648 : _GEN_2648; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4699 = _GEN_901 ? _GEN_2649 : _GEN_2649; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4700 = _GEN_901 ? _GEN_2650 : _GEN_2650; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4701 = _GEN_901 ? _GEN_2651 : _GEN_2651; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4702 = _GEN_901 ? _GEN_2652 : _GEN_2652; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4703 = _GEN_901 ? _GEN_2653 : _GEN_2653; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4704 = _GEN_901 ? _GEN_2654 : _GEN_2654; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4705 = _GEN_901 ? _GEN_2655 : _GEN_2655; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4706 = _GEN_901 ? _GEN_2656 : _GEN_2656; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4707 = _GEN_901 ? _GEN_2657 : _GEN_2657; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4708 = _GEN_901 ? _GEN_2658 : _GEN_2658; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4709 = _GEN_901 ? _GEN_2659 : _GEN_2659; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4710 = _GEN_901 ? _GEN_2660 : _GEN_2660; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4711 = _GEN_901 ? _GEN_2661 : _GEN_2661; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4712 = _GEN_901 ? _GEN_2662 : _GEN_2662; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4713 = _GEN_901 ? _GEN_2663 : _GEN_2663; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4714 = _GEN_901 ? _GEN_2664 : _GEN_2664; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4715 = _GEN_901 ? _GEN_2665 : _GEN_2665; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4716 = _GEN_901 ? _GEN_2666 : _GEN_2666; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4717 = _GEN_901 ? _GEN_2667 : _GEN_2667; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4718 = _GEN_901 ? _GEN_2668 : _GEN_2668; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4719 = _GEN_901 ? _GEN_2669 : _GEN_2669; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4720 = _GEN_901 ? _GEN_2670 : _GEN_2670; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4721 = _GEN_901 ? _GEN_2671 : _GEN_2671; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4722 = _GEN_901 ? _GEN_2672 : _GEN_2672; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4723 = _GEN_901 ? _GEN_2673 : _GEN_2673; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4724 = _GEN_901 ? _GEN_2674 : _GEN_2674; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4725 = _GEN_901 ? _GEN_2675 : _GEN_2675; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4726 = _GEN_901 ? _GEN_2676 : _GEN_2676; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4727 = _GEN_901 ? _GEN_2677 : _GEN_2677; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4728 = _GEN_901 ? _GEN_2678 : _GEN_2678; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4729 = _GEN_901 ? _GEN_2679 : _GEN_2679; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4730 = _GEN_901 ? _GEN_2680 : _GEN_2680; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4731 = _GEN_901 ? _GEN_2681 : _GEN_2681; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4732 = _GEN_901 ? _GEN_2682 : _GEN_2682; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4733 = _GEN_901 ? _GEN_2683 : _GEN_2683; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4734 = _GEN_901 ? _GEN_2684 : _GEN_2684; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4735 = _GEN_901 ? _GEN_2685 : _GEN_2685; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4736 = _GEN_901 ? _GEN_2686 : _GEN_2686; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4737 = _GEN_901 ? _GEN_2687 : _GEN_2687; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4738 = _GEN_901 ? _GEN_2688 : _GEN_2688; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4739 = _GEN_901 ? _GEN_2689 : _GEN_2689; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4740 = _GEN_901 ? _GEN_2690 : _GEN_2690; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4741 = _GEN_901 ? _GEN_2691 : _GEN_2691; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4742 = _GEN_901 ? _GEN_2692 : _GEN_2692; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4743 = _GEN_901 ? _GEN_2693 : _GEN_2693; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4744 = _GEN_901 ? _GEN_2694 : _GEN_2694; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4745 = _GEN_901 ? _GEN_2695 : _GEN_2695; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4746 = _GEN_901 ? _GEN_2696 : _GEN_2696; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4747 = _GEN_901 ? _GEN_2697 : _GEN_2697; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4748 = _GEN_901 ? _GEN_2698 : _GEN_2698; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4749 = _GEN_901 ? _GEN_2699 : _GEN_2699; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4750 = _GEN_901 ? _GEN_2700 : _GEN_2700; // @[d_cache.scala 149:47]
  wire [63:0] _GEN_4751 = _GEN_901 ? _GEN_2701 : _GEN_2701; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4752 = _GEN_901 ? _GEN_2702 : _GEN_2702; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4753 = _GEN_901 ? _GEN_2703 : _GEN_2703; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4754 = _GEN_901 ? _GEN_2704 : _GEN_2704; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4755 = _GEN_901 ? _GEN_2705 : _GEN_2705; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4756 = _GEN_901 ? _GEN_2706 : _GEN_2706; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4757 = _GEN_901 ? _GEN_2707 : _GEN_2707; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4758 = _GEN_901 ? _GEN_2708 : _GEN_2708; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4759 = _GEN_901 ? _GEN_2709 : _GEN_2709; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4760 = _GEN_901 ? _GEN_2710 : _GEN_2710; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4761 = _GEN_901 ? _GEN_2711 : _GEN_2711; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4762 = _GEN_901 ? _GEN_2712 : _GEN_2712; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4763 = _GEN_901 ? _GEN_2713 : _GEN_2713; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4764 = _GEN_901 ? _GEN_2714 : _GEN_2714; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4765 = _GEN_901 ? _GEN_2715 : _GEN_2715; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4766 = _GEN_901 ? _GEN_2716 : _GEN_2716; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4767 = _GEN_901 ? _GEN_2717 : _GEN_2717; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4768 = _GEN_901 ? _GEN_2718 : _GEN_2718; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4769 = _GEN_901 ? _GEN_2719 : _GEN_2719; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4770 = _GEN_901 ? _GEN_2720 : _GEN_2720; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4771 = _GEN_901 ? _GEN_2721 : _GEN_2721; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4772 = _GEN_901 ? _GEN_2722 : _GEN_2722; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4773 = _GEN_901 ? _GEN_2723 : _GEN_2723; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4774 = _GEN_901 ? _GEN_2724 : _GEN_2724; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4775 = _GEN_901 ? _GEN_2725 : _GEN_2725; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4776 = _GEN_901 ? _GEN_2726 : _GEN_2726; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4777 = _GEN_901 ? _GEN_2727 : _GEN_2727; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4778 = _GEN_901 ? _GEN_2728 : _GEN_2728; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4779 = _GEN_901 ? _GEN_2729 : _GEN_2729; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4780 = _GEN_901 ? _GEN_2730 : _GEN_2730; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4781 = _GEN_901 ? _GEN_2731 : _GEN_2731; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4782 = _GEN_901 ? _GEN_2732 : _GEN_2732; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4783 = _GEN_901 ? _GEN_2733 : _GEN_2733; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4784 = _GEN_901 ? _GEN_2734 : _GEN_2734; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4785 = _GEN_901 ? _GEN_2735 : _GEN_2735; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4786 = _GEN_901 ? _GEN_2736 : _GEN_2736; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4787 = _GEN_901 ? _GEN_2737 : _GEN_2737; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4788 = _GEN_901 ? _GEN_2738 : _GEN_2738; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4789 = _GEN_901 ? _GEN_2739 : _GEN_2739; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4790 = _GEN_901 ? _GEN_2740 : _GEN_2740; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4791 = _GEN_901 ? _GEN_2741 : _GEN_2741; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4792 = _GEN_901 ? _GEN_2742 : _GEN_2742; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4793 = _GEN_901 ? _GEN_2743 : _GEN_2743; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4794 = _GEN_901 ? _GEN_2744 : _GEN_2744; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4795 = _GEN_901 ? _GEN_2745 : _GEN_2745; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4796 = _GEN_901 ? _GEN_2746 : _GEN_2746; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4797 = _GEN_901 ? _GEN_2747 : _GEN_2747; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4798 = _GEN_901 ? _GEN_2748 : _GEN_2748; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4799 = _GEN_901 ? _GEN_2749 : _GEN_2749; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4800 = _GEN_901 ? _GEN_2750 : _GEN_2750; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4801 = _GEN_901 ? _GEN_2751 : _GEN_2751; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4802 = _GEN_901 ? _GEN_2752 : _GEN_2752; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4803 = _GEN_901 ? _GEN_2753 : _GEN_2753; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4804 = _GEN_901 ? _GEN_2754 : _GEN_2754; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4805 = _GEN_901 ? _GEN_2755 : _GEN_2755; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4806 = _GEN_901 ? _GEN_2756 : _GEN_2756; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4807 = _GEN_901 ? _GEN_2757 : _GEN_2757; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4808 = _GEN_901 ? _GEN_2758 : _GEN_2758; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4809 = _GEN_901 ? _GEN_2759 : _GEN_2759; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4810 = _GEN_901 ? _GEN_2760 : _GEN_2760; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4811 = _GEN_901 ? _GEN_2761 : _GEN_2761; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4812 = _GEN_901 ? _GEN_2762 : _GEN_2762; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4813 = _GEN_901 ? _GEN_2763 : _GEN_2763; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4814 = _GEN_901 ? _GEN_2764 : _GEN_2764; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4815 = _GEN_901 ? _GEN_2765 : _GEN_2765; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4816 = _GEN_901 ? _GEN_2766 : _GEN_2766; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4817 = _GEN_901 ? _GEN_2767 : _GEN_2767; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4818 = _GEN_901 ? _GEN_2768 : _GEN_2768; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4819 = _GEN_901 ? _GEN_2769 : _GEN_2769; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4820 = _GEN_901 ? _GEN_2770 : _GEN_2770; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4821 = _GEN_901 ? _GEN_2771 : _GEN_2771; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4822 = _GEN_901 ? _GEN_2772 : _GEN_2772; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4823 = _GEN_901 ? _GEN_2773 : _GEN_2773; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4824 = _GEN_901 ? _GEN_2774 : _GEN_2774; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4825 = _GEN_901 ? _GEN_2775 : _GEN_2775; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4826 = _GEN_901 ? _GEN_2776 : _GEN_2776; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4827 = _GEN_901 ? _GEN_2777 : _GEN_2777; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4828 = _GEN_901 ? _GEN_2778 : _GEN_2778; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4829 = _GEN_901 ? _GEN_2779 : _GEN_2779; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4830 = _GEN_901 ? _GEN_2780 : _GEN_2780; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4831 = _GEN_901 ? _GEN_2781 : _GEN_2781; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4832 = _GEN_901 ? _GEN_2782 : _GEN_2782; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4833 = _GEN_901 ? _GEN_2783 : _GEN_2783; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4834 = _GEN_901 ? _GEN_2784 : _GEN_2784; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4835 = _GEN_901 ? _GEN_2785 : _GEN_2785; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4836 = _GEN_901 ? _GEN_2786 : _GEN_2786; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4837 = _GEN_901 ? _GEN_2787 : _GEN_2787; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4838 = _GEN_901 ? _GEN_2788 : _GEN_2788; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4839 = _GEN_901 ? _GEN_2789 : _GEN_2789; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4840 = _GEN_901 ? _GEN_2790 : _GEN_2790; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4841 = _GEN_901 ? _GEN_2791 : _GEN_2791; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4842 = _GEN_901 ? _GEN_2792 : _GEN_2792; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4843 = _GEN_901 ? _GEN_2793 : _GEN_2793; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4844 = _GEN_901 ? _GEN_2794 : _GEN_2794; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4845 = _GEN_901 ? _GEN_2795 : _GEN_2795; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4846 = _GEN_901 ? _GEN_2796 : _GEN_2796; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4847 = _GEN_901 ? _GEN_2797 : _GEN_2797; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4848 = _GEN_901 ? _GEN_2798 : _GEN_2798; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4849 = _GEN_901 ? _GEN_2799 : _GEN_2799; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4850 = _GEN_901 ? _GEN_2800 : _GEN_2800; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4851 = _GEN_901 ? _GEN_2801 : _GEN_2801; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4852 = _GEN_901 ? _GEN_2802 : _GEN_2802; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4853 = _GEN_901 ? _GEN_2803 : _GEN_2803; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4854 = _GEN_901 ? _GEN_2804 : _GEN_2804; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4855 = _GEN_901 ? _GEN_2805 : _GEN_2805; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4856 = _GEN_901 ? _GEN_2806 : _GEN_2806; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4857 = _GEN_901 ? _GEN_2807 : _GEN_2807; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4858 = _GEN_901 ? _GEN_2808 : _GEN_2808; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4859 = _GEN_901 ? _GEN_2809 : _GEN_2809; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4860 = _GEN_901 ? _GEN_2810 : _GEN_2810; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4861 = _GEN_901 ? _GEN_2811 : _GEN_2811; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4862 = _GEN_901 ? _GEN_2812 : _GEN_2812; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4863 = _GEN_901 ? _GEN_2813 : _GEN_2813; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4864 = _GEN_901 ? _GEN_2814 : _GEN_2814; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4865 = _GEN_901 ? _GEN_2815 : _GEN_2815; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4866 = _GEN_901 ? _GEN_2816 : _GEN_2816; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4867 = _GEN_901 ? _GEN_2817 : _GEN_2817; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4868 = _GEN_901 ? _GEN_2818 : _GEN_2818; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4869 = _GEN_901 ? _GEN_2819 : _GEN_2819; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4870 = _GEN_901 ? _GEN_2820 : _GEN_2820; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4871 = _GEN_901 ? _GEN_2821 : _GEN_2821; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4872 = _GEN_901 ? _GEN_2822 : _GEN_2822; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4873 = _GEN_901 ? _GEN_2823 : _GEN_2823; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4874 = _GEN_901 ? _GEN_2824 : _GEN_2824; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4875 = _GEN_901 ? _GEN_2825 : _GEN_2825; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4876 = _GEN_901 ? _GEN_2826 : _GEN_2826; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4877 = _GEN_901 ? _GEN_2827 : _GEN_2827; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4878 = _GEN_901 ? _GEN_2828 : _GEN_2828; // @[d_cache.scala 149:47]
  wire [31:0] _GEN_4879 = _GEN_901 ? _GEN_2829 : _GEN_2829; // @[d_cache.scala 149:47]
  wire  _GEN_4880 = _GEN_901 ? _GEN_3982 : dirty_0_0; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4881 = _GEN_901 ? _GEN_3983 : dirty_0_1; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4882 = _GEN_901 ? _GEN_3984 : dirty_0_2; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4883 = _GEN_901 ? _GEN_3985 : dirty_0_3; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4884 = _GEN_901 ? _GEN_3986 : dirty_0_4; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4885 = _GEN_901 ? _GEN_3987 : dirty_0_5; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4886 = _GEN_901 ? _GEN_3988 : dirty_0_6; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4887 = _GEN_901 ? _GEN_3989 : dirty_0_7; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4888 = _GEN_901 ? _GEN_3990 : dirty_0_8; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4889 = _GEN_901 ? _GEN_3991 : dirty_0_9; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4890 = _GEN_901 ? _GEN_3992 : dirty_0_10; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4891 = _GEN_901 ? _GEN_3993 : dirty_0_11; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4892 = _GEN_901 ? _GEN_3994 : dirty_0_12; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4893 = _GEN_901 ? _GEN_3995 : dirty_0_13; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4894 = _GEN_901 ? _GEN_3996 : dirty_0_14; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4895 = _GEN_901 ? _GEN_3997 : dirty_0_15; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4896 = _GEN_901 ? _GEN_3998 : dirty_0_16; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4897 = _GEN_901 ? _GEN_3999 : dirty_0_17; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4898 = _GEN_901 ? _GEN_4000 : dirty_0_18; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4899 = _GEN_901 ? _GEN_4001 : dirty_0_19; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4900 = _GEN_901 ? _GEN_4002 : dirty_0_20; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4901 = _GEN_901 ? _GEN_4003 : dirty_0_21; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4902 = _GEN_901 ? _GEN_4004 : dirty_0_22; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4903 = _GEN_901 ? _GEN_4005 : dirty_0_23; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4904 = _GEN_901 ? _GEN_4006 : dirty_0_24; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4905 = _GEN_901 ? _GEN_4007 : dirty_0_25; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4906 = _GEN_901 ? _GEN_4008 : dirty_0_26; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4907 = _GEN_901 ? _GEN_4009 : dirty_0_27; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4908 = _GEN_901 ? _GEN_4010 : dirty_0_28; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4909 = _GEN_901 ? _GEN_4011 : dirty_0_29; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4910 = _GEN_901 ? _GEN_4012 : dirty_0_30; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4911 = _GEN_901 ? _GEN_4013 : dirty_0_31; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4912 = _GEN_901 ? _GEN_4014 : dirty_0_32; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4913 = _GEN_901 ? _GEN_4015 : dirty_0_33; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4914 = _GEN_901 ? _GEN_4016 : dirty_0_34; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4915 = _GEN_901 ? _GEN_4017 : dirty_0_35; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4916 = _GEN_901 ? _GEN_4018 : dirty_0_36; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4917 = _GEN_901 ? _GEN_4019 : dirty_0_37; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4918 = _GEN_901 ? _GEN_4020 : dirty_0_38; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4919 = _GEN_901 ? _GEN_4021 : dirty_0_39; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4920 = _GEN_901 ? _GEN_4022 : dirty_0_40; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4921 = _GEN_901 ? _GEN_4023 : dirty_0_41; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4922 = _GEN_901 ? _GEN_4024 : dirty_0_42; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4923 = _GEN_901 ? _GEN_4025 : dirty_0_43; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4924 = _GEN_901 ? _GEN_4026 : dirty_0_44; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4925 = _GEN_901 ? _GEN_4027 : dirty_0_45; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4926 = _GEN_901 ? _GEN_4028 : dirty_0_46; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4927 = _GEN_901 ? _GEN_4029 : dirty_0_47; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4928 = _GEN_901 ? _GEN_4030 : dirty_0_48; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4929 = _GEN_901 ? _GEN_4031 : dirty_0_49; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4930 = _GEN_901 ? _GEN_4032 : dirty_0_50; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4931 = _GEN_901 ? _GEN_4033 : dirty_0_51; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4932 = _GEN_901 ? _GEN_4034 : dirty_0_52; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4933 = _GEN_901 ? _GEN_4035 : dirty_0_53; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4934 = _GEN_901 ? _GEN_4036 : dirty_0_54; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4935 = _GEN_901 ? _GEN_4037 : dirty_0_55; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4936 = _GEN_901 ? _GEN_4038 : dirty_0_56; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4937 = _GEN_901 ? _GEN_4039 : dirty_0_57; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4938 = _GEN_901 ? _GEN_4040 : dirty_0_58; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4939 = _GEN_901 ? _GEN_4041 : dirty_0_59; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4940 = _GEN_901 ? _GEN_4042 : dirty_0_60; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4941 = _GEN_901 ? _GEN_4043 : dirty_0_61; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4942 = _GEN_901 ? _GEN_4044 : dirty_0_62; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4943 = _GEN_901 ? _GEN_4045 : dirty_0_63; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4944 = _GEN_901 ? _GEN_4046 : dirty_0_64; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4945 = _GEN_901 ? _GEN_4047 : dirty_0_65; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4946 = _GEN_901 ? _GEN_4048 : dirty_0_66; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4947 = _GEN_901 ? _GEN_4049 : dirty_0_67; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4948 = _GEN_901 ? _GEN_4050 : dirty_0_68; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4949 = _GEN_901 ? _GEN_4051 : dirty_0_69; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4950 = _GEN_901 ? _GEN_4052 : dirty_0_70; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4951 = _GEN_901 ? _GEN_4053 : dirty_0_71; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4952 = _GEN_901 ? _GEN_4054 : dirty_0_72; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4953 = _GEN_901 ? _GEN_4055 : dirty_0_73; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4954 = _GEN_901 ? _GEN_4056 : dirty_0_74; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4955 = _GEN_901 ? _GEN_4057 : dirty_0_75; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4956 = _GEN_901 ? _GEN_4058 : dirty_0_76; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4957 = _GEN_901 ? _GEN_4059 : dirty_0_77; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4958 = _GEN_901 ? _GEN_4060 : dirty_0_78; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4959 = _GEN_901 ? _GEN_4061 : dirty_0_79; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4960 = _GEN_901 ? _GEN_4062 : dirty_0_80; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4961 = _GEN_901 ? _GEN_4063 : dirty_0_81; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4962 = _GEN_901 ? _GEN_4064 : dirty_0_82; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4963 = _GEN_901 ? _GEN_4065 : dirty_0_83; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4964 = _GEN_901 ? _GEN_4066 : dirty_0_84; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4965 = _GEN_901 ? _GEN_4067 : dirty_0_85; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4966 = _GEN_901 ? _GEN_4068 : dirty_0_86; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4967 = _GEN_901 ? _GEN_4069 : dirty_0_87; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4968 = _GEN_901 ? _GEN_4070 : dirty_0_88; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4969 = _GEN_901 ? _GEN_4071 : dirty_0_89; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4970 = _GEN_901 ? _GEN_4072 : dirty_0_90; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4971 = _GEN_901 ? _GEN_4073 : dirty_0_91; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4972 = _GEN_901 ? _GEN_4074 : dirty_0_92; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4973 = _GEN_901 ? _GEN_4075 : dirty_0_93; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4974 = _GEN_901 ? _GEN_4076 : dirty_0_94; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4975 = _GEN_901 ? _GEN_4077 : dirty_0_95; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4976 = _GEN_901 ? _GEN_4078 : dirty_0_96; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4977 = _GEN_901 ? _GEN_4079 : dirty_0_97; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4978 = _GEN_901 ? _GEN_4080 : dirty_0_98; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4979 = _GEN_901 ? _GEN_4081 : dirty_0_99; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4980 = _GEN_901 ? _GEN_4082 : dirty_0_100; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4981 = _GEN_901 ? _GEN_4083 : dirty_0_101; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4982 = _GEN_901 ? _GEN_4084 : dirty_0_102; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4983 = _GEN_901 ? _GEN_4085 : dirty_0_103; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4984 = _GEN_901 ? _GEN_4086 : dirty_0_104; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4985 = _GEN_901 ? _GEN_4087 : dirty_0_105; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4986 = _GEN_901 ? _GEN_4088 : dirty_0_106; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4987 = _GEN_901 ? _GEN_4089 : dirty_0_107; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4988 = _GEN_901 ? _GEN_4090 : dirty_0_108; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4989 = _GEN_901 ? _GEN_4091 : dirty_0_109; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4990 = _GEN_901 ? _GEN_4092 : dirty_0_110; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4991 = _GEN_901 ? _GEN_4093 : dirty_0_111; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4992 = _GEN_901 ? _GEN_4094 : dirty_0_112; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4993 = _GEN_901 ? _GEN_4095 : dirty_0_113; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4994 = _GEN_901 ? _GEN_4096 : dirty_0_114; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4995 = _GEN_901 ? _GEN_4097 : dirty_0_115; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4996 = _GEN_901 ? _GEN_4098 : dirty_0_116; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4997 = _GEN_901 ? _GEN_4099 : dirty_0_117; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4998 = _GEN_901 ? _GEN_4100 : dirty_0_118; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_4999 = _GEN_901 ? _GEN_4101 : dirty_0_119; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_5000 = _GEN_901 ? _GEN_4102 : dirty_0_120; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_5001 = _GEN_901 ? _GEN_4103 : dirty_0_121; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_5002 = _GEN_901 ? _GEN_4104 : dirty_0_122; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_5003 = _GEN_901 ? _GEN_4105 : dirty_0_123; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_5004 = _GEN_901 ? _GEN_4106 : dirty_0_124; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_5005 = _GEN_901 ? _GEN_4107 : dirty_0_125; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_5006 = _GEN_901 ? _GEN_4108 : dirty_0_126; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_5007 = _GEN_901 ? _GEN_4109 : dirty_0_127; // @[d_cache.scala 149:47 24:26]
  wire  _GEN_5008 = _GEN_901 ? _GEN_2830 : _GEN_2830; // @[d_cache.scala 149:47]
  wire  _GEN_5009 = _GEN_901 ? _GEN_2831 : _GEN_2831; // @[d_cache.scala 149:47]
  wire  _GEN_5010 = _GEN_901 ? _GEN_2832 : _GEN_2832; // @[d_cache.scala 149:47]
  wire  _GEN_5011 = _GEN_901 ? _GEN_2833 : _GEN_2833; // @[d_cache.scala 149:47]
  wire  _GEN_5012 = _GEN_901 ? _GEN_2834 : _GEN_2834; // @[d_cache.scala 149:47]
  wire  _GEN_5013 = _GEN_901 ? _GEN_2835 : _GEN_2835; // @[d_cache.scala 149:47]
  wire  _GEN_5014 = _GEN_901 ? _GEN_2836 : _GEN_2836; // @[d_cache.scala 149:47]
  wire  _GEN_5015 = _GEN_901 ? _GEN_2837 : _GEN_2837; // @[d_cache.scala 149:47]
  wire  _GEN_5016 = _GEN_901 ? _GEN_2838 : _GEN_2838; // @[d_cache.scala 149:47]
  wire  _GEN_5017 = _GEN_901 ? _GEN_2839 : _GEN_2839; // @[d_cache.scala 149:47]
  wire  _GEN_5018 = _GEN_901 ? _GEN_2840 : _GEN_2840; // @[d_cache.scala 149:47]
  wire  _GEN_5019 = _GEN_901 ? _GEN_2841 : _GEN_2841; // @[d_cache.scala 149:47]
  wire  _GEN_5020 = _GEN_901 ? _GEN_2842 : _GEN_2842; // @[d_cache.scala 149:47]
  wire  _GEN_5021 = _GEN_901 ? _GEN_2843 : _GEN_2843; // @[d_cache.scala 149:47]
  wire  _GEN_5022 = _GEN_901 ? _GEN_2844 : _GEN_2844; // @[d_cache.scala 149:47]
  wire  _GEN_5023 = _GEN_901 ? _GEN_2845 : _GEN_2845; // @[d_cache.scala 149:47]
  wire  _GEN_5024 = _GEN_901 ? _GEN_2846 : _GEN_2846; // @[d_cache.scala 149:47]
  wire  _GEN_5025 = _GEN_901 ? _GEN_2847 : _GEN_2847; // @[d_cache.scala 149:47]
  wire  _GEN_5026 = _GEN_901 ? _GEN_2848 : _GEN_2848; // @[d_cache.scala 149:47]
  wire  _GEN_5027 = _GEN_901 ? _GEN_2849 : _GEN_2849; // @[d_cache.scala 149:47]
  wire  _GEN_5028 = _GEN_901 ? _GEN_2850 : _GEN_2850; // @[d_cache.scala 149:47]
  wire  _GEN_5029 = _GEN_901 ? _GEN_2851 : _GEN_2851; // @[d_cache.scala 149:47]
  wire  _GEN_5030 = _GEN_901 ? _GEN_2852 : _GEN_2852; // @[d_cache.scala 149:47]
  wire  _GEN_5031 = _GEN_901 ? _GEN_2853 : _GEN_2853; // @[d_cache.scala 149:47]
  wire  _GEN_5032 = _GEN_901 ? _GEN_2854 : _GEN_2854; // @[d_cache.scala 149:47]
  wire  _GEN_5033 = _GEN_901 ? _GEN_2855 : _GEN_2855; // @[d_cache.scala 149:47]
  wire  _GEN_5034 = _GEN_901 ? _GEN_2856 : _GEN_2856; // @[d_cache.scala 149:47]
  wire  _GEN_5035 = _GEN_901 ? _GEN_2857 : _GEN_2857; // @[d_cache.scala 149:47]
  wire  _GEN_5036 = _GEN_901 ? _GEN_2858 : _GEN_2858; // @[d_cache.scala 149:47]
  wire  _GEN_5037 = _GEN_901 ? _GEN_2859 : _GEN_2859; // @[d_cache.scala 149:47]
  wire  _GEN_5038 = _GEN_901 ? _GEN_2860 : _GEN_2860; // @[d_cache.scala 149:47]
  wire  _GEN_5039 = _GEN_901 ? _GEN_2861 : _GEN_2861; // @[d_cache.scala 149:47]
  wire  _GEN_5040 = _GEN_901 ? _GEN_2862 : _GEN_2862; // @[d_cache.scala 149:47]
  wire  _GEN_5041 = _GEN_901 ? _GEN_2863 : _GEN_2863; // @[d_cache.scala 149:47]
  wire  _GEN_5042 = _GEN_901 ? _GEN_2864 : _GEN_2864; // @[d_cache.scala 149:47]
  wire  _GEN_5043 = _GEN_901 ? _GEN_2865 : _GEN_2865; // @[d_cache.scala 149:47]
  wire  _GEN_5044 = _GEN_901 ? _GEN_2866 : _GEN_2866; // @[d_cache.scala 149:47]
  wire  _GEN_5045 = _GEN_901 ? _GEN_2867 : _GEN_2867; // @[d_cache.scala 149:47]
  wire  _GEN_5046 = _GEN_901 ? _GEN_2868 : _GEN_2868; // @[d_cache.scala 149:47]
  wire  _GEN_5047 = _GEN_901 ? _GEN_2869 : _GEN_2869; // @[d_cache.scala 149:47]
  wire  _GEN_5048 = _GEN_901 ? _GEN_2870 : _GEN_2870; // @[d_cache.scala 149:47]
  wire  _GEN_5049 = _GEN_901 ? _GEN_2871 : _GEN_2871; // @[d_cache.scala 149:47]
  wire  _GEN_5050 = _GEN_901 ? _GEN_2872 : _GEN_2872; // @[d_cache.scala 149:47]
  wire  _GEN_5051 = _GEN_901 ? _GEN_2873 : _GEN_2873; // @[d_cache.scala 149:47]
  wire  _GEN_5052 = _GEN_901 ? _GEN_2874 : _GEN_2874; // @[d_cache.scala 149:47]
  wire  _GEN_5053 = _GEN_901 ? _GEN_2875 : _GEN_2875; // @[d_cache.scala 149:47]
  wire  _GEN_5054 = _GEN_901 ? _GEN_2876 : _GEN_2876; // @[d_cache.scala 149:47]
  wire  _GEN_5055 = _GEN_901 ? _GEN_2877 : _GEN_2877; // @[d_cache.scala 149:47]
  wire  _GEN_5056 = _GEN_901 ? _GEN_2878 : _GEN_2878; // @[d_cache.scala 149:47]
  wire  _GEN_5057 = _GEN_901 ? _GEN_2879 : _GEN_2879; // @[d_cache.scala 149:47]
  wire  _GEN_5058 = _GEN_901 ? _GEN_2880 : _GEN_2880; // @[d_cache.scala 149:47]
  wire  _GEN_5059 = _GEN_901 ? _GEN_2881 : _GEN_2881; // @[d_cache.scala 149:47]
  wire  _GEN_5060 = _GEN_901 ? _GEN_2882 : _GEN_2882; // @[d_cache.scala 149:47]
  wire  _GEN_5061 = _GEN_901 ? _GEN_2883 : _GEN_2883; // @[d_cache.scala 149:47]
  wire  _GEN_5062 = _GEN_901 ? _GEN_2884 : _GEN_2884; // @[d_cache.scala 149:47]
  wire  _GEN_5063 = _GEN_901 ? _GEN_2885 : _GEN_2885; // @[d_cache.scala 149:47]
  wire  _GEN_5064 = _GEN_901 ? _GEN_2886 : _GEN_2886; // @[d_cache.scala 149:47]
  wire  _GEN_5065 = _GEN_901 ? _GEN_2887 : _GEN_2887; // @[d_cache.scala 149:47]
  wire  _GEN_5066 = _GEN_901 ? _GEN_2888 : _GEN_2888; // @[d_cache.scala 149:47]
  wire  _GEN_5067 = _GEN_901 ? _GEN_2889 : _GEN_2889; // @[d_cache.scala 149:47]
  wire  _GEN_5068 = _GEN_901 ? _GEN_2890 : _GEN_2890; // @[d_cache.scala 149:47]
  wire  _GEN_5069 = _GEN_901 ? _GEN_2891 : _GEN_2891; // @[d_cache.scala 149:47]
  wire  _GEN_5070 = _GEN_901 ? _GEN_2892 : _GEN_2892; // @[d_cache.scala 149:47]
  wire  _GEN_5071 = _GEN_901 ? _GEN_2893 : _GEN_2893; // @[d_cache.scala 149:47]
  wire  _GEN_5072 = _GEN_901 ? _GEN_2894 : _GEN_2894; // @[d_cache.scala 149:47]
  wire  _GEN_5073 = _GEN_901 ? _GEN_2895 : _GEN_2895; // @[d_cache.scala 149:47]
  wire  _GEN_5074 = _GEN_901 ? _GEN_2896 : _GEN_2896; // @[d_cache.scala 149:47]
  wire  _GEN_5075 = _GEN_901 ? _GEN_2897 : _GEN_2897; // @[d_cache.scala 149:47]
  wire  _GEN_5076 = _GEN_901 ? _GEN_2898 : _GEN_2898; // @[d_cache.scala 149:47]
  wire  _GEN_5077 = _GEN_901 ? _GEN_2899 : _GEN_2899; // @[d_cache.scala 149:47]
  wire  _GEN_5078 = _GEN_901 ? _GEN_2900 : _GEN_2900; // @[d_cache.scala 149:47]
  wire  _GEN_5079 = _GEN_901 ? _GEN_2901 : _GEN_2901; // @[d_cache.scala 149:47]
  wire  _GEN_5080 = _GEN_901 ? _GEN_2902 : _GEN_2902; // @[d_cache.scala 149:47]
  wire  _GEN_5081 = _GEN_901 ? _GEN_2903 : _GEN_2903; // @[d_cache.scala 149:47]
  wire  _GEN_5082 = _GEN_901 ? _GEN_2904 : _GEN_2904; // @[d_cache.scala 149:47]
  wire  _GEN_5083 = _GEN_901 ? _GEN_2905 : _GEN_2905; // @[d_cache.scala 149:47]
  wire  _GEN_5084 = _GEN_901 ? _GEN_2906 : _GEN_2906; // @[d_cache.scala 149:47]
  wire  _GEN_5085 = _GEN_901 ? _GEN_2907 : _GEN_2907; // @[d_cache.scala 149:47]
  wire  _GEN_5086 = _GEN_901 ? _GEN_2908 : _GEN_2908; // @[d_cache.scala 149:47]
  wire  _GEN_5087 = _GEN_901 ? _GEN_2909 : _GEN_2909; // @[d_cache.scala 149:47]
  wire  _GEN_5088 = _GEN_901 ? _GEN_2910 : _GEN_2910; // @[d_cache.scala 149:47]
  wire  _GEN_5089 = _GEN_901 ? _GEN_2911 : _GEN_2911; // @[d_cache.scala 149:47]
  wire  _GEN_5090 = _GEN_901 ? _GEN_2912 : _GEN_2912; // @[d_cache.scala 149:47]
  wire  _GEN_5091 = _GEN_901 ? _GEN_2913 : _GEN_2913; // @[d_cache.scala 149:47]
  wire  _GEN_5092 = _GEN_901 ? _GEN_2914 : _GEN_2914; // @[d_cache.scala 149:47]
  wire  _GEN_5093 = _GEN_901 ? _GEN_2915 : _GEN_2915; // @[d_cache.scala 149:47]
  wire  _GEN_5094 = _GEN_901 ? _GEN_2916 : _GEN_2916; // @[d_cache.scala 149:47]
  wire  _GEN_5095 = _GEN_901 ? _GEN_2917 : _GEN_2917; // @[d_cache.scala 149:47]
  wire  _GEN_5096 = _GEN_901 ? _GEN_2918 : _GEN_2918; // @[d_cache.scala 149:47]
  wire  _GEN_5097 = _GEN_901 ? _GEN_2919 : _GEN_2919; // @[d_cache.scala 149:47]
  wire  _GEN_5098 = _GEN_901 ? _GEN_2920 : _GEN_2920; // @[d_cache.scala 149:47]
  wire  _GEN_5099 = _GEN_901 ? _GEN_2921 : _GEN_2921; // @[d_cache.scala 149:47]
  wire  _GEN_5100 = _GEN_901 ? _GEN_2922 : _GEN_2922; // @[d_cache.scala 149:47]
  wire  _GEN_5101 = _GEN_901 ? _GEN_2923 : _GEN_2923; // @[d_cache.scala 149:47]
  wire  _GEN_5102 = _GEN_901 ? _GEN_2924 : _GEN_2924; // @[d_cache.scala 149:47]
  wire  _GEN_5103 = _GEN_901 ? _GEN_2925 : _GEN_2925; // @[d_cache.scala 149:47]
  wire  _GEN_5104 = _GEN_901 ? _GEN_2926 : _GEN_2926; // @[d_cache.scala 149:47]
  wire  _GEN_5105 = _GEN_901 ? _GEN_2927 : _GEN_2927; // @[d_cache.scala 149:47]
  wire  _GEN_5106 = _GEN_901 ? _GEN_2928 : _GEN_2928; // @[d_cache.scala 149:47]
  wire  _GEN_5107 = _GEN_901 ? _GEN_2929 : _GEN_2929; // @[d_cache.scala 149:47]
  wire  _GEN_5108 = _GEN_901 ? _GEN_2930 : _GEN_2930; // @[d_cache.scala 149:47]
  wire  _GEN_5109 = _GEN_901 ? _GEN_2931 : _GEN_2931; // @[d_cache.scala 149:47]
  wire  _GEN_5110 = _GEN_901 ? _GEN_2932 : _GEN_2932; // @[d_cache.scala 149:47]
  wire  _GEN_5111 = _GEN_901 ? _GEN_2933 : _GEN_2933; // @[d_cache.scala 149:47]
  wire  _GEN_5112 = _GEN_901 ? _GEN_2934 : _GEN_2934; // @[d_cache.scala 149:47]
  wire  _GEN_5113 = _GEN_901 ? _GEN_2935 : _GEN_2935; // @[d_cache.scala 149:47]
  wire  _GEN_5114 = _GEN_901 ? _GEN_2936 : _GEN_2936; // @[d_cache.scala 149:47]
  wire  _GEN_5115 = _GEN_901 ? _GEN_2937 : _GEN_2937; // @[d_cache.scala 149:47]
  wire  _GEN_5116 = _GEN_901 ? _GEN_2938 : _GEN_2938; // @[d_cache.scala 149:47]
  wire  _GEN_5117 = _GEN_901 ? _GEN_2939 : _GEN_2939; // @[d_cache.scala 149:47]
  wire  _GEN_5118 = _GEN_901 ? _GEN_2940 : _GEN_2940; // @[d_cache.scala 149:47]
  wire  _GEN_5119 = _GEN_901 ? _GEN_2941 : _GEN_2941; // @[d_cache.scala 149:47]
  wire  _GEN_5120 = _GEN_901 ? _GEN_2942 : _GEN_2942; // @[d_cache.scala 149:47]
  wire  _GEN_5121 = _GEN_901 ? _GEN_2943 : _GEN_2943; // @[d_cache.scala 149:47]
  wire  _GEN_5122 = _GEN_901 ? _GEN_2944 : _GEN_2944; // @[d_cache.scala 149:47]
  wire  _GEN_5123 = _GEN_901 ? _GEN_2945 : _GEN_2945; // @[d_cache.scala 149:47]
  wire  _GEN_5124 = _GEN_901 ? _GEN_2946 : _GEN_2946; // @[d_cache.scala 149:47]
  wire  _GEN_5125 = _GEN_901 ? _GEN_2947 : _GEN_2947; // @[d_cache.scala 149:47]
  wire  _GEN_5126 = _GEN_901 ? _GEN_2948 : _GEN_2948; // @[d_cache.scala 149:47]
  wire  _GEN_5127 = _GEN_901 ? _GEN_2949 : _GEN_2949; // @[d_cache.scala 149:47]
  wire  _GEN_5128 = _GEN_901 ? _GEN_2950 : _GEN_2950; // @[d_cache.scala 149:47]
  wire  _GEN_5129 = _GEN_901 ? _GEN_2951 : _GEN_2951; // @[d_cache.scala 149:47]
  wire  _GEN_5130 = _GEN_901 ? _GEN_2952 : _GEN_2952; // @[d_cache.scala 149:47]
  wire  _GEN_5131 = _GEN_901 ? _GEN_2953 : _GEN_2953; // @[d_cache.scala 149:47]
  wire  _GEN_5132 = _GEN_901 ? _GEN_2954 : _GEN_2954; // @[d_cache.scala 149:47]
  wire  _GEN_5133 = _GEN_901 ? _GEN_2955 : _GEN_2955; // @[d_cache.scala 149:47]
  wire  _GEN_5134 = _GEN_901 ? _GEN_2956 : _GEN_2956; // @[d_cache.scala 149:47]
  wire  _GEN_5135 = _GEN_901 ? _GEN_2957 : _GEN_2957; // @[d_cache.scala 149:47]
  wire [2:0] _GEN_5136 = _GEN_901 ? 3'h6 : 3'h7; // @[d_cache.scala 149:47 156:31 159:31]
  wire [63:0] _GEN_5267 = 7'h1 == index[6:0] ? ram_1_1 : ram_1_0; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5268 = 7'h2 == index[6:0] ? ram_1_2 : _GEN_5267; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5269 = 7'h3 == index[6:0] ? ram_1_3 : _GEN_5268; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5270 = 7'h4 == index[6:0] ? ram_1_4 : _GEN_5269; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5271 = 7'h5 == index[6:0] ? ram_1_5 : _GEN_5270; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5272 = 7'h6 == index[6:0] ? ram_1_6 : _GEN_5271; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5273 = 7'h7 == index[6:0] ? ram_1_7 : _GEN_5272; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5274 = 7'h8 == index[6:0] ? ram_1_8 : _GEN_5273; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5275 = 7'h9 == index[6:0] ? ram_1_9 : _GEN_5274; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5276 = 7'ha == index[6:0] ? ram_1_10 : _GEN_5275; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5277 = 7'hb == index[6:0] ? ram_1_11 : _GEN_5276; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5278 = 7'hc == index[6:0] ? ram_1_12 : _GEN_5277; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5279 = 7'hd == index[6:0] ? ram_1_13 : _GEN_5278; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5280 = 7'he == index[6:0] ? ram_1_14 : _GEN_5279; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5281 = 7'hf == index[6:0] ? ram_1_15 : _GEN_5280; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5282 = 7'h10 == index[6:0] ? ram_1_16 : _GEN_5281; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5283 = 7'h11 == index[6:0] ? ram_1_17 : _GEN_5282; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5284 = 7'h12 == index[6:0] ? ram_1_18 : _GEN_5283; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5285 = 7'h13 == index[6:0] ? ram_1_19 : _GEN_5284; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5286 = 7'h14 == index[6:0] ? ram_1_20 : _GEN_5285; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5287 = 7'h15 == index[6:0] ? ram_1_21 : _GEN_5286; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5288 = 7'h16 == index[6:0] ? ram_1_22 : _GEN_5287; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5289 = 7'h17 == index[6:0] ? ram_1_23 : _GEN_5288; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5290 = 7'h18 == index[6:0] ? ram_1_24 : _GEN_5289; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5291 = 7'h19 == index[6:0] ? ram_1_25 : _GEN_5290; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5292 = 7'h1a == index[6:0] ? ram_1_26 : _GEN_5291; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5293 = 7'h1b == index[6:0] ? ram_1_27 : _GEN_5292; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5294 = 7'h1c == index[6:0] ? ram_1_28 : _GEN_5293; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5295 = 7'h1d == index[6:0] ? ram_1_29 : _GEN_5294; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5296 = 7'h1e == index[6:0] ? ram_1_30 : _GEN_5295; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5297 = 7'h1f == index[6:0] ? ram_1_31 : _GEN_5296; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5298 = 7'h20 == index[6:0] ? ram_1_32 : _GEN_5297; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5299 = 7'h21 == index[6:0] ? ram_1_33 : _GEN_5298; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5300 = 7'h22 == index[6:0] ? ram_1_34 : _GEN_5299; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5301 = 7'h23 == index[6:0] ? ram_1_35 : _GEN_5300; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5302 = 7'h24 == index[6:0] ? ram_1_36 : _GEN_5301; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5303 = 7'h25 == index[6:0] ? ram_1_37 : _GEN_5302; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5304 = 7'h26 == index[6:0] ? ram_1_38 : _GEN_5303; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5305 = 7'h27 == index[6:0] ? ram_1_39 : _GEN_5304; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5306 = 7'h28 == index[6:0] ? ram_1_40 : _GEN_5305; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5307 = 7'h29 == index[6:0] ? ram_1_41 : _GEN_5306; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5308 = 7'h2a == index[6:0] ? ram_1_42 : _GEN_5307; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5309 = 7'h2b == index[6:0] ? ram_1_43 : _GEN_5308; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5310 = 7'h2c == index[6:0] ? ram_1_44 : _GEN_5309; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5311 = 7'h2d == index[6:0] ? ram_1_45 : _GEN_5310; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5312 = 7'h2e == index[6:0] ? ram_1_46 : _GEN_5311; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5313 = 7'h2f == index[6:0] ? ram_1_47 : _GEN_5312; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5314 = 7'h30 == index[6:0] ? ram_1_48 : _GEN_5313; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5315 = 7'h31 == index[6:0] ? ram_1_49 : _GEN_5314; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5316 = 7'h32 == index[6:0] ? ram_1_50 : _GEN_5315; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5317 = 7'h33 == index[6:0] ? ram_1_51 : _GEN_5316; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5318 = 7'h34 == index[6:0] ? ram_1_52 : _GEN_5317; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5319 = 7'h35 == index[6:0] ? ram_1_53 : _GEN_5318; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5320 = 7'h36 == index[6:0] ? ram_1_54 : _GEN_5319; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5321 = 7'h37 == index[6:0] ? ram_1_55 : _GEN_5320; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5322 = 7'h38 == index[6:0] ? ram_1_56 : _GEN_5321; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5323 = 7'h39 == index[6:0] ? ram_1_57 : _GEN_5322; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5324 = 7'h3a == index[6:0] ? ram_1_58 : _GEN_5323; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5325 = 7'h3b == index[6:0] ? ram_1_59 : _GEN_5324; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5326 = 7'h3c == index[6:0] ? ram_1_60 : _GEN_5325; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5327 = 7'h3d == index[6:0] ? ram_1_61 : _GEN_5326; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5328 = 7'h3e == index[6:0] ? ram_1_62 : _GEN_5327; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5329 = 7'h3f == index[6:0] ? ram_1_63 : _GEN_5328; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5330 = 7'h40 == index[6:0] ? ram_1_64 : _GEN_5329; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5331 = 7'h41 == index[6:0] ? ram_1_65 : _GEN_5330; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5332 = 7'h42 == index[6:0] ? ram_1_66 : _GEN_5331; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5333 = 7'h43 == index[6:0] ? ram_1_67 : _GEN_5332; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5334 = 7'h44 == index[6:0] ? ram_1_68 : _GEN_5333; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5335 = 7'h45 == index[6:0] ? ram_1_69 : _GEN_5334; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5336 = 7'h46 == index[6:0] ? ram_1_70 : _GEN_5335; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5337 = 7'h47 == index[6:0] ? ram_1_71 : _GEN_5336; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5338 = 7'h48 == index[6:0] ? ram_1_72 : _GEN_5337; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5339 = 7'h49 == index[6:0] ? ram_1_73 : _GEN_5338; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5340 = 7'h4a == index[6:0] ? ram_1_74 : _GEN_5339; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5341 = 7'h4b == index[6:0] ? ram_1_75 : _GEN_5340; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5342 = 7'h4c == index[6:0] ? ram_1_76 : _GEN_5341; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5343 = 7'h4d == index[6:0] ? ram_1_77 : _GEN_5342; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5344 = 7'h4e == index[6:0] ? ram_1_78 : _GEN_5343; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5345 = 7'h4f == index[6:0] ? ram_1_79 : _GEN_5344; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5346 = 7'h50 == index[6:0] ? ram_1_80 : _GEN_5345; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5347 = 7'h51 == index[6:0] ? ram_1_81 : _GEN_5346; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5348 = 7'h52 == index[6:0] ? ram_1_82 : _GEN_5347; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5349 = 7'h53 == index[6:0] ? ram_1_83 : _GEN_5348; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5350 = 7'h54 == index[6:0] ? ram_1_84 : _GEN_5349; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5351 = 7'h55 == index[6:0] ? ram_1_85 : _GEN_5350; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5352 = 7'h56 == index[6:0] ? ram_1_86 : _GEN_5351; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5353 = 7'h57 == index[6:0] ? ram_1_87 : _GEN_5352; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5354 = 7'h58 == index[6:0] ? ram_1_88 : _GEN_5353; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5355 = 7'h59 == index[6:0] ? ram_1_89 : _GEN_5354; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5356 = 7'h5a == index[6:0] ? ram_1_90 : _GEN_5355; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5357 = 7'h5b == index[6:0] ? ram_1_91 : _GEN_5356; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5358 = 7'h5c == index[6:0] ? ram_1_92 : _GEN_5357; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5359 = 7'h5d == index[6:0] ? ram_1_93 : _GEN_5358; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5360 = 7'h5e == index[6:0] ? ram_1_94 : _GEN_5359; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5361 = 7'h5f == index[6:0] ? ram_1_95 : _GEN_5360; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5362 = 7'h60 == index[6:0] ? ram_1_96 : _GEN_5361; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5363 = 7'h61 == index[6:0] ? ram_1_97 : _GEN_5362; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5364 = 7'h62 == index[6:0] ? ram_1_98 : _GEN_5363; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5365 = 7'h63 == index[6:0] ? ram_1_99 : _GEN_5364; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5366 = 7'h64 == index[6:0] ? ram_1_100 : _GEN_5365; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5367 = 7'h65 == index[6:0] ? ram_1_101 : _GEN_5366; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5368 = 7'h66 == index[6:0] ? ram_1_102 : _GEN_5367; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5369 = 7'h67 == index[6:0] ? ram_1_103 : _GEN_5368; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5370 = 7'h68 == index[6:0] ? ram_1_104 : _GEN_5369; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5371 = 7'h69 == index[6:0] ? ram_1_105 : _GEN_5370; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5372 = 7'h6a == index[6:0] ? ram_1_106 : _GEN_5371; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5373 = 7'h6b == index[6:0] ? ram_1_107 : _GEN_5372; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5374 = 7'h6c == index[6:0] ? ram_1_108 : _GEN_5373; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5375 = 7'h6d == index[6:0] ? ram_1_109 : _GEN_5374; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5376 = 7'h6e == index[6:0] ? ram_1_110 : _GEN_5375; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5377 = 7'h6f == index[6:0] ? ram_1_111 : _GEN_5376; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5378 = 7'h70 == index[6:0] ? ram_1_112 : _GEN_5377; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5379 = 7'h71 == index[6:0] ? ram_1_113 : _GEN_5378; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5380 = 7'h72 == index[6:0] ? ram_1_114 : _GEN_5379; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5381 = 7'h73 == index[6:0] ? ram_1_115 : _GEN_5380; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5382 = 7'h74 == index[6:0] ? ram_1_116 : _GEN_5381; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5383 = 7'h75 == index[6:0] ? ram_1_117 : _GEN_5382; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5384 = 7'h76 == index[6:0] ? ram_1_118 : _GEN_5383; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5385 = 7'h77 == index[6:0] ? ram_1_119 : _GEN_5384; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5386 = 7'h78 == index[6:0] ? ram_1_120 : _GEN_5385; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5387 = 7'h79 == index[6:0] ? ram_1_121 : _GEN_5386; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5388 = 7'h7a == index[6:0] ? ram_1_122 : _GEN_5387; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5389 = 7'h7b == index[6:0] ? ram_1_123 : _GEN_5388; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5390 = 7'h7c == index[6:0] ? ram_1_124 : _GEN_5389; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5391 = 7'h7d == index[6:0] ? ram_1_125 : _GEN_5390; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5392 = 7'h7e == index[6:0] ? ram_1_126 : _GEN_5391; // @[d_cache.scala 167:{41,41}]
  wire [63:0] _GEN_5393 = 7'h7f == index[6:0] ? ram_1_127 : _GEN_5392; // @[d_cache.scala 167:{41,41}]
  wire [41:0] _write_back_addr_T_5 = {_GEN_384, 10'h0}; // @[d_cache.scala 168:58]
  wire [41:0] _write_back_addr_T_7 = _write_back_addr_T_5 | _GEN_17319; // @[d_cache.scala 168:65]
  wire  _GEN_5778 = 7'h0 == index[6:0] ? 1'h0 : dirty_1_0; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5779 = 7'h1 == index[6:0] ? 1'h0 : dirty_1_1; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5780 = 7'h2 == index[6:0] ? 1'h0 : dirty_1_2; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5781 = 7'h3 == index[6:0] ? 1'h0 : dirty_1_3; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5782 = 7'h4 == index[6:0] ? 1'h0 : dirty_1_4; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5783 = 7'h5 == index[6:0] ? 1'h0 : dirty_1_5; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5784 = 7'h6 == index[6:0] ? 1'h0 : dirty_1_6; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5785 = 7'h7 == index[6:0] ? 1'h0 : dirty_1_7; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5786 = 7'h8 == index[6:0] ? 1'h0 : dirty_1_8; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5787 = 7'h9 == index[6:0] ? 1'h0 : dirty_1_9; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5788 = 7'ha == index[6:0] ? 1'h0 : dirty_1_10; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5789 = 7'hb == index[6:0] ? 1'h0 : dirty_1_11; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5790 = 7'hc == index[6:0] ? 1'h0 : dirty_1_12; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5791 = 7'hd == index[6:0] ? 1'h0 : dirty_1_13; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5792 = 7'he == index[6:0] ? 1'h0 : dirty_1_14; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5793 = 7'hf == index[6:0] ? 1'h0 : dirty_1_15; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5794 = 7'h10 == index[6:0] ? 1'h0 : dirty_1_16; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5795 = 7'h11 == index[6:0] ? 1'h0 : dirty_1_17; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5796 = 7'h12 == index[6:0] ? 1'h0 : dirty_1_18; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5797 = 7'h13 == index[6:0] ? 1'h0 : dirty_1_19; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5798 = 7'h14 == index[6:0] ? 1'h0 : dirty_1_20; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5799 = 7'h15 == index[6:0] ? 1'h0 : dirty_1_21; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5800 = 7'h16 == index[6:0] ? 1'h0 : dirty_1_22; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5801 = 7'h17 == index[6:0] ? 1'h0 : dirty_1_23; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5802 = 7'h18 == index[6:0] ? 1'h0 : dirty_1_24; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5803 = 7'h19 == index[6:0] ? 1'h0 : dirty_1_25; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5804 = 7'h1a == index[6:0] ? 1'h0 : dirty_1_26; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5805 = 7'h1b == index[6:0] ? 1'h0 : dirty_1_27; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5806 = 7'h1c == index[6:0] ? 1'h0 : dirty_1_28; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5807 = 7'h1d == index[6:0] ? 1'h0 : dirty_1_29; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5808 = 7'h1e == index[6:0] ? 1'h0 : dirty_1_30; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5809 = 7'h1f == index[6:0] ? 1'h0 : dirty_1_31; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5810 = 7'h20 == index[6:0] ? 1'h0 : dirty_1_32; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5811 = 7'h21 == index[6:0] ? 1'h0 : dirty_1_33; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5812 = 7'h22 == index[6:0] ? 1'h0 : dirty_1_34; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5813 = 7'h23 == index[6:0] ? 1'h0 : dirty_1_35; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5814 = 7'h24 == index[6:0] ? 1'h0 : dirty_1_36; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5815 = 7'h25 == index[6:0] ? 1'h0 : dirty_1_37; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5816 = 7'h26 == index[6:0] ? 1'h0 : dirty_1_38; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5817 = 7'h27 == index[6:0] ? 1'h0 : dirty_1_39; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5818 = 7'h28 == index[6:0] ? 1'h0 : dirty_1_40; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5819 = 7'h29 == index[6:0] ? 1'h0 : dirty_1_41; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5820 = 7'h2a == index[6:0] ? 1'h0 : dirty_1_42; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5821 = 7'h2b == index[6:0] ? 1'h0 : dirty_1_43; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5822 = 7'h2c == index[6:0] ? 1'h0 : dirty_1_44; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5823 = 7'h2d == index[6:0] ? 1'h0 : dirty_1_45; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5824 = 7'h2e == index[6:0] ? 1'h0 : dirty_1_46; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5825 = 7'h2f == index[6:0] ? 1'h0 : dirty_1_47; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5826 = 7'h30 == index[6:0] ? 1'h0 : dirty_1_48; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5827 = 7'h31 == index[6:0] ? 1'h0 : dirty_1_49; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5828 = 7'h32 == index[6:0] ? 1'h0 : dirty_1_50; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5829 = 7'h33 == index[6:0] ? 1'h0 : dirty_1_51; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5830 = 7'h34 == index[6:0] ? 1'h0 : dirty_1_52; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5831 = 7'h35 == index[6:0] ? 1'h0 : dirty_1_53; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5832 = 7'h36 == index[6:0] ? 1'h0 : dirty_1_54; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5833 = 7'h37 == index[6:0] ? 1'h0 : dirty_1_55; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5834 = 7'h38 == index[6:0] ? 1'h0 : dirty_1_56; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5835 = 7'h39 == index[6:0] ? 1'h0 : dirty_1_57; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5836 = 7'h3a == index[6:0] ? 1'h0 : dirty_1_58; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5837 = 7'h3b == index[6:0] ? 1'h0 : dirty_1_59; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5838 = 7'h3c == index[6:0] ? 1'h0 : dirty_1_60; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5839 = 7'h3d == index[6:0] ? 1'h0 : dirty_1_61; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5840 = 7'h3e == index[6:0] ? 1'h0 : dirty_1_62; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5841 = 7'h3f == index[6:0] ? 1'h0 : dirty_1_63; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5842 = 7'h40 == index[6:0] ? 1'h0 : dirty_1_64; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5843 = 7'h41 == index[6:0] ? 1'h0 : dirty_1_65; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5844 = 7'h42 == index[6:0] ? 1'h0 : dirty_1_66; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5845 = 7'h43 == index[6:0] ? 1'h0 : dirty_1_67; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5846 = 7'h44 == index[6:0] ? 1'h0 : dirty_1_68; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5847 = 7'h45 == index[6:0] ? 1'h0 : dirty_1_69; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5848 = 7'h46 == index[6:0] ? 1'h0 : dirty_1_70; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5849 = 7'h47 == index[6:0] ? 1'h0 : dirty_1_71; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5850 = 7'h48 == index[6:0] ? 1'h0 : dirty_1_72; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5851 = 7'h49 == index[6:0] ? 1'h0 : dirty_1_73; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5852 = 7'h4a == index[6:0] ? 1'h0 : dirty_1_74; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5853 = 7'h4b == index[6:0] ? 1'h0 : dirty_1_75; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5854 = 7'h4c == index[6:0] ? 1'h0 : dirty_1_76; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5855 = 7'h4d == index[6:0] ? 1'h0 : dirty_1_77; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5856 = 7'h4e == index[6:0] ? 1'h0 : dirty_1_78; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5857 = 7'h4f == index[6:0] ? 1'h0 : dirty_1_79; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5858 = 7'h50 == index[6:0] ? 1'h0 : dirty_1_80; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5859 = 7'h51 == index[6:0] ? 1'h0 : dirty_1_81; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5860 = 7'h52 == index[6:0] ? 1'h0 : dirty_1_82; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5861 = 7'h53 == index[6:0] ? 1'h0 : dirty_1_83; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5862 = 7'h54 == index[6:0] ? 1'h0 : dirty_1_84; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5863 = 7'h55 == index[6:0] ? 1'h0 : dirty_1_85; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5864 = 7'h56 == index[6:0] ? 1'h0 : dirty_1_86; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5865 = 7'h57 == index[6:0] ? 1'h0 : dirty_1_87; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5866 = 7'h58 == index[6:0] ? 1'h0 : dirty_1_88; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5867 = 7'h59 == index[6:0] ? 1'h0 : dirty_1_89; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5868 = 7'h5a == index[6:0] ? 1'h0 : dirty_1_90; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5869 = 7'h5b == index[6:0] ? 1'h0 : dirty_1_91; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5870 = 7'h5c == index[6:0] ? 1'h0 : dirty_1_92; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5871 = 7'h5d == index[6:0] ? 1'h0 : dirty_1_93; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5872 = 7'h5e == index[6:0] ? 1'h0 : dirty_1_94; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5873 = 7'h5f == index[6:0] ? 1'h0 : dirty_1_95; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5874 = 7'h60 == index[6:0] ? 1'h0 : dirty_1_96; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5875 = 7'h61 == index[6:0] ? 1'h0 : dirty_1_97; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5876 = 7'h62 == index[6:0] ? 1'h0 : dirty_1_98; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5877 = 7'h63 == index[6:0] ? 1'h0 : dirty_1_99; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5878 = 7'h64 == index[6:0] ? 1'h0 : dirty_1_100; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5879 = 7'h65 == index[6:0] ? 1'h0 : dirty_1_101; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5880 = 7'h66 == index[6:0] ? 1'h0 : dirty_1_102; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5881 = 7'h67 == index[6:0] ? 1'h0 : dirty_1_103; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5882 = 7'h68 == index[6:0] ? 1'h0 : dirty_1_104; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5883 = 7'h69 == index[6:0] ? 1'h0 : dirty_1_105; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5884 = 7'h6a == index[6:0] ? 1'h0 : dirty_1_106; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5885 = 7'h6b == index[6:0] ? 1'h0 : dirty_1_107; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5886 = 7'h6c == index[6:0] ? 1'h0 : dirty_1_108; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5887 = 7'h6d == index[6:0] ? 1'h0 : dirty_1_109; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5888 = 7'h6e == index[6:0] ? 1'h0 : dirty_1_110; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5889 = 7'h6f == index[6:0] ? 1'h0 : dirty_1_111; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5890 = 7'h70 == index[6:0] ? 1'h0 : dirty_1_112; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5891 = 7'h71 == index[6:0] ? 1'h0 : dirty_1_113; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5892 = 7'h72 == index[6:0] ? 1'h0 : dirty_1_114; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5893 = 7'h73 == index[6:0] ? 1'h0 : dirty_1_115; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5894 = 7'h74 == index[6:0] ? 1'h0 : dirty_1_116; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5895 = 7'h75 == index[6:0] ? 1'h0 : dirty_1_117; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5896 = 7'h76 == index[6:0] ? 1'h0 : dirty_1_118; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5897 = 7'h77 == index[6:0] ? 1'h0 : dirty_1_119; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5898 = 7'h78 == index[6:0] ? 1'h0 : dirty_1_120; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5899 = 7'h79 == index[6:0] ? 1'h0 : dirty_1_121; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5900 = 7'h7a == index[6:0] ? 1'h0 : dirty_1_122; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5901 = 7'h7b == index[6:0] ? 1'h0 : dirty_1_123; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5902 = 7'h7c == index[6:0] ? 1'h0 : dirty_1_124; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5903 = 7'h7d == index[6:0] ? 1'h0 : dirty_1_125; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5904 = 7'h7e == index[6:0] ? 1'h0 : dirty_1_126; // @[d_cache.scala 171:{40,40} 25:26]
  wire  _GEN_5905 = 7'h7f == index[6:0] ? 1'h0 : dirty_1_127; // @[d_cache.scala 171:{40,40} 25:26]
  wire [63:0] _GEN_6418 = _GEN_1030 ? _GEN_5393 : write_back_data; // @[d_cache.scala 166:47 167:41 29:34]
  wire [41:0] _GEN_6419 = _GEN_1030 ? _write_back_addr_T_7 : {{10'd0}, write_back_addr}; // @[d_cache.scala 166:47 168:41 30:34]
  wire [63:0] _GEN_6420 = _GEN_1030 ? _GEN_2958 : _GEN_2958; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6421 = _GEN_1030 ? _GEN_2959 : _GEN_2959; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6422 = _GEN_1030 ? _GEN_2960 : _GEN_2960; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6423 = _GEN_1030 ? _GEN_2961 : _GEN_2961; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6424 = _GEN_1030 ? _GEN_2962 : _GEN_2962; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6425 = _GEN_1030 ? _GEN_2963 : _GEN_2963; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6426 = _GEN_1030 ? _GEN_2964 : _GEN_2964; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6427 = _GEN_1030 ? _GEN_2965 : _GEN_2965; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6428 = _GEN_1030 ? _GEN_2966 : _GEN_2966; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6429 = _GEN_1030 ? _GEN_2967 : _GEN_2967; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6430 = _GEN_1030 ? _GEN_2968 : _GEN_2968; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6431 = _GEN_1030 ? _GEN_2969 : _GEN_2969; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6432 = _GEN_1030 ? _GEN_2970 : _GEN_2970; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6433 = _GEN_1030 ? _GEN_2971 : _GEN_2971; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6434 = _GEN_1030 ? _GEN_2972 : _GEN_2972; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6435 = _GEN_1030 ? _GEN_2973 : _GEN_2973; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6436 = _GEN_1030 ? _GEN_2974 : _GEN_2974; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6437 = _GEN_1030 ? _GEN_2975 : _GEN_2975; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6438 = _GEN_1030 ? _GEN_2976 : _GEN_2976; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6439 = _GEN_1030 ? _GEN_2977 : _GEN_2977; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6440 = _GEN_1030 ? _GEN_2978 : _GEN_2978; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6441 = _GEN_1030 ? _GEN_2979 : _GEN_2979; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6442 = _GEN_1030 ? _GEN_2980 : _GEN_2980; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6443 = _GEN_1030 ? _GEN_2981 : _GEN_2981; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6444 = _GEN_1030 ? _GEN_2982 : _GEN_2982; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6445 = _GEN_1030 ? _GEN_2983 : _GEN_2983; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6446 = _GEN_1030 ? _GEN_2984 : _GEN_2984; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6447 = _GEN_1030 ? _GEN_2985 : _GEN_2985; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6448 = _GEN_1030 ? _GEN_2986 : _GEN_2986; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6449 = _GEN_1030 ? _GEN_2987 : _GEN_2987; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6450 = _GEN_1030 ? _GEN_2988 : _GEN_2988; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6451 = _GEN_1030 ? _GEN_2989 : _GEN_2989; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6452 = _GEN_1030 ? _GEN_2990 : _GEN_2990; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6453 = _GEN_1030 ? _GEN_2991 : _GEN_2991; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6454 = _GEN_1030 ? _GEN_2992 : _GEN_2992; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6455 = _GEN_1030 ? _GEN_2993 : _GEN_2993; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6456 = _GEN_1030 ? _GEN_2994 : _GEN_2994; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6457 = _GEN_1030 ? _GEN_2995 : _GEN_2995; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6458 = _GEN_1030 ? _GEN_2996 : _GEN_2996; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6459 = _GEN_1030 ? _GEN_2997 : _GEN_2997; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6460 = _GEN_1030 ? _GEN_2998 : _GEN_2998; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6461 = _GEN_1030 ? _GEN_2999 : _GEN_2999; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6462 = _GEN_1030 ? _GEN_3000 : _GEN_3000; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6463 = _GEN_1030 ? _GEN_3001 : _GEN_3001; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6464 = _GEN_1030 ? _GEN_3002 : _GEN_3002; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6465 = _GEN_1030 ? _GEN_3003 : _GEN_3003; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6466 = _GEN_1030 ? _GEN_3004 : _GEN_3004; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6467 = _GEN_1030 ? _GEN_3005 : _GEN_3005; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6468 = _GEN_1030 ? _GEN_3006 : _GEN_3006; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6469 = _GEN_1030 ? _GEN_3007 : _GEN_3007; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6470 = _GEN_1030 ? _GEN_3008 : _GEN_3008; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6471 = _GEN_1030 ? _GEN_3009 : _GEN_3009; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6472 = _GEN_1030 ? _GEN_3010 : _GEN_3010; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6473 = _GEN_1030 ? _GEN_3011 : _GEN_3011; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6474 = _GEN_1030 ? _GEN_3012 : _GEN_3012; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6475 = _GEN_1030 ? _GEN_3013 : _GEN_3013; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6476 = _GEN_1030 ? _GEN_3014 : _GEN_3014; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6477 = _GEN_1030 ? _GEN_3015 : _GEN_3015; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6478 = _GEN_1030 ? _GEN_3016 : _GEN_3016; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6479 = _GEN_1030 ? _GEN_3017 : _GEN_3017; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6480 = _GEN_1030 ? _GEN_3018 : _GEN_3018; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6481 = _GEN_1030 ? _GEN_3019 : _GEN_3019; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6482 = _GEN_1030 ? _GEN_3020 : _GEN_3020; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6483 = _GEN_1030 ? _GEN_3021 : _GEN_3021; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6484 = _GEN_1030 ? _GEN_3022 : _GEN_3022; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6485 = _GEN_1030 ? _GEN_3023 : _GEN_3023; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6486 = _GEN_1030 ? _GEN_3024 : _GEN_3024; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6487 = _GEN_1030 ? _GEN_3025 : _GEN_3025; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6488 = _GEN_1030 ? _GEN_3026 : _GEN_3026; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6489 = _GEN_1030 ? _GEN_3027 : _GEN_3027; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6490 = _GEN_1030 ? _GEN_3028 : _GEN_3028; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6491 = _GEN_1030 ? _GEN_3029 : _GEN_3029; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6492 = _GEN_1030 ? _GEN_3030 : _GEN_3030; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6493 = _GEN_1030 ? _GEN_3031 : _GEN_3031; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6494 = _GEN_1030 ? _GEN_3032 : _GEN_3032; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6495 = _GEN_1030 ? _GEN_3033 : _GEN_3033; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6496 = _GEN_1030 ? _GEN_3034 : _GEN_3034; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6497 = _GEN_1030 ? _GEN_3035 : _GEN_3035; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6498 = _GEN_1030 ? _GEN_3036 : _GEN_3036; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6499 = _GEN_1030 ? _GEN_3037 : _GEN_3037; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6500 = _GEN_1030 ? _GEN_3038 : _GEN_3038; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6501 = _GEN_1030 ? _GEN_3039 : _GEN_3039; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6502 = _GEN_1030 ? _GEN_3040 : _GEN_3040; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6503 = _GEN_1030 ? _GEN_3041 : _GEN_3041; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6504 = _GEN_1030 ? _GEN_3042 : _GEN_3042; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6505 = _GEN_1030 ? _GEN_3043 : _GEN_3043; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6506 = _GEN_1030 ? _GEN_3044 : _GEN_3044; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6507 = _GEN_1030 ? _GEN_3045 : _GEN_3045; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6508 = _GEN_1030 ? _GEN_3046 : _GEN_3046; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6509 = _GEN_1030 ? _GEN_3047 : _GEN_3047; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6510 = _GEN_1030 ? _GEN_3048 : _GEN_3048; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6511 = _GEN_1030 ? _GEN_3049 : _GEN_3049; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6512 = _GEN_1030 ? _GEN_3050 : _GEN_3050; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6513 = _GEN_1030 ? _GEN_3051 : _GEN_3051; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6514 = _GEN_1030 ? _GEN_3052 : _GEN_3052; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6515 = _GEN_1030 ? _GEN_3053 : _GEN_3053; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6516 = _GEN_1030 ? _GEN_3054 : _GEN_3054; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6517 = _GEN_1030 ? _GEN_3055 : _GEN_3055; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6518 = _GEN_1030 ? _GEN_3056 : _GEN_3056; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6519 = _GEN_1030 ? _GEN_3057 : _GEN_3057; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6520 = _GEN_1030 ? _GEN_3058 : _GEN_3058; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6521 = _GEN_1030 ? _GEN_3059 : _GEN_3059; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6522 = _GEN_1030 ? _GEN_3060 : _GEN_3060; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6523 = _GEN_1030 ? _GEN_3061 : _GEN_3061; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6524 = _GEN_1030 ? _GEN_3062 : _GEN_3062; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6525 = _GEN_1030 ? _GEN_3063 : _GEN_3063; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6526 = _GEN_1030 ? _GEN_3064 : _GEN_3064; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6527 = _GEN_1030 ? _GEN_3065 : _GEN_3065; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6528 = _GEN_1030 ? _GEN_3066 : _GEN_3066; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6529 = _GEN_1030 ? _GEN_3067 : _GEN_3067; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6530 = _GEN_1030 ? _GEN_3068 : _GEN_3068; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6531 = _GEN_1030 ? _GEN_3069 : _GEN_3069; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6532 = _GEN_1030 ? _GEN_3070 : _GEN_3070; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6533 = _GEN_1030 ? _GEN_3071 : _GEN_3071; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6534 = _GEN_1030 ? _GEN_3072 : _GEN_3072; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6535 = _GEN_1030 ? _GEN_3073 : _GEN_3073; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6536 = _GEN_1030 ? _GEN_3074 : _GEN_3074; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6537 = _GEN_1030 ? _GEN_3075 : _GEN_3075; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6538 = _GEN_1030 ? _GEN_3076 : _GEN_3076; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6539 = _GEN_1030 ? _GEN_3077 : _GEN_3077; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6540 = _GEN_1030 ? _GEN_3078 : _GEN_3078; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6541 = _GEN_1030 ? _GEN_3079 : _GEN_3079; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6542 = _GEN_1030 ? _GEN_3080 : _GEN_3080; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6543 = _GEN_1030 ? _GEN_3081 : _GEN_3081; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6544 = _GEN_1030 ? _GEN_3082 : _GEN_3082; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6545 = _GEN_1030 ? _GEN_3083 : _GEN_3083; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6546 = _GEN_1030 ? _GEN_3084 : _GEN_3084; // @[d_cache.scala 166:47]
  wire [63:0] _GEN_6547 = _GEN_1030 ? _GEN_3085 : _GEN_3085; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6548 = _GEN_1030 ? _GEN_3086 : _GEN_3086; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6549 = _GEN_1030 ? _GEN_3087 : _GEN_3087; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6550 = _GEN_1030 ? _GEN_3088 : _GEN_3088; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6551 = _GEN_1030 ? _GEN_3089 : _GEN_3089; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6552 = _GEN_1030 ? _GEN_3090 : _GEN_3090; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6553 = _GEN_1030 ? _GEN_3091 : _GEN_3091; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6554 = _GEN_1030 ? _GEN_3092 : _GEN_3092; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6555 = _GEN_1030 ? _GEN_3093 : _GEN_3093; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6556 = _GEN_1030 ? _GEN_3094 : _GEN_3094; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6557 = _GEN_1030 ? _GEN_3095 : _GEN_3095; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6558 = _GEN_1030 ? _GEN_3096 : _GEN_3096; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6559 = _GEN_1030 ? _GEN_3097 : _GEN_3097; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6560 = _GEN_1030 ? _GEN_3098 : _GEN_3098; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6561 = _GEN_1030 ? _GEN_3099 : _GEN_3099; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6562 = _GEN_1030 ? _GEN_3100 : _GEN_3100; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6563 = _GEN_1030 ? _GEN_3101 : _GEN_3101; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6564 = _GEN_1030 ? _GEN_3102 : _GEN_3102; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6565 = _GEN_1030 ? _GEN_3103 : _GEN_3103; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6566 = _GEN_1030 ? _GEN_3104 : _GEN_3104; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6567 = _GEN_1030 ? _GEN_3105 : _GEN_3105; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6568 = _GEN_1030 ? _GEN_3106 : _GEN_3106; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6569 = _GEN_1030 ? _GEN_3107 : _GEN_3107; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6570 = _GEN_1030 ? _GEN_3108 : _GEN_3108; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6571 = _GEN_1030 ? _GEN_3109 : _GEN_3109; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6572 = _GEN_1030 ? _GEN_3110 : _GEN_3110; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6573 = _GEN_1030 ? _GEN_3111 : _GEN_3111; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6574 = _GEN_1030 ? _GEN_3112 : _GEN_3112; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6575 = _GEN_1030 ? _GEN_3113 : _GEN_3113; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6576 = _GEN_1030 ? _GEN_3114 : _GEN_3114; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6577 = _GEN_1030 ? _GEN_3115 : _GEN_3115; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6578 = _GEN_1030 ? _GEN_3116 : _GEN_3116; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6579 = _GEN_1030 ? _GEN_3117 : _GEN_3117; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6580 = _GEN_1030 ? _GEN_3118 : _GEN_3118; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6581 = _GEN_1030 ? _GEN_3119 : _GEN_3119; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6582 = _GEN_1030 ? _GEN_3120 : _GEN_3120; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6583 = _GEN_1030 ? _GEN_3121 : _GEN_3121; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6584 = _GEN_1030 ? _GEN_3122 : _GEN_3122; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6585 = _GEN_1030 ? _GEN_3123 : _GEN_3123; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6586 = _GEN_1030 ? _GEN_3124 : _GEN_3124; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6587 = _GEN_1030 ? _GEN_3125 : _GEN_3125; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6588 = _GEN_1030 ? _GEN_3126 : _GEN_3126; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6589 = _GEN_1030 ? _GEN_3127 : _GEN_3127; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6590 = _GEN_1030 ? _GEN_3128 : _GEN_3128; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6591 = _GEN_1030 ? _GEN_3129 : _GEN_3129; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6592 = _GEN_1030 ? _GEN_3130 : _GEN_3130; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6593 = _GEN_1030 ? _GEN_3131 : _GEN_3131; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6594 = _GEN_1030 ? _GEN_3132 : _GEN_3132; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6595 = _GEN_1030 ? _GEN_3133 : _GEN_3133; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6596 = _GEN_1030 ? _GEN_3134 : _GEN_3134; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6597 = _GEN_1030 ? _GEN_3135 : _GEN_3135; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6598 = _GEN_1030 ? _GEN_3136 : _GEN_3136; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6599 = _GEN_1030 ? _GEN_3137 : _GEN_3137; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6600 = _GEN_1030 ? _GEN_3138 : _GEN_3138; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6601 = _GEN_1030 ? _GEN_3139 : _GEN_3139; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6602 = _GEN_1030 ? _GEN_3140 : _GEN_3140; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6603 = _GEN_1030 ? _GEN_3141 : _GEN_3141; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6604 = _GEN_1030 ? _GEN_3142 : _GEN_3142; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6605 = _GEN_1030 ? _GEN_3143 : _GEN_3143; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6606 = _GEN_1030 ? _GEN_3144 : _GEN_3144; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6607 = _GEN_1030 ? _GEN_3145 : _GEN_3145; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6608 = _GEN_1030 ? _GEN_3146 : _GEN_3146; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6609 = _GEN_1030 ? _GEN_3147 : _GEN_3147; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6610 = _GEN_1030 ? _GEN_3148 : _GEN_3148; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6611 = _GEN_1030 ? _GEN_3149 : _GEN_3149; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6612 = _GEN_1030 ? _GEN_3150 : _GEN_3150; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6613 = _GEN_1030 ? _GEN_3151 : _GEN_3151; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6614 = _GEN_1030 ? _GEN_3152 : _GEN_3152; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6615 = _GEN_1030 ? _GEN_3153 : _GEN_3153; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6616 = _GEN_1030 ? _GEN_3154 : _GEN_3154; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6617 = _GEN_1030 ? _GEN_3155 : _GEN_3155; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6618 = _GEN_1030 ? _GEN_3156 : _GEN_3156; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6619 = _GEN_1030 ? _GEN_3157 : _GEN_3157; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6620 = _GEN_1030 ? _GEN_3158 : _GEN_3158; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6621 = _GEN_1030 ? _GEN_3159 : _GEN_3159; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6622 = _GEN_1030 ? _GEN_3160 : _GEN_3160; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6623 = _GEN_1030 ? _GEN_3161 : _GEN_3161; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6624 = _GEN_1030 ? _GEN_3162 : _GEN_3162; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6625 = _GEN_1030 ? _GEN_3163 : _GEN_3163; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6626 = _GEN_1030 ? _GEN_3164 : _GEN_3164; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6627 = _GEN_1030 ? _GEN_3165 : _GEN_3165; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6628 = _GEN_1030 ? _GEN_3166 : _GEN_3166; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6629 = _GEN_1030 ? _GEN_3167 : _GEN_3167; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6630 = _GEN_1030 ? _GEN_3168 : _GEN_3168; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6631 = _GEN_1030 ? _GEN_3169 : _GEN_3169; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6632 = _GEN_1030 ? _GEN_3170 : _GEN_3170; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6633 = _GEN_1030 ? _GEN_3171 : _GEN_3171; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6634 = _GEN_1030 ? _GEN_3172 : _GEN_3172; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6635 = _GEN_1030 ? _GEN_3173 : _GEN_3173; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6636 = _GEN_1030 ? _GEN_3174 : _GEN_3174; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6637 = _GEN_1030 ? _GEN_3175 : _GEN_3175; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6638 = _GEN_1030 ? _GEN_3176 : _GEN_3176; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6639 = _GEN_1030 ? _GEN_3177 : _GEN_3177; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6640 = _GEN_1030 ? _GEN_3178 : _GEN_3178; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6641 = _GEN_1030 ? _GEN_3179 : _GEN_3179; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6642 = _GEN_1030 ? _GEN_3180 : _GEN_3180; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6643 = _GEN_1030 ? _GEN_3181 : _GEN_3181; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6644 = _GEN_1030 ? _GEN_3182 : _GEN_3182; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6645 = _GEN_1030 ? _GEN_3183 : _GEN_3183; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6646 = _GEN_1030 ? _GEN_3184 : _GEN_3184; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6647 = _GEN_1030 ? _GEN_3185 : _GEN_3185; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6648 = _GEN_1030 ? _GEN_3186 : _GEN_3186; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6649 = _GEN_1030 ? _GEN_3187 : _GEN_3187; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6650 = _GEN_1030 ? _GEN_3188 : _GEN_3188; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6651 = _GEN_1030 ? _GEN_3189 : _GEN_3189; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6652 = _GEN_1030 ? _GEN_3190 : _GEN_3190; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6653 = _GEN_1030 ? _GEN_3191 : _GEN_3191; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6654 = _GEN_1030 ? _GEN_3192 : _GEN_3192; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6655 = _GEN_1030 ? _GEN_3193 : _GEN_3193; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6656 = _GEN_1030 ? _GEN_3194 : _GEN_3194; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6657 = _GEN_1030 ? _GEN_3195 : _GEN_3195; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6658 = _GEN_1030 ? _GEN_3196 : _GEN_3196; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6659 = _GEN_1030 ? _GEN_3197 : _GEN_3197; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6660 = _GEN_1030 ? _GEN_3198 : _GEN_3198; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6661 = _GEN_1030 ? _GEN_3199 : _GEN_3199; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6662 = _GEN_1030 ? _GEN_3200 : _GEN_3200; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6663 = _GEN_1030 ? _GEN_3201 : _GEN_3201; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6664 = _GEN_1030 ? _GEN_3202 : _GEN_3202; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6665 = _GEN_1030 ? _GEN_3203 : _GEN_3203; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6666 = _GEN_1030 ? _GEN_3204 : _GEN_3204; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6667 = _GEN_1030 ? _GEN_3205 : _GEN_3205; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6668 = _GEN_1030 ? _GEN_3206 : _GEN_3206; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6669 = _GEN_1030 ? _GEN_3207 : _GEN_3207; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6670 = _GEN_1030 ? _GEN_3208 : _GEN_3208; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6671 = _GEN_1030 ? _GEN_3209 : _GEN_3209; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6672 = _GEN_1030 ? _GEN_3210 : _GEN_3210; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6673 = _GEN_1030 ? _GEN_3211 : _GEN_3211; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6674 = _GEN_1030 ? _GEN_3212 : _GEN_3212; // @[d_cache.scala 166:47]
  wire [31:0] _GEN_6675 = _GEN_1030 ? _GEN_3213 : _GEN_3213; // @[d_cache.scala 166:47]
  wire  _GEN_6676 = _GEN_1030 ? _GEN_5778 : dirty_1_0; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6677 = _GEN_1030 ? _GEN_5779 : dirty_1_1; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6678 = _GEN_1030 ? _GEN_5780 : dirty_1_2; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6679 = _GEN_1030 ? _GEN_5781 : dirty_1_3; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6680 = _GEN_1030 ? _GEN_5782 : dirty_1_4; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6681 = _GEN_1030 ? _GEN_5783 : dirty_1_5; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6682 = _GEN_1030 ? _GEN_5784 : dirty_1_6; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6683 = _GEN_1030 ? _GEN_5785 : dirty_1_7; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6684 = _GEN_1030 ? _GEN_5786 : dirty_1_8; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6685 = _GEN_1030 ? _GEN_5787 : dirty_1_9; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6686 = _GEN_1030 ? _GEN_5788 : dirty_1_10; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6687 = _GEN_1030 ? _GEN_5789 : dirty_1_11; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6688 = _GEN_1030 ? _GEN_5790 : dirty_1_12; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6689 = _GEN_1030 ? _GEN_5791 : dirty_1_13; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6690 = _GEN_1030 ? _GEN_5792 : dirty_1_14; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6691 = _GEN_1030 ? _GEN_5793 : dirty_1_15; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6692 = _GEN_1030 ? _GEN_5794 : dirty_1_16; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6693 = _GEN_1030 ? _GEN_5795 : dirty_1_17; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6694 = _GEN_1030 ? _GEN_5796 : dirty_1_18; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6695 = _GEN_1030 ? _GEN_5797 : dirty_1_19; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6696 = _GEN_1030 ? _GEN_5798 : dirty_1_20; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6697 = _GEN_1030 ? _GEN_5799 : dirty_1_21; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6698 = _GEN_1030 ? _GEN_5800 : dirty_1_22; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6699 = _GEN_1030 ? _GEN_5801 : dirty_1_23; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6700 = _GEN_1030 ? _GEN_5802 : dirty_1_24; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6701 = _GEN_1030 ? _GEN_5803 : dirty_1_25; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6702 = _GEN_1030 ? _GEN_5804 : dirty_1_26; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6703 = _GEN_1030 ? _GEN_5805 : dirty_1_27; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6704 = _GEN_1030 ? _GEN_5806 : dirty_1_28; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6705 = _GEN_1030 ? _GEN_5807 : dirty_1_29; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6706 = _GEN_1030 ? _GEN_5808 : dirty_1_30; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6707 = _GEN_1030 ? _GEN_5809 : dirty_1_31; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6708 = _GEN_1030 ? _GEN_5810 : dirty_1_32; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6709 = _GEN_1030 ? _GEN_5811 : dirty_1_33; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6710 = _GEN_1030 ? _GEN_5812 : dirty_1_34; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6711 = _GEN_1030 ? _GEN_5813 : dirty_1_35; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6712 = _GEN_1030 ? _GEN_5814 : dirty_1_36; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6713 = _GEN_1030 ? _GEN_5815 : dirty_1_37; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6714 = _GEN_1030 ? _GEN_5816 : dirty_1_38; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6715 = _GEN_1030 ? _GEN_5817 : dirty_1_39; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6716 = _GEN_1030 ? _GEN_5818 : dirty_1_40; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6717 = _GEN_1030 ? _GEN_5819 : dirty_1_41; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6718 = _GEN_1030 ? _GEN_5820 : dirty_1_42; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6719 = _GEN_1030 ? _GEN_5821 : dirty_1_43; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6720 = _GEN_1030 ? _GEN_5822 : dirty_1_44; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6721 = _GEN_1030 ? _GEN_5823 : dirty_1_45; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6722 = _GEN_1030 ? _GEN_5824 : dirty_1_46; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6723 = _GEN_1030 ? _GEN_5825 : dirty_1_47; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6724 = _GEN_1030 ? _GEN_5826 : dirty_1_48; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6725 = _GEN_1030 ? _GEN_5827 : dirty_1_49; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6726 = _GEN_1030 ? _GEN_5828 : dirty_1_50; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6727 = _GEN_1030 ? _GEN_5829 : dirty_1_51; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6728 = _GEN_1030 ? _GEN_5830 : dirty_1_52; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6729 = _GEN_1030 ? _GEN_5831 : dirty_1_53; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6730 = _GEN_1030 ? _GEN_5832 : dirty_1_54; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6731 = _GEN_1030 ? _GEN_5833 : dirty_1_55; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6732 = _GEN_1030 ? _GEN_5834 : dirty_1_56; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6733 = _GEN_1030 ? _GEN_5835 : dirty_1_57; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6734 = _GEN_1030 ? _GEN_5836 : dirty_1_58; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6735 = _GEN_1030 ? _GEN_5837 : dirty_1_59; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6736 = _GEN_1030 ? _GEN_5838 : dirty_1_60; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6737 = _GEN_1030 ? _GEN_5839 : dirty_1_61; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6738 = _GEN_1030 ? _GEN_5840 : dirty_1_62; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6739 = _GEN_1030 ? _GEN_5841 : dirty_1_63; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6740 = _GEN_1030 ? _GEN_5842 : dirty_1_64; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6741 = _GEN_1030 ? _GEN_5843 : dirty_1_65; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6742 = _GEN_1030 ? _GEN_5844 : dirty_1_66; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6743 = _GEN_1030 ? _GEN_5845 : dirty_1_67; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6744 = _GEN_1030 ? _GEN_5846 : dirty_1_68; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6745 = _GEN_1030 ? _GEN_5847 : dirty_1_69; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6746 = _GEN_1030 ? _GEN_5848 : dirty_1_70; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6747 = _GEN_1030 ? _GEN_5849 : dirty_1_71; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6748 = _GEN_1030 ? _GEN_5850 : dirty_1_72; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6749 = _GEN_1030 ? _GEN_5851 : dirty_1_73; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6750 = _GEN_1030 ? _GEN_5852 : dirty_1_74; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6751 = _GEN_1030 ? _GEN_5853 : dirty_1_75; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6752 = _GEN_1030 ? _GEN_5854 : dirty_1_76; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6753 = _GEN_1030 ? _GEN_5855 : dirty_1_77; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6754 = _GEN_1030 ? _GEN_5856 : dirty_1_78; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6755 = _GEN_1030 ? _GEN_5857 : dirty_1_79; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6756 = _GEN_1030 ? _GEN_5858 : dirty_1_80; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6757 = _GEN_1030 ? _GEN_5859 : dirty_1_81; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6758 = _GEN_1030 ? _GEN_5860 : dirty_1_82; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6759 = _GEN_1030 ? _GEN_5861 : dirty_1_83; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6760 = _GEN_1030 ? _GEN_5862 : dirty_1_84; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6761 = _GEN_1030 ? _GEN_5863 : dirty_1_85; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6762 = _GEN_1030 ? _GEN_5864 : dirty_1_86; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6763 = _GEN_1030 ? _GEN_5865 : dirty_1_87; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6764 = _GEN_1030 ? _GEN_5866 : dirty_1_88; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6765 = _GEN_1030 ? _GEN_5867 : dirty_1_89; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6766 = _GEN_1030 ? _GEN_5868 : dirty_1_90; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6767 = _GEN_1030 ? _GEN_5869 : dirty_1_91; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6768 = _GEN_1030 ? _GEN_5870 : dirty_1_92; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6769 = _GEN_1030 ? _GEN_5871 : dirty_1_93; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6770 = _GEN_1030 ? _GEN_5872 : dirty_1_94; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6771 = _GEN_1030 ? _GEN_5873 : dirty_1_95; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6772 = _GEN_1030 ? _GEN_5874 : dirty_1_96; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6773 = _GEN_1030 ? _GEN_5875 : dirty_1_97; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6774 = _GEN_1030 ? _GEN_5876 : dirty_1_98; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6775 = _GEN_1030 ? _GEN_5877 : dirty_1_99; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6776 = _GEN_1030 ? _GEN_5878 : dirty_1_100; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6777 = _GEN_1030 ? _GEN_5879 : dirty_1_101; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6778 = _GEN_1030 ? _GEN_5880 : dirty_1_102; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6779 = _GEN_1030 ? _GEN_5881 : dirty_1_103; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6780 = _GEN_1030 ? _GEN_5882 : dirty_1_104; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6781 = _GEN_1030 ? _GEN_5883 : dirty_1_105; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6782 = _GEN_1030 ? _GEN_5884 : dirty_1_106; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6783 = _GEN_1030 ? _GEN_5885 : dirty_1_107; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6784 = _GEN_1030 ? _GEN_5886 : dirty_1_108; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6785 = _GEN_1030 ? _GEN_5887 : dirty_1_109; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6786 = _GEN_1030 ? _GEN_5888 : dirty_1_110; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6787 = _GEN_1030 ? _GEN_5889 : dirty_1_111; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6788 = _GEN_1030 ? _GEN_5890 : dirty_1_112; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6789 = _GEN_1030 ? _GEN_5891 : dirty_1_113; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6790 = _GEN_1030 ? _GEN_5892 : dirty_1_114; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6791 = _GEN_1030 ? _GEN_5893 : dirty_1_115; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6792 = _GEN_1030 ? _GEN_5894 : dirty_1_116; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6793 = _GEN_1030 ? _GEN_5895 : dirty_1_117; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6794 = _GEN_1030 ? _GEN_5896 : dirty_1_118; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6795 = _GEN_1030 ? _GEN_5897 : dirty_1_119; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6796 = _GEN_1030 ? _GEN_5898 : dirty_1_120; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6797 = _GEN_1030 ? _GEN_5899 : dirty_1_121; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6798 = _GEN_1030 ? _GEN_5900 : dirty_1_122; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6799 = _GEN_1030 ? _GEN_5901 : dirty_1_123; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6800 = _GEN_1030 ? _GEN_5902 : dirty_1_124; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6801 = _GEN_1030 ? _GEN_5903 : dirty_1_125; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6802 = _GEN_1030 ? _GEN_5904 : dirty_1_126; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6803 = _GEN_1030 ? _GEN_5905 : dirty_1_127; // @[d_cache.scala 166:47 25:26]
  wire  _GEN_6804 = _GEN_1030 ? _GEN_3214 : _GEN_3214; // @[d_cache.scala 166:47]
  wire  _GEN_6805 = _GEN_1030 ? _GEN_3215 : _GEN_3215; // @[d_cache.scala 166:47]
  wire  _GEN_6806 = _GEN_1030 ? _GEN_3216 : _GEN_3216; // @[d_cache.scala 166:47]
  wire  _GEN_6807 = _GEN_1030 ? _GEN_3217 : _GEN_3217; // @[d_cache.scala 166:47]
  wire  _GEN_6808 = _GEN_1030 ? _GEN_3218 : _GEN_3218; // @[d_cache.scala 166:47]
  wire  _GEN_6809 = _GEN_1030 ? _GEN_3219 : _GEN_3219; // @[d_cache.scala 166:47]
  wire  _GEN_6810 = _GEN_1030 ? _GEN_3220 : _GEN_3220; // @[d_cache.scala 166:47]
  wire  _GEN_6811 = _GEN_1030 ? _GEN_3221 : _GEN_3221; // @[d_cache.scala 166:47]
  wire  _GEN_6812 = _GEN_1030 ? _GEN_3222 : _GEN_3222; // @[d_cache.scala 166:47]
  wire  _GEN_6813 = _GEN_1030 ? _GEN_3223 : _GEN_3223; // @[d_cache.scala 166:47]
  wire  _GEN_6814 = _GEN_1030 ? _GEN_3224 : _GEN_3224; // @[d_cache.scala 166:47]
  wire  _GEN_6815 = _GEN_1030 ? _GEN_3225 : _GEN_3225; // @[d_cache.scala 166:47]
  wire  _GEN_6816 = _GEN_1030 ? _GEN_3226 : _GEN_3226; // @[d_cache.scala 166:47]
  wire  _GEN_6817 = _GEN_1030 ? _GEN_3227 : _GEN_3227; // @[d_cache.scala 166:47]
  wire  _GEN_6818 = _GEN_1030 ? _GEN_3228 : _GEN_3228; // @[d_cache.scala 166:47]
  wire  _GEN_6819 = _GEN_1030 ? _GEN_3229 : _GEN_3229; // @[d_cache.scala 166:47]
  wire  _GEN_6820 = _GEN_1030 ? _GEN_3230 : _GEN_3230; // @[d_cache.scala 166:47]
  wire  _GEN_6821 = _GEN_1030 ? _GEN_3231 : _GEN_3231; // @[d_cache.scala 166:47]
  wire  _GEN_6822 = _GEN_1030 ? _GEN_3232 : _GEN_3232; // @[d_cache.scala 166:47]
  wire  _GEN_6823 = _GEN_1030 ? _GEN_3233 : _GEN_3233; // @[d_cache.scala 166:47]
  wire  _GEN_6824 = _GEN_1030 ? _GEN_3234 : _GEN_3234; // @[d_cache.scala 166:47]
  wire  _GEN_6825 = _GEN_1030 ? _GEN_3235 : _GEN_3235; // @[d_cache.scala 166:47]
  wire  _GEN_6826 = _GEN_1030 ? _GEN_3236 : _GEN_3236; // @[d_cache.scala 166:47]
  wire  _GEN_6827 = _GEN_1030 ? _GEN_3237 : _GEN_3237; // @[d_cache.scala 166:47]
  wire  _GEN_6828 = _GEN_1030 ? _GEN_3238 : _GEN_3238; // @[d_cache.scala 166:47]
  wire  _GEN_6829 = _GEN_1030 ? _GEN_3239 : _GEN_3239; // @[d_cache.scala 166:47]
  wire  _GEN_6830 = _GEN_1030 ? _GEN_3240 : _GEN_3240; // @[d_cache.scala 166:47]
  wire  _GEN_6831 = _GEN_1030 ? _GEN_3241 : _GEN_3241; // @[d_cache.scala 166:47]
  wire  _GEN_6832 = _GEN_1030 ? _GEN_3242 : _GEN_3242; // @[d_cache.scala 166:47]
  wire  _GEN_6833 = _GEN_1030 ? _GEN_3243 : _GEN_3243; // @[d_cache.scala 166:47]
  wire  _GEN_6834 = _GEN_1030 ? _GEN_3244 : _GEN_3244; // @[d_cache.scala 166:47]
  wire  _GEN_6835 = _GEN_1030 ? _GEN_3245 : _GEN_3245; // @[d_cache.scala 166:47]
  wire  _GEN_6836 = _GEN_1030 ? _GEN_3246 : _GEN_3246; // @[d_cache.scala 166:47]
  wire  _GEN_6837 = _GEN_1030 ? _GEN_3247 : _GEN_3247; // @[d_cache.scala 166:47]
  wire  _GEN_6838 = _GEN_1030 ? _GEN_3248 : _GEN_3248; // @[d_cache.scala 166:47]
  wire  _GEN_6839 = _GEN_1030 ? _GEN_3249 : _GEN_3249; // @[d_cache.scala 166:47]
  wire  _GEN_6840 = _GEN_1030 ? _GEN_3250 : _GEN_3250; // @[d_cache.scala 166:47]
  wire  _GEN_6841 = _GEN_1030 ? _GEN_3251 : _GEN_3251; // @[d_cache.scala 166:47]
  wire  _GEN_6842 = _GEN_1030 ? _GEN_3252 : _GEN_3252; // @[d_cache.scala 166:47]
  wire  _GEN_6843 = _GEN_1030 ? _GEN_3253 : _GEN_3253; // @[d_cache.scala 166:47]
  wire  _GEN_6844 = _GEN_1030 ? _GEN_3254 : _GEN_3254; // @[d_cache.scala 166:47]
  wire  _GEN_6845 = _GEN_1030 ? _GEN_3255 : _GEN_3255; // @[d_cache.scala 166:47]
  wire  _GEN_6846 = _GEN_1030 ? _GEN_3256 : _GEN_3256; // @[d_cache.scala 166:47]
  wire  _GEN_6847 = _GEN_1030 ? _GEN_3257 : _GEN_3257; // @[d_cache.scala 166:47]
  wire  _GEN_6848 = _GEN_1030 ? _GEN_3258 : _GEN_3258; // @[d_cache.scala 166:47]
  wire  _GEN_6849 = _GEN_1030 ? _GEN_3259 : _GEN_3259; // @[d_cache.scala 166:47]
  wire  _GEN_6850 = _GEN_1030 ? _GEN_3260 : _GEN_3260; // @[d_cache.scala 166:47]
  wire  _GEN_6851 = _GEN_1030 ? _GEN_3261 : _GEN_3261; // @[d_cache.scala 166:47]
  wire  _GEN_6852 = _GEN_1030 ? _GEN_3262 : _GEN_3262; // @[d_cache.scala 166:47]
  wire  _GEN_6853 = _GEN_1030 ? _GEN_3263 : _GEN_3263; // @[d_cache.scala 166:47]
  wire  _GEN_6854 = _GEN_1030 ? _GEN_3264 : _GEN_3264; // @[d_cache.scala 166:47]
  wire  _GEN_6855 = _GEN_1030 ? _GEN_3265 : _GEN_3265; // @[d_cache.scala 166:47]
  wire  _GEN_6856 = _GEN_1030 ? _GEN_3266 : _GEN_3266; // @[d_cache.scala 166:47]
  wire  _GEN_6857 = _GEN_1030 ? _GEN_3267 : _GEN_3267; // @[d_cache.scala 166:47]
  wire  _GEN_6858 = _GEN_1030 ? _GEN_3268 : _GEN_3268; // @[d_cache.scala 166:47]
  wire  _GEN_6859 = _GEN_1030 ? _GEN_3269 : _GEN_3269; // @[d_cache.scala 166:47]
  wire  _GEN_6860 = _GEN_1030 ? _GEN_3270 : _GEN_3270; // @[d_cache.scala 166:47]
  wire  _GEN_6861 = _GEN_1030 ? _GEN_3271 : _GEN_3271; // @[d_cache.scala 166:47]
  wire  _GEN_6862 = _GEN_1030 ? _GEN_3272 : _GEN_3272; // @[d_cache.scala 166:47]
  wire  _GEN_6863 = _GEN_1030 ? _GEN_3273 : _GEN_3273; // @[d_cache.scala 166:47]
  wire  _GEN_6864 = _GEN_1030 ? _GEN_3274 : _GEN_3274; // @[d_cache.scala 166:47]
  wire  _GEN_6865 = _GEN_1030 ? _GEN_3275 : _GEN_3275; // @[d_cache.scala 166:47]
  wire  _GEN_6866 = _GEN_1030 ? _GEN_3276 : _GEN_3276; // @[d_cache.scala 166:47]
  wire  _GEN_6867 = _GEN_1030 ? _GEN_3277 : _GEN_3277; // @[d_cache.scala 166:47]
  wire  _GEN_6868 = _GEN_1030 ? _GEN_3278 : _GEN_3278; // @[d_cache.scala 166:47]
  wire  _GEN_6869 = _GEN_1030 ? _GEN_3279 : _GEN_3279; // @[d_cache.scala 166:47]
  wire  _GEN_6870 = _GEN_1030 ? _GEN_3280 : _GEN_3280; // @[d_cache.scala 166:47]
  wire  _GEN_6871 = _GEN_1030 ? _GEN_3281 : _GEN_3281; // @[d_cache.scala 166:47]
  wire  _GEN_6872 = _GEN_1030 ? _GEN_3282 : _GEN_3282; // @[d_cache.scala 166:47]
  wire  _GEN_6873 = _GEN_1030 ? _GEN_3283 : _GEN_3283; // @[d_cache.scala 166:47]
  wire  _GEN_6874 = _GEN_1030 ? _GEN_3284 : _GEN_3284; // @[d_cache.scala 166:47]
  wire  _GEN_6875 = _GEN_1030 ? _GEN_3285 : _GEN_3285; // @[d_cache.scala 166:47]
  wire  _GEN_6876 = _GEN_1030 ? _GEN_3286 : _GEN_3286; // @[d_cache.scala 166:47]
  wire  _GEN_6877 = _GEN_1030 ? _GEN_3287 : _GEN_3287; // @[d_cache.scala 166:47]
  wire  _GEN_6878 = _GEN_1030 ? _GEN_3288 : _GEN_3288; // @[d_cache.scala 166:47]
  wire  _GEN_6879 = _GEN_1030 ? _GEN_3289 : _GEN_3289; // @[d_cache.scala 166:47]
  wire  _GEN_6880 = _GEN_1030 ? _GEN_3290 : _GEN_3290; // @[d_cache.scala 166:47]
  wire  _GEN_6881 = _GEN_1030 ? _GEN_3291 : _GEN_3291; // @[d_cache.scala 166:47]
  wire  _GEN_6882 = _GEN_1030 ? _GEN_3292 : _GEN_3292; // @[d_cache.scala 166:47]
  wire  _GEN_6883 = _GEN_1030 ? _GEN_3293 : _GEN_3293; // @[d_cache.scala 166:47]
  wire  _GEN_6884 = _GEN_1030 ? _GEN_3294 : _GEN_3294; // @[d_cache.scala 166:47]
  wire  _GEN_6885 = _GEN_1030 ? _GEN_3295 : _GEN_3295; // @[d_cache.scala 166:47]
  wire  _GEN_6886 = _GEN_1030 ? _GEN_3296 : _GEN_3296; // @[d_cache.scala 166:47]
  wire  _GEN_6887 = _GEN_1030 ? _GEN_3297 : _GEN_3297; // @[d_cache.scala 166:47]
  wire  _GEN_6888 = _GEN_1030 ? _GEN_3298 : _GEN_3298; // @[d_cache.scala 166:47]
  wire  _GEN_6889 = _GEN_1030 ? _GEN_3299 : _GEN_3299; // @[d_cache.scala 166:47]
  wire  _GEN_6890 = _GEN_1030 ? _GEN_3300 : _GEN_3300; // @[d_cache.scala 166:47]
  wire  _GEN_6891 = _GEN_1030 ? _GEN_3301 : _GEN_3301; // @[d_cache.scala 166:47]
  wire  _GEN_6892 = _GEN_1030 ? _GEN_3302 : _GEN_3302; // @[d_cache.scala 166:47]
  wire  _GEN_6893 = _GEN_1030 ? _GEN_3303 : _GEN_3303; // @[d_cache.scala 166:47]
  wire  _GEN_6894 = _GEN_1030 ? _GEN_3304 : _GEN_3304; // @[d_cache.scala 166:47]
  wire  _GEN_6895 = _GEN_1030 ? _GEN_3305 : _GEN_3305; // @[d_cache.scala 166:47]
  wire  _GEN_6896 = _GEN_1030 ? _GEN_3306 : _GEN_3306; // @[d_cache.scala 166:47]
  wire  _GEN_6897 = _GEN_1030 ? _GEN_3307 : _GEN_3307; // @[d_cache.scala 166:47]
  wire  _GEN_6898 = _GEN_1030 ? _GEN_3308 : _GEN_3308; // @[d_cache.scala 166:47]
  wire  _GEN_6899 = _GEN_1030 ? _GEN_3309 : _GEN_3309; // @[d_cache.scala 166:47]
  wire  _GEN_6900 = _GEN_1030 ? _GEN_3310 : _GEN_3310; // @[d_cache.scala 166:47]
  wire  _GEN_6901 = _GEN_1030 ? _GEN_3311 : _GEN_3311; // @[d_cache.scala 166:47]
  wire  _GEN_6902 = _GEN_1030 ? _GEN_3312 : _GEN_3312; // @[d_cache.scala 166:47]
  wire  _GEN_6903 = _GEN_1030 ? _GEN_3313 : _GEN_3313; // @[d_cache.scala 166:47]
  wire  _GEN_6904 = _GEN_1030 ? _GEN_3314 : _GEN_3314; // @[d_cache.scala 166:47]
  wire  _GEN_6905 = _GEN_1030 ? _GEN_3315 : _GEN_3315; // @[d_cache.scala 166:47]
  wire  _GEN_6906 = _GEN_1030 ? _GEN_3316 : _GEN_3316; // @[d_cache.scala 166:47]
  wire  _GEN_6907 = _GEN_1030 ? _GEN_3317 : _GEN_3317; // @[d_cache.scala 166:47]
  wire  _GEN_6908 = _GEN_1030 ? _GEN_3318 : _GEN_3318; // @[d_cache.scala 166:47]
  wire  _GEN_6909 = _GEN_1030 ? _GEN_3319 : _GEN_3319; // @[d_cache.scala 166:47]
  wire  _GEN_6910 = _GEN_1030 ? _GEN_3320 : _GEN_3320; // @[d_cache.scala 166:47]
  wire  _GEN_6911 = _GEN_1030 ? _GEN_3321 : _GEN_3321; // @[d_cache.scala 166:47]
  wire  _GEN_6912 = _GEN_1030 ? _GEN_3322 : _GEN_3322; // @[d_cache.scala 166:47]
  wire  _GEN_6913 = _GEN_1030 ? _GEN_3323 : _GEN_3323; // @[d_cache.scala 166:47]
  wire  _GEN_6914 = _GEN_1030 ? _GEN_3324 : _GEN_3324; // @[d_cache.scala 166:47]
  wire  _GEN_6915 = _GEN_1030 ? _GEN_3325 : _GEN_3325; // @[d_cache.scala 166:47]
  wire  _GEN_6916 = _GEN_1030 ? _GEN_3326 : _GEN_3326; // @[d_cache.scala 166:47]
  wire  _GEN_6917 = _GEN_1030 ? _GEN_3327 : _GEN_3327; // @[d_cache.scala 166:47]
  wire  _GEN_6918 = _GEN_1030 ? _GEN_3328 : _GEN_3328; // @[d_cache.scala 166:47]
  wire  _GEN_6919 = _GEN_1030 ? _GEN_3329 : _GEN_3329; // @[d_cache.scala 166:47]
  wire  _GEN_6920 = _GEN_1030 ? _GEN_3330 : _GEN_3330; // @[d_cache.scala 166:47]
  wire  _GEN_6921 = _GEN_1030 ? _GEN_3331 : _GEN_3331; // @[d_cache.scala 166:47]
  wire  _GEN_6922 = _GEN_1030 ? _GEN_3332 : _GEN_3332; // @[d_cache.scala 166:47]
  wire  _GEN_6923 = _GEN_1030 ? _GEN_3333 : _GEN_3333; // @[d_cache.scala 166:47]
  wire  _GEN_6924 = _GEN_1030 ? _GEN_3334 : _GEN_3334; // @[d_cache.scala 166:47]
  wire  _GEN_6925 = _GEN_1030 ? _GEN_3335 : _GEN_3335; // @[d_cache.scala 166:47]
  wire  _GEN_6926 = _GEN_1030 ? _GEN_3336 : _GEN_3336; // @[d_cache.scala 166:47]
  wire  _GEN_6927 = _GEN_1030 ? _GEN_3337 : _GEN_3337; // @[d_cache.scala 166:47]
  wire  _GEN_6928 = _GEN_1030 ? _GEN_3338 : _GEN_3338; // @[d_cache.scala 166:47]
  wire  _GEN_6929 = _GEN_1030 ? _GEN_3339 : _GEN_3339; // @[d_cache.scala 166:47]
  wire  _GEN_6930 = _GEN_1030 ? _GEN_3340 : _GEN_3340; // @[d_cache.scala 166:47]
  wire  _GEN_6931 = _GEN_1030 ? _GEN_3341 : _GEN_3341; // @[d_cache.scala 166:47]
  wire [2:0] _GEN_6932 = _GEN_1030 ? 3'h6 : 3'h7; // @[d_cache.scala 166:47 173:31 176:31]
  wire [63:0] _GEN_6934 = ~quene ? _GEN_4622 : _GEN_6418; // @[d_cache.scala 147:34]
  wire [41:0] _GEN_6935 = ~quene ? _GEN_4623 : _GEN_6419; // @[d_cache.scala 147:34]
  wire [63:0] _GEN_6936 = ~quene ? _GEN_4624 : ram_0_0; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6937 = ~quene ? _GEN_4625 : ram_0_1; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6938 = ~quene ? _GEN_4626 : ram_0_2; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6939 = ~quene ? _GEN_4627 : ram_0_3; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6940 = ~quene ? _GEN_4628 : ram_0_4; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6941 = ~quene ? _GEN_4629 : ram_0_5; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6942 = ~quene ? _GEN_4630 : ram_0_6; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6943 = ~quene ? _GEN_4631 : ram_0_7; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6944 = ~quene ? _GEN_4632 : ram_0_8; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6945 = ~quene ? _GEN_4633 : ram_0_9; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6946 = ~quene ? _GEN_4634 : ram_0_10; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6947 = ~quene ? _GEN_4635 : ram_0_11; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6948 = ~quene ? _GEN_4636 : ram_0_12; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6949 = ~quene ? _GEN_4637 : ram_0_13; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6950 = ~quene ? _GEN_4638 : ram_0_14; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6951 = ~quene ? _GEN_4639 : ram_0_15; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6952 = ~quene ? _GEN_4640 : ram_0_16; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6953 = ~quene ? _GEN_4641 : ram_0_17; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6954 = ~quene ? _GEN_4642 : ram_0_18; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6955 = ~quene ? _GEN_4643 : ram_0_19; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6956 = ~quene ? _GEN_4644 : ram_0_20; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6957 = ~quene ? _GEN_4645 : ram_0_21; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6958 = ~quene ? _GEN_4646 : ram_0_22; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6959 = ~quene ? _GEN_4647 : ram_0_23; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6960 = ~quene ? _GEN_4648 : ram_0_24; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6961 = ~quene ? _GEN_4649 : ram_0_25; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6962 = ~quene ? _GEN_4650 : ram_0_26; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6963 = ~quene ? _GEN_4651 : ram_0_27; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6964 = ~quene ? _GEN_4652 : ram_0_28; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6965 = ~quene ? _GEN_4653 : ram_0_29; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6966 = ~quene ? _GEN_4654 : ram_0_30; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6967 = ~quene ? _GEN_4655 : ram_0_31; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6968 = ~quene ? _GEN_4656 : ram_0_32; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6969 = ~quene ? _GEN_4657 : ram_0_33; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6970 = ~quene ? _GEN_4658 : ram_0_34; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6971 = ~quene ? _GEN_4659 : ram_0_35; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6972 = ~quene ? _GEN_4660 : ram_0_36; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6973 = ~quene ? _GEN_4661 : ram_0_37; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6974 = ~quene ? _GEN_4662 : ram_0_38; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6975 = ~quene ? _GEN_4663 : ram_0_39; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6976 = ~quene ? _GEN_4664 : ram_0_40; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6977 = ~quene ? _GEN_4665 : ram_0_41; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6978 = ~quene ? _GEN_4666 : ram_0_42; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6979 = ~quene ? _GEN_4667 : ram_0_43; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6980 = ~quene ? _GEN_4668 : ram_0_44; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6981 = ~quene ? _GEN_4669 : ram_0_45; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6982 = ~quene ? _GEN_4670 : ram_0_46; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6983 = ~quene ? _GEN_4671 : ram_0_47; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6984 = ~quene ? _GEN_4672 : ram_0_48; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6985 = ~quene ? _GEN_4673 : ram_0_49; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6986 = ~quene ? _GEN_4674 : ram_0_50; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6987 = ~quene ? _GEN_4675 : ram_0_51; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6988 = ~quene ? _GEN_4676 : ram_0_52; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6989 = ~quene ? _GEN_4677 : ram_0_53; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6990 = ~quene ? _GEN_4678 : ram_0_54; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6991 = ~quene ? _GEN_4679 : ram_0_55; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6992 = ~quene ? _GEN_4680 : ram_0_56; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6993 = ~quene ? _GEN_4681 : ram_0_57; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6994 = ~quene ? _GEN_4682 : ram_0_58; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6995 = ~quene ? _GEN_4683 : ram_0_59; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6996 = ~quene ? _GEN_4684 : ram_0_60; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6997 = ~quene ? _GEN_4685 : ram_0_61; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6998 = ~quene ? _GEN_4686 : ram_0_62; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_6999 = ~quene ? _GEN_4687 : ram_0_63; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7000 = ~quene ? _GEN_4688 : ram_0_64; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7001 = ~quene ? _GEN_4689 : ram_0_65; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7002 = ~quene ? _GEN_4690 : ram_0_66; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7003 = ~quene ? _GEN_4691 : ram_0_67; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7004 = ~quene ? _GEN_4692 : ram_0_68; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7005 = ~quene ? _GEN_4693 : ram_0_69; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7006 = ~quene ? _GEN_4694 : ram_0_70; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7007 = ~quene ? _GEN_4695 : ram_0_71; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7008 = ~quene ? _GEN_4696 : ram_0_72; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7009 = ~quene ? _GEN_4697 : ram_0_73; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7010 = ~quene ? _GEN_4698 : ram_0_74; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7011 = ~quene ? _GEN_4699 : ram_0_75; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7012 = ~quene ? _GEN_4700 : ram_0_76; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7013 = ~quene ? _GEN_4701 : ram_0_77; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7014 = ~quene ? _GEN_4702 : ram_0_78; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7015 = ~quene ? _GEN_4703 : ram_0_79; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7016 = ~quene ? _GEN_4704 : ram_0_80; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7017 = ~quene ? _GEN_4705 : ram_0_81; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7018 = ~quene ? _GEN_4706 : ram_0_82; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7019 = ~quene ? _GEN_4707 : ram_0_83; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7020 = ~quene ? _GEN_4708 : ram_0_84; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7021 = ~quene ? _GEN_4709 : ram_0_85; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7022 = ~quene ? _GEN_4710 : ram_0_86; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7023 = ~quene ? _GEN_4711 : ram_0_87; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7024 = ~quene ? _GEN_4712 : ram_0_88; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7025 = ~quene ? _GEN_4713 : ram_0_89; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7026 = ~quene ? _GEN_4714 : ram_0_90; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7027 = ~quene ? _GEN_4715 : ram_0_91; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7028 = ~quene ? _GEN_4716 : ram_0_92; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7029 = ~quene ? _GEN_4717 : ram_0_93; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7030 = ~quene ? _GEN_4718 : ram_0_94; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7031 = ~quene ? _GEN_4719 : ram_0_95; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7032 = ~quene ? _GEN_4720 : ram_0_96; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7033 = ~quene ? _GEN_4721 : ram_0_97; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7034 = ~quene ? _GEN_4722 : ram_0_98; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7035 = ~quene ? _GEN_4723 : ram_0_99; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7036 = ~quene ? _GEN_4724 : ram_0_100; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7037 = ~quene ? _GEN_4725 : ram_0_101; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7038 = ~quene ? _GEN_4726 : ram_0_102; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7039 = ~quene ? _GEN_4727 : ram_0_103; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7040 = ~quene ? _GEN_4728 : ram_0_104; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7041 = ~quene ? _GEN_4729 : ram_0_105; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7042 = ~quene ? _GEN_4730 : ram_0_106; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7043 = ~quene ? _GEN_4731 : ram_0_107; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7044 = ~quene ? _GEN_4732 : ram_0_108; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7045 = ~quene ? _GEN_4733 : ram_0_109; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7046 = ~quene ? _GEN_4734 : ram_0_110; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7047 = ~quene ? _GEN_4735 : ram_0_111; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7048 = ~quene ? _GEN_4736 : ram_0_112; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7049 = ~quene ? _GEN_4737 : ram_0_113; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7050 = ~quene ? _GEN_4738 : ram_0_114; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7051 = ~quene ? _GEN_4739 : ram_0_115; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7052 = ~quene ? _GEN_4740 : ram_0_116; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7053 = ~quene ? _GEN_4741 : ram_0_117; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7054 = ~quene ? _GEN_4742 : ram_0_118; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7055 = ~quene ? _GEN_4743 : ram_0_119; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7056 = ~quene ? _GEN_4744 : ram_0_120; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7057 = ~quene ? _GEN_4745 : ram_0_121; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7058 = ~quene ? _GEN_4746 : ram_0_122; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7059 = ~quene ? _GEN_4747 : ram_0_123; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7060 = ~quene ? _GEN_4748 : ram_0_124; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7061 = ~quene ? _GEN_4749 : ram_0_125; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7062 = ~quene ? _GEN_4750 : ram_0_126; // @[d_cache.scala 147:34 18:24]
  wire [63:0] _GEN_7063 = ~quene ? _GEN_4751 : ram_0_127; // @[d_cache.scala 147:34 18:24]
  wire [31:0] _GEN_7064 = ~quene ? _GEN_4752 : tag_0_0; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7065 = ~quene ? _GEN_4753 : tag_0_1; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7066 = ~quene ? _GEN_4754 : tag_0_2; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7067 = ~quene ? _GEN_4755 : tag_0_3; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7068 = ~quene ? _GEN_4756 : tag_0_4; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7069 = ~quene ? _GEN_4757 : tag_0_5; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7070 = ~quene ? _GEN_4758 : tag_0_6; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7071 = ~quene ? _GEN_4759 : tag_0_7; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7072 = ~quene ? _GEN_4760 : tag_0_8; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7073 = ~quene ? _GEN_4761 : tag_0_9; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7074 = ~quene ? _GEN_4762 : tag_0_10; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7075 = ~quene ? _GEN_4763 : tag_0_11; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7076 = ~quene ? _GEN_4764 : tag_0_12; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7077 = ~quene ? _GEN_4765 : tag_0_13; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7078 = ~quene ? _GEN_4766 : tag_0_14; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7079 = ~quene ? _GEN_4767 : tag_0_15; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7080 = ~quene ? _GEN_4768 : tag_0_16; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7081 = ~quene ? _GEN_4769 : tag_0_17; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7082 = ~quene ? _GEN_4770 : tag_0_18; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7083 = ~quene ? _GEN_4771 : tag_0_19; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7084 = ~quene ? _GEN_4772 : tag_0_20; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7085 = ~quene ? _GEN_4773 : tag_0_21; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7086 = ~quene ? _GEN_4774 : tag_0_22; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7087 = ~quene ? _GEN_4775 : tag_0_23; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7088 = ~quene ? _GEN_4776 : tag_0_24; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7089 = ~quene ? _GEN_4777 : tag_0_25; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7090 = ~quene ? _GEN_4778 : tag_0_26; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7091 = ~quene ? _GEN_4779 : tag_0_27; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7092 = ~quene ? _GEN_4780 : tag_0_28; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7093 = ~quene ? _GEN_4781 : tag_0_29; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7094 = ~quene ? _GEN_4782 : tag_0_30; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7095 = ~quene ? _GEN_4783 : tag_0_31; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7096 = ~quene ? _GEN_4784 : tag_0_32; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7097 = ~quene ? _GEN_4785 : tag_0_33; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7098 = ~quene ? _GEN_4786 : tag_0_34; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7099 = ~quene ? _GEN_4787 : tag_0_35; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7100 = ~quene ? _GEN_4788 : tag_0_36; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7101 = ~quene ? _GEN_4789 : tag_0_37; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7102 = ~quene ? _GEN_4790 : tag_0_38; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7103 = ~quene ? _GEN_4791 : tag_0_39; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7104 = ~quene ? _GEN_4792 : tag_0_40; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7105 = ~quene ? _GEN_4793 : tag_0_41; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7106 = ~quene ? _GEN_4794 : tag_0_42; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7107 = ~quene ? _GEN_4795 : tag_0_43; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7108 = ~quene ? _GEN_4796 : tag_0_44; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7109 = ~quene ? _GEN_4797 : tag_0_45; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7110 = ~quene ? _GEN_4798 : tag_0_46; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7111 = ~quene ? _GEN_4799 : tag_0_47; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7112 = ~quene ? _GEN_4800 : tag_0_48; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7113 = ~quene ? _GEN_4801 : tag_0_49; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7114 = ~quene ? _GEN_4802 : tag_0_50; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7115 = ~quene ? _GEN_4803 : tag_0_51; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7116 = ~quene ? _GEN_4804 : tag_0_52; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7117 = ~quene ? _GEN_4805 : tag_0_53; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7118 = ~quene ? _GEN_4806 : tag_0_54; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7119 = ~quene ? _GEN_4807 : tag_0_55; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7120 = ~quene ? _GEN_4808 : tag_0_56; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7121 = ~quene ? _GEN_4809 : tag_0_57; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7122 = ~quene ? _GEN_4810 : tag_0_58; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7123 = ~quene ? _GEN_4811 : tag_0_59; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7124 = ~quene ? _GEN_4812 : tag_0_60; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7125 = ~quene ? _GEN_4813 : tag_0_61; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7126 = ~quene ? _GEN_4814 : tag_0_62; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7127 = ~quene ? _GEN_4815 : tag_0_63; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7128 = ~quene ? _GEN_4816 : tag_0_64; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7129 = ~quene ? _GEN_4817 : tag_0_65; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7130 = ~quene ? _GEN_4818 : tag_0_66; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7131 = ~quene ? _GEN_4819 : tag_0_67; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7132 = ~quene ? _GEN_4820 : tag_0_68; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7133 = ~quene ? _GEN_4821 : tag_0_69; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7134 = ~quene ? _GEN_4822 : tag_0_70; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7135 = ~quene ? _GEN_4823 : tag_0_71; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7136 = ~quene ? _GEN_4824 : tag_0_72; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7137 = ~quene ? _GEN_4825 : tag_0_73; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7138 = ~quene ? _GEN_4826 : tag_0_74; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7139 = ~quene ? _GEN_4827 : tag_0_75; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7140 = ~quene ? _GEN_4828 : tag_0_76; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7141 = ~quene ? _GEN_4829 : tag_0_77; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7142 = ~quene ? _GEN_4830 : tag_0_78; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7143 = ~quene ? _GEN_4831 : tag_0_79; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7144 = ~quene ? _GEN_4832 : tag_0_80; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7145 = ~quene ? _GEN_4833 : tag_0_81; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7146 = ~quene ? _GEN_4834 : tag_0_82; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7147 = ~quene ? _GEN_4835 : tag_0_83; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7148 = ~quene ? _GEN_4836 : tag_0_84; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7149 = ~quene ? _GEN_4837 : tag_0_85; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7150 = ~quene ? _GEN_4838 : tag_0_86; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7151 = ~quene ? _GEN_4839 : tag_0_87; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7152 = ~quene ? _GEN_4840 : tag_0_88; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7153 = ~quene ? _GEN_4841 : tag_0_89; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7154 = ~quene ? _GEN_4842 : tag_0_90; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7155 = ~quene ? _GEN_4843 : tag_0_91; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7156 = ~quene ? _GEN_4844 : tag_0_92; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7157 = ~quene ? _GEN_4845 : tag_0_93; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7158 = ~quene ? _GEN_4846 : tag_0_94; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7159 = ~quene ? _GEN_4847 : tag_0_95; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7160 = ~quene ? _GEN_4848 : tag_0_96; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7161 = ~quene ? _GEN_4849 : tag_0_97; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7162 = ~quene ? _GEN_4850 : tag_0_98; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7163 = ~quene ? _GEN_4851 : tag_0_99; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7164 = ~quene ? _GEN_4852 : tag_0_100; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7165 = ~quene ? _GEN_4853 : tag_0_101; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7166 = ~quene ? _GEN_4854 : tag_0_102; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7167 = ~quene ? _GEN_4855 : tag_0_103; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7168 = ~quene ? _GEN_4856 : tag_0_104; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7169 = ~quene ? _GEN_4857 : tag_0_105; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7170 = ~quene ? _GEN_4858 : tag_0_106; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7171 = ~quene ? _GEN_4859 : tag_0_107; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7172 = ~quene ? _GEN_4860 : tag_0_108; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7173 = ~quene ? _GEN_4861 : tag_0_109; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7174 = ~quene ? _GEN_4862 : tag_0_110; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7175 = ~quene ? _GEN_4863 : tag_0_111; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7176 = ~quene ? _GEN_4864 : tag_0_112; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7177 = ~quene ? _GEN_4865 : tag_0_113; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7178 = ~quene ? _GEN_4866 : tag_0_114; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7179 = ~quene ? _GEN_4867 : tag_0_115; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7180 = ~quene ? _GEN_4868 : tag_0_116; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7181 = ~quene ? _GEN_4869 : tag_0_117; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7182 = ~quene ? _GEN_4870 : tag_0_118; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7183 = ~quene ? _GEN_4871 : tag_0_119; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7184 = ~quene ? _GEN_4872 : tag_0_120; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7185 = ~quene ? _GEN_4873 : tag_0_121; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7186 = ~quene ? _GEN_4874 : tag_0_122; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7187 = ~quene ? _GEN_4875 : tag_0_123; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7188 = ~quene ? _GEN_4876 : tag_0_124; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7189 = ~quene ? _GEN_4877 : tag_0_125; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7190 = ~quene ? _GEN_4878 : tag_0_126; // @[d_cache.scala 147:34 20:24]
  wire [31:0] _GEN_7191 = ~quene ? _GEN_4879 : tag_0_127; // @[d_cache.scala 147:34 20:24]
  wire  _GEN_7192 = ~quene ? _GEN_4880 : dirty_0_0; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7193 = ~quene ? _GEN_4881 : dirty_0_1; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7194 = ~quene ? _GEN_4882 : dirty_0_2; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7195 = ~quene ? _GEN_4883 : dirty_0_3; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7196 = ~quene ? _GEN_4884 : dirty_0_4; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7197 = ~quene ? _GEN_4885 : dirty_0_5; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7198 = ~quene ? _GEN_4886 : dirty_0_6; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7199 = ~quene ? _GEN_4887 : dirty_0_7; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7200 = ~quene ? _GEN_4888 : dirty_0_8; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7201 = ~quene ? _GEN_4889 : dirty_0_9; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7202 = ~quene ? _GEN_4890 : dirty_0_10; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7203 = ~quene ? _GEN_4891 : dirty_0_11; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7204 = ~quene ? _GEN_4892 : dirty_0_12; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7205 = ~quene ? _GEN_4893 : dirty_0_13; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7206 = ~quene ? _GEN_4894 : dirty_0_14; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7207 = ~quene ? _GEN_4895 : dirty_0_15; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7208 = ~quene ? _GEN_4896 : dirty_0_16; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7209 = ~quene ? _GEN_4897 : dirty_0_17; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7210 = ~quene ? _GEN_4898 : dirty_0_18; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7211 = ~quene ? _GEN_4899 : dirty_0_19; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7212 = ~quene ? _GEN_4900 : dirty_0_20; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7213 = ~quene ? _GEN_4901 : dirty_0_21; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7214 = ~quene ? _GEN_4902 : dirty_0_22; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7215 = ~quene ? _GEN_4903 : dirty_0_23; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7216 = ~quene ? _GEN_4904 : dirty_0_24; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7217 = ~quene ? _GEN_4905 : dirty_0_25; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7218 = ~quene ? _GEN_4906 : dirty_0_26; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7219 = ~quene ? _GEN_4907 : dirty_0_27; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7220 = ~quene ? _GEN_4908 : dirty_0_28; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7221 = ~quene ? _GEN_4909 : dirty_0_29; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7222 = ~quene ? _GEN_4910 : dirty_0_30; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7223 = ~quene ? _GEN_4911 : dirty_0_31; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7224 = ~quene ? _GEN_4912 : dirty_0_32; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7225 = ~quene ? _GEN_4913 : dirty_0_33; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7226 = ~quene ? _GEN_4914 : dirty_0_34; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7227 = ~quene ? _GEN_4915 : dirty_0_35; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7228 = ~quene ? _GEN_4916 : dirty_0_36; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7229 = ~quene ? _GEN_4917 : dirty_0_37; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7230 = ~quene ? _GEN_4918 : dirty_0_38; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7231 = ~quene ? _GEN_4919 : dirty_0_39; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7232 = ~quene ? _GEN_4920 : dirty_0_40; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7233 = ~quene ? _GEN_4921 : dirty_0_41; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7234 = ~quene ? _GEN_4922 : dirty_0_42; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7235 = ~quene ? _GEN_4923 : dirty_0_43; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7236 = ~quene ? _GEN_4924 : dirty_0_44; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7237 = ~quene ? _GEN_4925 : dirty_0_45; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7238 = ~quene ? _GEN_4926 : dirty_0_46; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7239 = ~quene ? _GEN_4927 : dirty_0_47; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7240 = ~quene ? _GEN_4928 : dirty_0_48; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7241 = ~quene ? _GEN_4929 : dirty_0_49; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7242 = ~quene ? _GEN_4930 : dirty_0_50; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7243 = ~quene ? _GEN_4931 : dirty_0_51; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7244 = ~quene ? _GEN_4932 : dirty_0_52; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7245 = ~quene ? _GEN_4933 : dirty_0_53; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7246 = ~quene ? _GEN_4934 : dirty_0_54; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7247 = ~quene ? _GEN_4935 : dirty_0_55; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7248 = ~quene ? _GEN_4936 : dirty_0_56; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7249 = ~quene ? _GEN_4937 : dirty_0_57; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7250 = ~quene ? _GEN_4938 : dirty_0_58; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7251 = ~quene ? _GEN_4939 : dirty_0_59; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7252 = ~quene ? _GEN_4940 : dirty_0_60; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7253 = ~quene ? _GEN_4941 : dirty_0_61; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7254 = ~quene ? _GEN_4942 : dirty_0_62; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7255 = ~quene ? _GEN_4943 : dirty_0_63; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7256 = ~quene ? _GEN_4944 : dirty_0_64; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7257 = ~quene ? _GEN_4945 : dirty_0_65; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7258 = ~quene ? _GEN_4946 : dirty_0_66; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7259 = ~quene ? _GEN_4947 : dirty_0_67; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7260 = ~quene ? _GEN_4948 : dirty_0_68; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7261 = ~quene ? _GEN_4949 : dirty_0_69; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7262 = ~quene ? _GEN_4950 : dirty_0_70; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7263 = ~quene ? _GEN_4951 : dirty_0_71; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7264 = ~quene ? _GEN_4952 : dirty_0_72; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7265 = ~quene ? _GEN_4953 : dirty_0_73; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7266 = ~quene ? _GEN_4954 : dirty_0_74; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7267 = ~quene ? _GEN_4955 : dirty_0_75; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7268 = ~quene ? _GEN_4956 : dirty_0_76; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7269 = ~quene ? _GEN_4957 : dirty_0_77; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7270 = ~quene ? _GEN_4958 : dirty_0_78; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7271 = ~quene ? _GEN_4959 : dirty_0_79; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7272 = ~quene ? _GEN_4960 : dirty_0_80; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7273 = ~quene ? _GEN_4961 : dirty_0_81; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7274 = ~quene ? _GEN_4962 : dirty_0_82; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7275 = ~quene ? _GEN_4963 : dirty_0_83; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7276 = ~quene ? _GEN_4964 : dirty_0_84; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7277 = ~quene ? _GEN_4965 : dirty_0_85; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7278 = ~quene ? _GEN_4966 : dirty_0_86; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7279 = ~quene ? _GEN_4967 : dirty_0_87; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7280 = ~quene ? _GEN_4968 : dirty_0_88; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7281 = ~quene ? _GEN_4969 : dirty_0_89; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7282 = ~quene ? _GEN_4970 : dirty_0_90; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7283 = ~quene ? _GEN_4971 : dirty_0_91; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7284 = ~quene ? _GEN_4972 : dirty_0_92; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7285 = ~quene ? _GEN_4973 : dirty_0_93; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7286 = ~quene ? _GEN_4974 : dirty_0_94; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7287 = ~quene ? _GEN_4975 : dirty_0_95; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7288 = ~quene ? _GEN_4976 : dirty_0_96; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7289 = ~quene ? _GEN_4977 : dirty_0_97; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7290 = ~quene ? _GEN_4978 : dirty_0_98; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7291 = ~quene ? _GEN_4979 : dirty_0_99; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7292 = ~quene ? _GEN_4980 : dirty_0_100; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7293 = ~quene ? _GEN_4981 : dirty_0_101; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7294 = ~quene ? _GEN_4982 : dirty_0_102; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7295 = ~quene ? _GEN_4983 : dirty_0_103; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7296 = ~quene ? _GEN_4984 : dirty_0_104; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7297 = ~quene ? _GEN_4985 : dirty_0_105; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7298 = ~quene ? _GEN_4986 : dirty_0_106; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7299 = ~quene ? _GEN_4987 : dirty_0_107; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7300 = ~quene ? _GEN_4988 : dirty_0_108; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7301 = ~quene ? _GEN_4989 : dirty_0_109; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7302 = ~quene ? _GEN_4990 : dirty_0_110; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7303 = ~quene ? _GEN_4991 : dirty_0_111; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7304 = ~quene ? _GEN_4992 : dirty_0_112; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7305 = ~quene ? _GEN_4993 : dirty_0_113; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7306 = ~quene ? _GEN_4994 : dirty_0_114; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7307 = ~quene ? _GEN_4995 : dirty_0_115; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7308 = ~quene ? _GEN_4996 : dirty_0_116; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7309 = ~quene ? _GEN_4997 : dirty_0_117; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7310 = ~quene ? _GEN_4998 : dirty_0_118; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7311 = ~quene ? _GEN_4999 : dirty_0_119; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7312 = ~quene ? _GEN_5000 : dirty_0_120; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7313 = ~quene ? _GEN_5001 : dirty_0_121; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7314 = ~quene ? _GEN_5002 : dirty_0_122; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7315 = ~quene ? _GEN_5003 : dirty_0_123; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7316 = ~quene ? _GEN_5004 : dirty_0_124; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7317 = ~quene ? _GEN_5005 : dirty_0_125; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7318 = ~quene ? _GEN_5006 : dirty_0_126; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7319 = ~quene ? _GEN_5007 : dirty_0_127; // @[d_cache.scala 147:34 24:26]
  wire  _GEN_7320 = ~quene ? _GEN_5008 : valid_0_0; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7321 = ~quene ? _GEN_5009 : valid_0_1; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7322 = ~quene ? _GEN_5010 : valid_0_2; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7323 = ~quene ? _GEN_5011 : valid_0_3; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7324 = ~quene ? _GEN_5012 : valid_0_4; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7325 = ~quene ? _GEN_5013 : valid_0_5; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7326 = ~quene ? _GEN_5014 : valid_0_6; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7327 = ~quene ? _GEN_5015 : valid_0_7; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7328 = ~quene ? _GEN_5016 : valid_0_8; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7329 = ~quene ? _GEN_5017 : valid_0_9; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7330 = ~quene ? _GEN_5018 : valid_0_10; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7331 = ~quene ? _GEN_5019 : valid_0_11; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7332 = ~quene ? _GEN_5020 : valid_0_12; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7333 = ~quene ? _GEN_5021 : valid_0_13; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7334 = ~quene ? _GEN_5022 : valid_0_14; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7335 = ~quene ? _GEN_5023 : valid_0_15; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7336 = ~quene ? _GEN_5024 : valid_0_16; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7337 = ~quene ? _GEN_5025 : valid_0_17; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7338 = ~quene ? _GEN_5026 : valid_0_18; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7339 = ~quene ? _GEN_5027 : valid_0_19; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7340 = ~quene ? _GEN_5028 : valid_0_20; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7341 = ~quene ? _GEN_5029 : valid_0_21; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7342 = ~quene ? _GEN_5030 : valid_0_22; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7343 = ~quene ? _GEN_5031 : valid_0_23; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7344 = ~quene ? _GEN_5032 : valid_0_24; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7345 = ~quene ? _GEN_5033 : valid_0_25; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7346 = ~quene ? _GEN_5034 : valid_0_26; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7347 = ~quene ? _GEN_5035 : valid_0_27; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7348 = ~quene ? _GEN_5036 : valid_0_28; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7349 = ~quene ? _GEN_5037 : valid_0_29; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7350 = ~quene ? _GEN_5038 : valid_0_30; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7351 = ~quene ? _GEN_5039 : valid_0_31; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7352 = ~quene ? _GEN_5040 : valid_0_32; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7353 = ~quene ? _GEN_5041 : valid_0_33; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7354 = ~quene ? _GEN_5042 : valid_0_34; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7355 = ~quene ? _GEN_5043 : valid_0_35; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7356 = ~quene ? _GEN_5044 : valid_0_36; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7357 = ~quene ? _GEN_5045 : valid_0_37; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7358 = ~quene ? _GEN_5046 : valid_0_38; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7359 = ~quene ? _GEN_5047 : valid_0_39; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7360 = ~quene ? _GEN_5048 : valid_0_40; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7361 = ~quene ? _GEN_5049 : valid_0_41; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7362 = ~quene ? _GEN_5050 : valid_0_42; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7363 = ~quene ? _GEN_5051 : valid_0_43; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7364 = ~quene ? _GEN_5052 : valid_0_44; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7365 = ~quene ? _GEN_5053 : valid_0_45; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7366 = ~quene ? _GEN_5054 : valid_0_46; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7367 = ~quene ? _GEN_5055 : valid_0_47; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7368 = ~quene ? _GEN_5056 : valid_0_48; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7369 = ~quene ? _GEN_5057 : valid_0_49; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7370 = ~quene ? _GEN_5058 : valid_0_50; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7371 = ~quene ? _GEN_5059 : valid_0_51; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7372 = ~quene ? _GEN_5060 : valid_0_52; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7373 = ~quene ? _GEN_5061 : valid_0_53; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7374 = ~quene ? _GEN_5062 : valid_0_54; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7375 = ~quene ? _GEN_5063 : valid_0_55; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7376 = ~quene ? _GEN_5064 : valid_0_56; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7377 = ~quene ? _GEN_5065 : valid_0_57; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7378 = ~quene ? _GEN_5066 : valid_0_58; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7379 = ~quene ? _GEN_5067 : valid_0_59; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7380 = ~quene ? _GEN_5068 : valid_0_60; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7381 = ~quene ? _GEN_5069 : valid_0_61; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7382 = ~quene ? _GEN_5070 : valid_0_62; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7383 = ~quene ? _GEN_5071 : valid_0_63; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7384 = ~quene ? _GEN_5072 : valid_0_64; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7385 = ~quene ? _GEN_5073 : valid_0_65; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7386 = ~quene ? _GEN_5074 : valid_0_66; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7387 = ~quene ? _GEN_5075 : valid_0_67; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7388 = ~quene ? _GEN_5076 : valid_0_68; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7389 = ~quene ? _GEN_5077 : valid_0_69; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7390 = ~quene ? _GEN_5078 : valid_0_70; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7391 = ~quene ? _GEN_5079 : valid_0_71; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7392 = ~quene ? _GEN_5080 : valid_0_72; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7393 = ~quene ? _GEN_5081 : valid_0_73; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7394 = ~quene ? _GEN_5082 : valid_0_74; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7395 = ~quene ? _GEN_5083 : valid_0_75; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7396 = ~quene ? _GEN_5084 : valid_0_76; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7397 = ~quene ? _GEN_5085 : valid_0_77; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7398 = ~quene ? _GEN_5086 : valid_0_78; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7399 = ~quene ? _GEN_5087 : valid_0_79; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7400 = ~quene ? _GEN_5088 : valid_0_80; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7401 = ~quene ? _GEN_5089 : valid_0_81; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7402 = ~quene ? _GEN_5090 : valid_0_82; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7403 = ~quene ? _GEN_5091 : valid_0_83; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7404 = ~quene ? _GEN_5092 : valid_0_84; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7405 = ~quene ? _GEN_5093 : valid_0_85; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7406 = ~quene ? _GEN_5094 : valid_0_86; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7407 = ~quene ? _GEN_5095 : valid_0_87; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7408 = ~quene ? _GEN_5096 : valid_0_88; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7409 = ~quene ? _GEN_5097 : valid_0_89; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7410 = ~quene ? _GEN_5098 : valid_0_90; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7411 = ~quene ? _GEN_5099 : valid_0_91; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7412 = ~quene ? _GEN_5100 : valid_0_92; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7413 = ~quene ? _GEN_5101 : valid_0_93; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7414 = ~quene ? _GEN_5102 : valid_0_94; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7415 = ~quene ? _GEN_5103 : valid_0_95; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7416 = ~quene ? _GEN_5104 : valid_0_96; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7417 = ~quene ? _GEN_5105 : valid_0_97; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7418 = ~quene ? _GEN_5106 : valid_0_98; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7419 = ~quene ? _GEN_5107 : valid_0_99; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7420 = ~quene ? _GEN_5108 : valid_0_100; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7421 = ~quene ? _GEN_5109 : valid_0_101; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7422 = ~quene ? _GEN_5110 : valid_0_102; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7423 = ~quene ? _GEN_5111 : valid_0_103; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7424 = ~quene ? _GEN_5112 : valid_0_104; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7425 = ~quene ? _GEN_5113 : valid_0_105; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7426 = ~quene ? _GEN_5114 : valid_0_106; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7427 = ~quene ? _GEN_5115 : valid_0_107; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7428 = ~quene ? _GEN_5116 : valid_0_108; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7429 = ~quene ? _GEN_5117 : valid_0_109; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7430 = ~quene ? _GEN_5118 : valid_0_110; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7431 = ~quene ? _GEN_5119 : valid_0_111; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7432 = ~quene ? _GEN_5120 : valid_0_112; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7433 = ~quene ? _GEN_5121 : valid_0_113; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7434 = ~quene ? _GEN_5122 : valid_0_114; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7435 = ~quene ? _GEN_5123 : valid_0_115; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7436 = ~quene ? _GEN_5124 : valid_0_116; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7437 = ~quene ? _GEN_5125 : valid_0_117; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7438 = ~quene ? _GEN_5126 : valid_0_118; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7439 = ~quene ? _GEN_5127 : valid_0_119; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7440 = ~quene ? _GEN_5128 : valid_0_120; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7441 = ~quene ? _GEN_5129 : valid_0_121; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7442 = ~quene ? _GEN_5130 : valid_0_122; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7443 = ~quene ? _GEN_5131 : valid_0_123; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7444 = ~quene ? _GEN_5132 : valid_0_124; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7445 = ~quene ? _GEN_5133 : valid_0_125; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7446 = ~quene ? _GEN_5134 : valid_0_126; // @[d_cache.scala 147:34 22:26]
  wire  _GEN_7447 = ~quene ? _GEN_5135 : valid_0_127; // @[d_cache.scala 147:34 22:26]
  wire [2:0] _GEN_7448 = ~quene ? _GEN_5136 : _GEN_6932; // @[d_cache.scala 147:34]
  wire [63:0] _GEN_7450 = ~quene ? ram_1_0 : _GEN_6420; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7451 = ~quene ? ram_1_1 : _GEN_6421; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7452 = ~quene ? ram_1_2 : _GEN_6422; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7453 = ~quene ? ram_1_3 : _GEN_6423; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7454 = ~quene ? ram_1_4 : _GEN_6424; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7455 = ~quene ? ram_1_5 : _GEN_6425; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7456 = ~quene ? ram_1_6 : _GEN_6426; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7457 = ~quene ? ram_1_7 : _GEN_6427; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7458 = ~quene ? ram_1_8 : _GEN_6428; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7459 = ~quene ? ram_1_9 : _GEN_6429; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7460 = ~quene ? ram_1_10 : _GEN_6430; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7461 = ~quene ? ram_1_11 : _GEN_6431; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7462 = ~quene ? ram_1_12 : _GEN_6432; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7463 = ~quene ? ram_1_13 : _GEN_6433; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7464 = ~quene ? ram_1_14 : _GEN_6434; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7465 = ~quene ? ram_1_15 : _GEN_6435; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7466 = ~quene ? ram_1_16 : _GEN_6436; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7467 = ~quene ? ram_1_17 : _GEN_6437; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7468 = ~quene ? ram_1_18 : _GEN_6438; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7469 = ~quene ? ram_1_19 : _GEN_6439; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7470 = ~quene ? ram_1_20 : _GEN_6440; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7471 = ~quene ? ram_1_21 : _GEN_6441; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7472 = ~quene ? ram_1_22 : _GEN_6442; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7473 = ~quene ? ram_1_23 : _GEN_6443; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7474 = ~quene ? ram_1_24 : _GEN_6444; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7475 = ~quene ? ram_1_25 : _GEN_6445; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7476 = ~quene ? ram_1_26 : _GEN_6446; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7477 = ~quene ? ram_1_27 : _GEN_6447; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7478 = ~quene ? ram_1_28 : _GEN_6448; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7479 = ~quene ? ram_1_29 : _GEN_6449; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7480 = ~quene ? ram_1_30 : _GEN_6450; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7481 = ~quene ? ram_1_31 : _GEN_6451; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7482 = ~quene ? ram_1_32 : _GEN_6452; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7483 = ~quene ? ram_1_33 : _GEN_6453; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7484 = ~quene ? ram_1_34 : _GEN_6454; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7485 = ~quene ? ram_1_35 : _GEN_6455; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7486 = ~quene ? ram_1_36 : _GEN_6456; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7487 = ~quene ? ram_1_37 : _GEN_6457; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7488 = ~quene ? ram_1_38 : _GEN_6458; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7489 = ~quene ? ram_1_39 : _GEN_6459; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7490 = ~quene ? ram_1_40 : _GEN_6460; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7491 = ~quene ? ram_1_41 : _GEN_6461; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7492 = ~quene ? ram_1_42 : _GEN_6462; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7493 = ~quene ? ram_1_43 : _GEN_6463; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7494 = ~quene ? ram_1_44 : _GEN_6464; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7495 = ~quene ? ram_1_45 : _GEN_6465; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7496 = ~quene ? ram_1_46 : _GEN_6466; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7497 = ~quene ? ram_1_47 : _GEN_6467; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7498 = ~quene ? ram_1_48 : _GEN_6468; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7499 = ~quene ? ram_1_49 : _GEN_6469; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7500 = ~quene ? ram_1_50 : _GEN_6470; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7501 = ~quene ? ram_1_51 : _GEN_6471; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7502 = ~quene ? ram_1_52 : _GEN_6472; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7503 = ~quene ? ram_1_53 : _GEN_6473; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7504 = ~quene ? ram_1_54 : _GEN_6474; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7505 = ~quene ? ram_1_55 : _GEN_6475; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7506 = ~quene ? ram_1_56 : _GEN_6476; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7507 = ~quene ? ram_1_57 : _GEN_6477; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7508 = ~quene ? ram_1_58 : _GEN_6478; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7509 = ~quene ? ram_1_59 : _GEN_6479; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7510 = ~quene ? ram_1_60 : _GEN_6480; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7511 = ~quene ? ram_1_61 : _GEN_6481; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7512 = ~quene ? ram_1_62 : _GEN_6482; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7513 = ~quene ? ram_1_63 : _GEN_6483; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7514 = ~quene ? ram_1_64 : _GEN_6484; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7515 = ~quene ? ram_1_65 : _GEN_6485; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7516 = ~quene ? ram_1_66 : _GEN_6486; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7517 = ~quene ? ram_1_67 : _GEN_6487; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7518 = ~quene ? ram_1_68 : _GEN_6488; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7519 = ~quene ? ram_1_69 : _GEN_6489; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7520 = ~quene ? ram_1_70 : _GEN_6490; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7521 = ~quene ? ram_1_71 : _GEN_6491; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7522 = ~quene ? ram_1_72 : _GEN_6492; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7523 = ~quene ? ram_1_73 : _GEN_6493; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7524 = ~quene ? ram_1_74 : _GEN_6494; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7525 = ~quene ? ram_1_75 : _GEN_6495; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7526 = ~quene ? ram_1_76 : _GEN_6496; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7527 = ~quene ? ram_1_77 : _GEN_6497; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7528 = ~quene ? ram_1_78 : _GEN_6498; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7529 = ~quene ? ram_1_79 : _GEN_6499; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7530 = ~quene ? ram_1_80 : _GEN_6500; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7531 = ~quene ? ram_1_81 : _GEN_6501; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7532 = ~quene ? ram_1_82 : _GEN_6502; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7533 = ~quene ? ram_1_83 : _GEN_6503; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7534 = ~quene ? ram_1_84 : _GEN_6504; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7535 = ~quene ? ram_1_85 : _GEN_6505; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7536 = ~quene ? ram_1_86 : _GEN_6506; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7537 = ~quene ? ram_1_87 : _GEN_6507; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7538 = ~quene ? ram_1_88 : _GEN_6508; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7539 = ~quene ? ram_1_89 : _GEN_6509; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7540 = ~quene ? ram_1_90 : _GEN_6510; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7541 = ~quene ? ram_1_91 : _GEN_6511; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7542 = ~quene ? ram_1_92 : _GEN_6512; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7543 = ~quene ? ram_1_93 : _GEN_6513; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7544 = ~quene ? ram_1_94 : _GEN_6514; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7545 = ~quene ? ram_1_95 : _GEN_6515; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7546 = ~quene ? ram_1_96 : _GEN_6516; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7547 = ~quene ? ram_1_97 : _GEN_6517; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7548 = ~quene ? ram_1_98 : _GEN_6518; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7549 = ~quene ? ram_1_99 : _GEN_6519; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7550 = ~quene ? ram_1_100 : _GEN_6520; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7551 = ~quene ? ram_1_101 : _GEN_6521; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7552 = ~quene ? ram_1_102 : _GEN_6522; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7553 = ~quene ? ram_1_103 : _GEN_6523; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7554 = ~quene ? ram_1_104 : _GEN_6524; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7555 = ~quene ? ram_1_105 : _GEN_6525; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7556 = ~quene ? ram_1_106 : _GEN_6526; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7557 = ~quene ? ram_1_107 : _GEN_6527; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7558 = ~quene ? ram_1_108 : _GEN_6528; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7559 = ~quene ? ram_1_109 : _GEN_6529; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7560 = ~quene ? ram_1_110 : _GEN_6530; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7561 = ~quene ? ram_1_111 : _GEN_6531; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7562 = ~quene ? ram_1_112 : _GEN_6532; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7563 = ~quene ? ram_1_113 : _GEN_6533; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7564 = ~quene ? ram_1_114 : _GEN_6534; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7565 = ~quene ? ram_1_115 : _GEN_6535; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7566 = ~quene ? ram_1_116 : _GEN_6536; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7567 = ~quene ? ram_1_117 : _GEN_6537; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7568 = ~quene ? ram_1_118 : _GEN_6538; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7569 = ~quene ? ram_1_119 : _GEN_6539; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7570 = ~quene ? ram_1_120 : _GEN_6540; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7571 = ~quene ? ram_1_121 : _GEN_6541; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7572 = ~quene ? ram_1_122 : _GEN_6542; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7573 = ~quene ? ram_1_123 : _GEN_6543; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7574 = ~quene ? ram_1_124 : _GEN_6544; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7575 = ~quene ? ram_1_125 : _GEN_6545; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7576 = ~quene ? ram_1_126 : _GEN_6546; // @[d_cache.scala 147:34 19:24]
  wire [63:0] _GEN_7577 = ~quene ? ram_1_127 : _GEN_6547; // @[d_cache.scala 147:34 19:24]
  wire [31:0] _GEN_7578 = ~quene ? tag_1_0 : _GEN_6548; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7579 = ~quene ? tag_1_1 : _GEN_6549; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7580 = ~quene ? tag_1_2 : _GEN_6550; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7581 = ~quene ? tag_1_3 : _GEN_6551; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7582 = ~quene ? tag_1_4 : _GEN_6552; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7583 = ~quene ? tag_1_5 : _GEN_6553; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7584 = ~quene ? tag_1_6 : _GEN_6554; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7585 = ~quene ? tag_1_7 : _GEN_6555; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7586 = ~quene ? tag_1_8 : _GEN_6556; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7587 = ~quene ? tag_1_9 : _GEN_6557; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7588 = ~quene ? tag_1_10 : _GEN_6558; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7589 = ~quene ? tag_1_11 : _GEN_6559; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7590 = ~quene ? tag_1_12 : _GEN_6560; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7591 = ~quene ? tag_1_13 : _GEN_6561; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7592 = ~quene ? tag_1_14 : _GEN_6562; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7593 = ~quene ? tag_1_15 : _GEN_6563; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7594 = ~quene ? tag_1_16 : _GEN_6564; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7595 = ~quene ? tag_1_17 : _GEN_6565; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7596 = ~quene ? tag_1_18 : _GEN_6566; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7597 = ~quene ? tag_1_19 : _GEN_6567; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7598 = ~quene ? tag_1_20 : _GEN_6568; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7599 = ~quene ? tag_1_21 : _GEN_6569; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7600 = ~quene ? tag_1_22 : _GEN_6570; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7601 = ~quene ? tag_1_23 : _GEN_6571; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7602 = ~quene ? tag_1_24 : _GEN_6572; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7603 = ~quene ? tag_1_25 : _GEN_6573; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7604 = ~quene ? tag_1_26 : _GEN_6574; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7605 = ~quene ? tag_1_27 : _GEN_6575; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7606 = ~quene ? tag_1_28 : _GEN_6576; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7607 = ~quene ? tag_1_29 : _GEN_6577; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7608 = ~quene ? tag_1_30 : _GEN_6578; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7609 = ~quene ? tag_1_31 : _GEN_6579; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7610 = ~quene ? tag_1_32 : _GEN_6580; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7611 = ~quene ? tag_1_33 : _GEN_6581; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7612 = ~quene ? tag_1_34 : _GEN_6582; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7613 = ~quene ? tag_1_35 : _GEN_6583; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7614 = ~quene ? tag_1_36 : _GEN_6584; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7615 = ~quene ? tag_1_37 : _GEN_6585; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7616 = ~quene ? tag_1_38 : _GEN_6586; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7617 = ~quene ? tag_1_39 : _GEN_6587; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7618 = ~quene ? tag_1_40 : _GEN_6588; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7619 = ~quene ? tag_1_41 : _GEN_6589; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7620 = ~quene ? tag_1_42 : _GEN_6590; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7621 = ~quene ? tag_1_43 : _GEN_6591; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7622 = ~quene ? tag_1_44 : _GEN_6592; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7623 = ~quene ? tag_1_45 : _GEN_6593; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7624 = ~quene ? tag_1_46 : _GEN_6594; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7625 = ~quene ? tag_1_47 : _GEN_6595; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7626 = ~quene ? tag_1_48 : _GEN_6596; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7627 = ~quene ? tag_1_49 : _GEN_6597; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7628 = ~quene ? tag_1_50 : _GEN_6598; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7629 = ~quene ? tag_1_51 : _GEN_6599; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7630 = ~quene ? tag_1_52 : _GEN_6600; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7631 = ~quene ? tag_1_53 : _GEN_6601; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7632 = ~quene ? tag_1_54 : _GEN_6602; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7633 = ~quene ? tag_1_55 : _GEN_6603; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7634 = ~quene ? tag_1_56 : _GEN_6604; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7635 = ~quene ? tag_1_57 : _GEN_6605; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7636 = ~quene ? tag_1_58 : _GEN_6606; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7637 = ~quene ? tag_1_59 : _GEN_6607; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7638 = ~quene ? tag_1_60 : _GEN_6608; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7639 = ~quene ? tag_1_61 : _GEN_6609; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7640 = ~quene ? tag_1_62 : _GEN_6610; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7641 = ~quene ? tag_1_63 : _GEN_6611; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7642 = ~quene ? tag_1_64 : _GEN_6612; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7643 = ~quene ? tag_1_65 : _GEN_6613; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7644 = ~quene ? tag_1_66 : _GEN_6614; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7645 = ~quene ? tag_1_67 : _GEN_6615; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7646 = ~quene ? tag_1_68 : _GEN_6616; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7647 = ~quene ? tag_1_69 : _GEN_6617; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7648 = ~quene ? tag_1_70 : _GEN_6618; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7649 = ~quene ? tag_1_71 : _GEN_6619; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7650 = ~quene ? tag_1_72 : _GEN_6620; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7651 = ~quene ? tag_1_73 : _GEN_6621; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7652 = ~quene ? tag_1_74 : _GEN_6622; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7653 = ~quene ? tag_1_75 : _GEN_6623; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7654 = ~quene ? tag_1_76 : _GEN_6624; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7655 = ~quene ? tag_1_77 : _GEN_6625; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7656 = ~quene ? tag_1_78 : _GEN_6626; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7657 = ~quene ? tag_1_79 : _GEN_6627; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7658 = ~quene ? tag_1_80 : _GEN_6628; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7659 = ~quene ? tag_1_81 : _GEN_6629; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7660 = ~quene ? tag_1_82 : _GEN_6630; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7661 = ~quene ? tag_1_83 : _GEN_6631; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7662 = ~quene ? tag_1_84 : _GEN_6632; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7663 = ~quene ? tag_1_85 : _GEN_6633; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7664 = ~quene ? tag_1_86 : _GEN_6634; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7665 = ~quene ? tag_1_87 : _GEN_6635; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7666 = ~quene ? tag_1_88 : _GEN_6636; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7667 = ~quene ? tag_1_89 : _GEN_6637; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7668 = ~quene ? tag_1_90 : _GEN_6638; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7669 = ~quene ? tag_1_91 : _GEN_6639; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7670 = ~quene ? tag_1_92 : _GEN_6640; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7671 = ~quene ? tag_1_93 : _GEN_6641; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7672 = ~quene ? tag_1_94 : _GEN_6642; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7673 = ~quene ? tag_1_95 : _GEN_6643; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7674 = ~quene ? tag_1_96 : _GEN_6644; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7675 = ~quene ? tag_1_97 : _GEN_6645; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7676 = ~quene ? tag_1_98 : _GEN_6646; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7677 = ~quene ? tag_1_99 : _GEN_6647; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7678 = ~quene ? tag_1_100 : _GEN_6648; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7679 = ~quene ? tag_1_101 : _GEN_6649; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7680 = ~quene ? tag_1_102 : _GEN_6650; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7681 = ~quene ? tag_1_103 : _GEN_6651; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7682 = ~quene ? tag_1_104 : _GEN_6652; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7683 = ~quene ? tag_1_105 : _GEN_6653; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7684 = ~quene ? tag_1_106 : _GEN_6654; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7685 = ~quene ? tag_1_107 : _GEN_6655; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7686 = ~quene ? tag_1_108 : _GEN_6656; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7687 = ~quene ? tag_1_109 : _GEN_6657; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7688 = ~quene ? tag_1_110 : _GEN_6658; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7689 = ~quene ? tag_1_111 : _GEN_6659; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7690 = ~quene ? tag_1_112 : _GEN_6660; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7691 = ~quene ? tag_1_113 : _GEN_6661; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7692 = ~quene ? tag_1_114 : _GEN_6662; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7693 = ~quene ? tag_1_115 : _GEN_6663; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7694 = ~quene ? tag_1_116 : _GEN_6664; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7695 = ~quene ? tag_1_117 : _GEN_6665; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7696 = ~quene ? tag_1_118 : _GEN_6666; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7697 = ~quene ? tag_1_119 : _GEN_6667; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7698 = ~quene ? tag_1_120 : _GEN_6668; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7699 = ~quene ? tag_1_121 : _GEN_6669; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7700 = ~quene ? tag_1_122 : _GEN_6670; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7701 = ~quene ? tag_1_123 : _GEN_6671; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7702 = ~quene ? tag_1_124 : _GEN_6672; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7703 = ~quene ? tag_1_125 : _GEN_6673; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7704 = ~quene ? tag_1_126 : _GEN_6674; // @[d_cache.scala 147:34 21:24]
  wire [31:0] _GEN_7705 = ~quene ? tag_1_127 : _GEN_6675; // @[d_cache.scala 147:34 21:24]
  wire  _GEN_7706 = ~quene ? dirty_1_0 : _GEN_6676; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7707 = ~quene ? dirty_1_1 : _GEN_6677; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7708 = ~quene ? dirty_1_2 : _GEN_6678; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7709 = ~quene ? dirty_1_3 : _GEN_6679; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7710 = ~quene ? dirty_1_4 : _GEN_6680; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7711 = ~quene ? dirty_1_5 : _GEN_6681; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7712 = ~quene ? dirty_1_6 : _GEN_6682; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7713 = ~quene ? dirty_1_7 : _GEN_6683; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7714 = ~quene ? dirty_1_8 : _GEN_6684; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7715 = ~quene ? dirty_1_9 : _GEN_6685; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7716 = ~quene ? dirty_1_10 : _GEN_6686; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7717 = ~quene ? dirty_1_11 : _GEN_6687; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7718 = ~quene ? dirty_1_12 : _GEN_6688; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7719 = ~quene ? dirty_1_13 : _GEN_6689; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7720 = ~quene ? dirty_1_14 : _GEN_6690; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7721 = ~quene ? dirty_1_15 : _GEN_6691; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7722 = ~quene ? dirty_1_16 : _GEN_6692; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7723 = ~quene ? dirty_1_17 : _GEN_6693; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7724 = ~quene ? dirty_1_18 : _GEN_6694; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7725 = ~quene ? dirty_1_19 : _GEN_6695; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7726 = ~quene ? dirty_1_20 : _GEN_6696; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7727 = ~quene ? dirty_1_21 : _GEN_6697; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7728 = ~quene ? dirty_1_22 : _GEN_6698; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7729 = ~quene ? dirty_1_23 : _GEN_6699; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7730 = ~quene ? dirty_1_24 : _GEN_6700; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7731 = ~quene ? dirty_1_25 : _GEN_6701; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7732 = ~quene ? dirty_1_26 : _GEN_6702; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7733 = ~quene ? dirty_1_27 : _GEN_6703; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7734 = ~quene ? dirty_1_28 : _GEN_6704; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7735 = ~quene ? dirty_1_29 : _GEN_6705; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7736 = ~quene ? dirty_1_30 : _GEN_6706; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7737 = ~quene ? dirty_1_31 : _GEN_6707; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7738 = ~quene ? dirty_1_32 : _GEN_6708; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7739 = ~quene ? dirty_1_33 : _GEN_6709; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7740 = ~quene ? dirty_1_34 : _GEN_6710; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7741 = ~quene ? dirty_1_35 : _GEN_6711; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7742 = ~quene ? dirty_1_36 : _GEN_6712; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7743 = ~quene ? dirty_1_37 : _GEN_6713; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7744 = ~quene ? dirty_1_38 : _GEN_6714; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7745 = ~quene ? dirty_1_39 : _GEN_6715; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7746 = ~quene ? dirty_1_40 : _GEN_6716; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7747 = ~quene ? dirty_1_41 : _GEN_6717; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7748 = ~quene ? dirty_1_42 : _GEN_6718; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7749 = ~quene ? dirty_1_43 : _GEN_6719; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7750 = ~quene ? dirty_1_44 : _GEN_6720; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7751 = ~quene ? dirty_1_45 : _GEN_6721; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7752 = ~quene ? dirty_1_46 : _GEN_6722; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7753 = ~quene ? dirty_1_47 : _GEN_6723; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7754 = ~quene ? dirty_1_48 : _GEN_6724; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7755 = ~quene ? dirty_1_49 : _GEN_6725; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7756 = ~quene ? dirty_1_50 : _GEN_6726; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7757 = ~quene ? dirty_1_51 : _GEN_6727; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7758 = ~quene ? dirty_1_52 : _GEN_6728; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7759 = ~quene ? dirty_1_53 : _GEN_6729; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7760 = ~quene ? dirty_1_54 : _GEN_6730; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7761 = ~quene ? dirty_1_55 : _GEN_6731; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7762 = ~quene ? dirty_1_56 : _GEN_6732; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7763 = ~quene ? dirty_1_57 : _GEN_6733; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7764 = ~quene ? dirty_1_58 : _GEN_6734; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7765 = ~quene ? dirty_1_59 : _GEN_6735; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7766 = ~quene ? dirty_1_60 : _GEN_6736; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7767 = ~quene ? dirty_1_61 : _GEN_6737; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7768 = ~quene ? dirty_1_62 : _GEN_6738; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7769 = ~quene ? dirty_1_63 : _GEN_6739; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7770 = ~quene ? dirty_1_64 : _GEN_6740; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7771 = ~quene ? dirty_1_65 : _GEN_6741; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7772 = ~quene ? dirty_1_66 : _GEN_6742; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7773 = ~quene ? dirty_1_67 : _GEN_6743; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7774 = ~quene ? dirty_1_68 : _GEN_6744; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7775 = ~quene ? dirty_1_69 : _GEN_6745; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7776 = ~quene ? dirty_1_70 : _GEN_6746; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7777 = ~quene ? dirty_1_71 : _GEN_6747; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7778 = ~quene ? dirty_1_72 : _GEN_6748; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7779 = ~quene ? dirty_1_73 : _GEN_6749; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7780 = ~quene ? dirty_1_74 : _GEN_6750; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7781 = ~quene ? dirty_1_75 : _GEN_6751; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7782 = ~quene ? dirty_1_76 : _GEN_6752; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7783 = ~quene ? dirty_1_77 : _GEN_6753; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7784 = ~quene ? dirty_1_78 : _GEN_6754; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7785 = ~quene ? dirty_1_79 : _GEN_6755; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7786 = ~quene ? dirty_1_80 : _GEN_6756; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7787 = ~quene ? dirty_1_81 : _GEN_6757; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7788 = ~quene ? dirty_1_82 : _GEN_6758; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7789 = ~quene ? dirty_1_83 : _GEN_6759; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7790 = ~quene ? dirty_1_84 : _GEN_6760; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7791 = ~quene ? dirty_1_85 : _GEN_6761; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7792 = ~quene ? dirty_1_86 : _GEN_6762; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7793 = ~quene ? dirty_1_87 : _GEN_6763; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7794 = ~quene ? dirty_1_88 : _GEN_6764; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7795 = ~quene ? dirty_1_89 : _GEN_6765; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7796 = ~quene ? dirty_1_90 : _GEN_6766; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7797 = ~quene ? dirty_1_91 : _GEN_6767; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7798 = ~quene ? dirty_1_92 : _GEN_6768; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7799 = ~quene ? dirty_1_93 : _GEN_6769; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7800 = ~quene ? dirty_1_94 : _GEN_6770; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7801 = ~quene ? dirty_1_95 : _GEN_6771; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7802 = ~quene ? dirty_1_96 : _GEN_6772; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7803 = ~quene ? dirty_1_97 : _GEN_6773; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7804 = ~quene ? dirty_1_98 : _GEN_6774; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7805 = ~quene ? dirty_1_99 : _GEN_6775; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7806 = ~quene ? dirty_1_100 : _GEN_6776; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7807 = ~quene ? dirty_1_101 : _GEN_6777; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7808 = ~quene ? dirty_1_102 : _GEN_6778; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7809 = ~quene ? dirty_1_103 : _GEN_6779; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7810 = ~quene ? dirty_1_104 : _GEN_6780; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7811 = ~quene ? dirty_1_105 : _GEN_6781; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7812 = ~quene ? dirty_1_106 : _GEN_6782; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7813 = ~quene ? dirty_1_107 : _GEN_6783; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7814 = ~quene ? dirty_1_108 : _GEN_6784; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7815 = ~quene ? dirty_1_109 : _GEN_6785; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7816 = ~quene ? dirty_1_110 : _GEN_6786; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7817 = ~quene ? dirty_1_111 : _GEN_6787; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7818 = ~quene ? dirty_1_112 : _GEN_6788; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7819 = ~quene ? dirty_1_113 : _GEN_6789; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7820 = ~quene ? dirty_1_114 : _GEN_6790; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7821 = ~quene ? dirty_1_115 : _GEN_6791; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7822 = ~quene ? dirty_1_116 : _GEN_6792; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7823 = ~quene ? dirty_1_117 : _GEN_6793; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7824 = ~quene ? dirty_1_118 : _GEN_6794; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7825 = ~quene ? dirty_1_119 : _GEN_6795; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7826 = ~quene ? dirty_1_120 : _GEN_6796; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7827 = ~quene ? dirty_1_121 : _GEN_6797; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7828 = ~quene ? dirty_1_122 : _GEN_6798; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7829 = ~quene ? dirty_1_123 : _GEN_6799; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7830 = ~quene ? dirty_1_124 : _GEN_6800; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7831 = ~quene ? dirty_1_125 : _GEN_6801; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7832 = ~quene ? dirty_1_126 : _GEN_6802; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7833 = ~quene ? dirty_1_127 : _GEN_6803; // @[d_cache.scala 147:34 25:26]
  wire  _GEN_7834 = ~quene ? valid_1_0 : _GEN_6804; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7835 = ~quene ? valid_1_1 : _GEN_6805; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7836 = ~quene ? valid_1_2 : _GEN_6806; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7837 = ~quene ? valid_1_3 : _GEN_6807; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7838 = ~quene ? valid_1_4 : _GEN_6808; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7839 = ~quene ? valid_1_5 : _GEN_6809; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7840 = ~quene ? valid_1_6 : _GEN_6810; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7841 = ~quene ? valid_1_7 : _GEN_6811; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7842 = ~quene ? valid_1_8 : _GEN_6812; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7843 = ~quene ? valid_1_9 : _GEN_6813; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7844 = ~quene ? valid_1_10 : _GEN_6814; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7845 = ~quene ? valid_1_11 : _GEN_6815; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7846 = ~quene ? valid_1_12 : _GEN_6816; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7847 = ~quene ? valid_1_13 : _GEN_6817; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7848 = ~quene ? valid_1_14 : _GEN_6818; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7849 = ~quene ? valid_1_15 : _GEN_6819; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7850 = ~quene ? valid_1_16 : _GEN_6820; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7851 = ~quene ? valid_1_17 : _GEN_6821; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7852 = ~quene ? valid_1_18 : _GEN_6822; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7853 = ~quene ? valid_1_19 : _GEN_6823; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7854 = ~quene ? valid_1_20 : _GEN_6824; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7855 = ~quene ? valid_1_21 : _GEN_6825; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7856 = ~quene ? valid_1_22 : _GEN_6826; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7857 = ~quene ? valid_1_23 : _GEN_6827; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7858 = ~quene ? valid_1_24 : _GEN_6828; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7859 = ~quene ? valid_1_25 : _GEN_6829; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7860 = ~quene ? valid_1_26 : _GEN_6830; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7861 = ~quene ? valid_1_27 : _GEN_6831; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7862 = ~quene ? valid_1_28 : _GEN_6832; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7863 = ~quene ? valid_1_29 : _GEN_6833; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7864 = ~quene ? valid_1_30 : _GEN_6834; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7865 = ~quene ? valid_1_31 : _GEN_6835; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7866 = ~quene ? valid_1_32 : _GEN_6836; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7867 = ~quene ? valid_1_33 : _GEN_6837; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7868 = ~quene ? valid_1_34 : _GEN_6838; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7869 = ~quene ? valid_1_35 : _GEN_6839; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7870 = ~quene ? valid_1_36 : _GEN_6840; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7871 = ~quene ? valid_1_37 : _GEN_6841; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7872 = ~quene ? valid_1_38 : _GEN_6842; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7873 = ~quene ? valid_1_39 : _GEN_6843; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7874 = ~quene ? valid_1_40 : _GEN_6844; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7875 = ~quene ? valid_1_41 : _GEN_6845; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7876 = ~quene ? valid_1_42 : _GEN_6846; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7877 = ~quene ? valid_1_43 : _GEN_6847; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7878 = ~quene ? valid_1_44 : _GEN_6848; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7879 = ~quene ? valid_1_45 : _GEN_6849; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7880 = ~quene ? valid_1_46 : _GEN_6850; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7881 = ~quene ? valid_1_47 : _GEN_6851; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7882 = ~quene ? valid_1_48 : _GEN_6852; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7883 = ~quene ? valid_1_49 : _GEN_6853; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7884 = ~quene ? valid_1_50 : _GEN_6854; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7885 = ~quene ? valid_1_51 : _GEN_6855; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7886 = ~quene ? valid_1_52 : _GEN_6856; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7887 = ~quene ? valid_1_53 : _GEN_6857; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7888 = ~quene ? valid_1_54 : _GEN_6858; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7889 = ~quene ? valid_1_55 : _GEN_6859; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7890 = ~quene ? valid_1_56 : _GEN_6860; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7891 = ~quene ? valid_1_57 : _GEN_6861; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7892 = ~quene ? valid_1_58 : _GEN_6862; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7893 = ~quene ? valid_1_59 : _GEN_6863; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7894 = ~quene ? valid_1_60 : _GEN_6864; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7895 = ~quene ? valid_1_61 : _GEN_6865; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7896 = ~quene ? valid_1_62 : _GEN_6866; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7897 = ~quene ? valid_1_63 : _GEN_6867; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7898 = ~quene ? valid_1_64 : _GEN_6868; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7899 = ~quene ? valid_1_65 : _GEN_6869; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7900 = ~quene ? valid_1_66 : _GEN_6870; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7901 = ~quene ? valid_1_67 : _GEN_6871; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7902 = ~quene ? valid_1_68 : _GEN_6872; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7903 = ~quene ? valid_1_69 : _GEN_6873; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7904 = ~quene ? valid_1_70 : _GEN_6874; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7905 = ~quene ? valid_1_71 : _GEN_6875; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7906 = ~quene ? valid_1_72 : _GEN_6876; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7907 = ~quene ? valid_1_73 : _GEN_6877; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7908 = ~quene ? valid_1_74 : _GEN_6878; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7909 = ~quene ? valid_1_75 : _GEN_6879; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7910 = ~quene ? valid_1_76 : _GEN_6880; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7911 = ~quene ? valid_1_77 : _GEN_6881; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7912 = ~quene ? valid_1_78 : _GEN_6882; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7913 = ~quene ? valid_1_79 : _GEN_6883; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7914 = ~quene ? valid_1_80 : _GEN_6884; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7915 = ~quene ? valid_1_81 : _GEN_6885; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7916 = ~quene ? valid_1_82 : _GEN_6886; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7917 = ~quene ? valid_1_83 : _GEN_6887; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7918 = ~quene ? valid_1_84 : _GEN_6888; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7919 = ~quene ? valid_1_85 : _GEN_6889; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7920 = ~quene ? valid_1_86 : _GEN_6890; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7921 = ~quene ? valid_1_87 : _GEN_6891; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7922 = ~quene ? valid_1_88 : _GEN_6892; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7923 = ~quene ? valid_1_89 : _GEN_6893; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7924 = ~quene ? valid_1_90 : _GEN_6894; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7925 = ~quene ? valid_1_91 : _GEN_6895; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7926 = ~quene ? valid_1_92 : _GEN_6896; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7927 = ~quene ? valid_1_93 : _GEN_6897; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7928 = ~quene ? valid_1_94 : _GEN_6898; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7929 = ~quene ? valid_1_95 : _GEN_6899; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7930 = ~quene ? valid_1_96 : _GEN_6900; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7931 = ~quene ? valid_1_97 : _GEN_6901; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7932 = ~quene ? valid_1_98 : _GEN_6902; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7933 = ~quene ? valid_1_99 : _GEN_6903; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7934 = ~quene ? valid_1_100 : _GEN_6904; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7935 = ~quene ? valid_1_101 : _GEN_6905; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7936 = ~quene ? valid_1_102 : _GEN_6906; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7937 = ~quene ? valid_1_103 : _GEN_6907; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7938 = ~quene ? valid_1_104 : _GEN_6908; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7939 = ~quene ? valid_1_105 : _GEN_6909; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7940 = ~quene ? valid_1_106 : _GEN_6910; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7941 = ~quene ? valid_1_107 : _GEN_6911; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7942 = ~quene ? valid_1_108 : _GEN_6912; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7943 = ~quene ? valid_1_109 : _GEN_6913; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7944 = ~quene ? valid_1_110 : _GEN_6914; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7945 = ~quene ? valid_1_111 : _GEN_6915; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7946 = ~quene ? valid_1_112 : _GEN_6916; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7947 = ~quene ? valid_1_113 : _GEN_6917; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7948 = ~quene ? valid_1_114 : _GEN_6918; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7949 = ~quene ? valid_1_115 : _GEN_6919; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7950 = ~quene ? valid_1_116 : _GEN_6920; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7951 = ~quene ? valid_1_117 : _GEN_6921; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7952 = ~quene ? valid_1_118 : _GEN_6922; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7953 = ~quene ? valid_1_119 : _GEN_6923; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7954 = ~quene ? valid_1_120 : _GEN_6924; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7955 = ~quene ? valid_1_121 : _GEN_6925; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7956 = ~quene ? valid_1_122 : _GEN_6926; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7957 = ~quene ? valid_1_123 : _GEN_6927; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7958 = ~quene ? valid_1_124 : _GEN_6928; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7959 = ~quene ? valid_1_125 : _GEN_6929; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7960 = ~quene ? valid_1_126 : _GEN_6930; // @[d_cache.scala 147:34 23:26]
  wire  _GEN_7961 = ~quene ? valid_1_127 : _GEN_6931; // @[d_cache.scala 147:34 23:26]
  wire [2:0] _GEN_7962 = unuse_way == 2'h2 ? 3'h7 : _GEN_7448; // @[d_cache.scala 140:40 141:23]
  wire [63:0] _GEN_7963 = unuse_way == 2'h2 ? _GEN_2958 : _GEN_7450; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7964 = unuse_way == 2'h2 ? _GEN_2959 : _GEN_7451; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7965 = unuse_way == 2'h2 ? _GEN_2960 : _GEN_7452; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7966 = unuse_way == 2'h2 ? _GEN_2961 : _GEN_7453; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7967 = unuse_way == 2'h2 ? _GEN_2962 : _GEN_7454; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7968 = unuse_way == 2'h2 ? _GEN_2963 : _GEN_7455; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7969 = unuse_way == 2'h2 ? _GEN_2964 : _GEN_7456; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7970 = unuse_way == 2'h2 ? _GEN_2965 : _GEN_7457; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7971 = unuse_way == 2'h2 ? _GEN_2966 : _GEN_7458; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7972 = unuse_way == 2'h2 ? _GEN_2967 : _GEN_7459; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7973 = unuse_way == 2'h2 ? _GEN_2968 : _GEN_7460; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7974 = unuse_way == 2'h2 ? _GEN_2969 : _GEN_7461; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7975 = unuse_way == 2'h2 ? _GEN_2970 : _GEN_7462; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7976 = unuse_way == 2'h2 ? _GEN_2971 : _GEN_7463; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7977 = unuse_way == 2'h2 ? _GEN_2972 : _GEN_7464; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7978 = unuse_way == 2'h2 ? _GEN_2973 : _GEN_7465; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7979 = unuse_way == 2'h2 ? _GEN_2974 : _GEN_7466; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7980 = unuse_way == 2'h2 ? _GEN_2975 : _GEN_7467; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7981 = unuse_way == 2'h2 ? _GEN_2976 : _GEN_7468; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7982 = unuse_way == 2'h2 ? _GEN_2977 : _GEN_7469; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7983 = unuse_way == 2'h2 ? _GEN_2978 : _GEN_7470; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7984 = unuse_way == 2'h2 ? _GEN_2979 : _GEN_7471; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7985 = unuse_way == 2'h2 ? _GEN_2980 : _GEN_7472; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7986 = unuse_way == 2'h2 ? _GEN_2981 : _GEN_7473; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7987 = unuse_way == 2'h2 ? _GEN_2982 : _GEN_7474; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7988 = unuse_way == 2'h2 ? _GEN_2983 : _GEN_7475; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7989 = unuse_way == 2'h2 ? _GEN_2984 : _GEN_7476; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7990 = unuse_way == 2'h2 ? _GEN_2985 : _GEN_7477; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7991 = unuse_way == 2'h2 ? _GEN_2986 : _GEN_7478; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7992 = unuse_way == 2'h2 ? _GEN_2987 : _GEN_7479; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7993 = unuse_way == 2'h2 ? _GEN_2988 : _GEN_7480; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7994 = unuse_way == 2'h2 ? _GEN_2989 : _GEN_7481; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7995 = unuse_way == 2'h2 ? _GEN_2990 : _GEN_7482; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7996 = unuse_way == 2'h2 ? _GEN_2991 : _GEN_7483; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7997 = unuse_way == 2'h2 ? _GEN_2992 : _GEN_7484; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7998 = unuse_way == 2'h2 ? _GEN_2993 : _GEN_7485; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_7999 = unuse_way == 2'h2 ? _GEN_2994 : _GEN_7486; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8000 = unuse_way == 2'h2 ? _GEN_2995 : _GEN_7487; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8001 = unuse_way == 2'h2 ? _GEN_2996 : _GEN_7488; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8002 = unuse_way == 2'h2 ? _GEN_2997 : _GEN_7489; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8003 = unuse_way == 2'h2 ? _GEN_2998 : _GEN_7490; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8004 = unuse_way == 2'h2 ? _GEN_2999 : _GEN_7491; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8005 = unuse_way == 2'h2 ? _GEN_3000 : _GEN_7492; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8006 = unuse_way == 2'h2 ? _GEN_3001 : _GEN_7493; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8007 = unuse_way == 2'h2 ? _GEN_3002 : _GEN_7494; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8008 = unuse_way == 2'h2 ? _GEN_3003 : _GEN_7495; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8009 = unuse_way == 2'h2 ? _GEN_3004 : _GEN_7496; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8010 = unuse_way == 2'h2 ? _GEN_3005 : _GEN_7497; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8011 = unuse_way == 2'h2 ? _GEN_3006 : _GEN_7498; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8012 = unuse_way == 2'h2 ? _GEN_3007 : _GEN_7499; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8013 = unuse_way == 2'h2 ? _GEN_3008 : _GEN_7500; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8014 = unuse_way == 2'h2 ? _GEN_3009 : _GEN_7501; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8015 = unuse_way == 2'h2 ? _GEN_3010 : _GEN_7502; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8016 = unuse_way == 2'h2 ? _GEN_3011 : _GEN_7503; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8017 = unuse_way == 2'h2 ? _GEN_3012 : _GEN_7504; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8018 = unuse_way == 2'h2 ? _GEN_3013 : _GEN_7505; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8019 = unuse_way == 2'h2 ? _GEN_3014 : _GEN_7506; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8020 = unuse_way == 2'h2 ? _GEN_3015 : _GEN_7507; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8021 = unuse_way == 2'h2 ? _GEN_3016 : _GEN_7508; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8022 = unuse_way == 2'h2 ? _GEN_3017 : _GEN_7509; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8023 = unuse_way == 2'h2 ? _GEN_3018 : _GEN_7510; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8024 = unuse_way == 2'h2 ? _GEN_3019 : _GEN_7511; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8025 = unuse_way == 2'h2 ? _GEN_3020 : _GEN_7512; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8026 = unuse_way == 2'h2 ? _GEN_3021 : _GEN_7513; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8027 = unuse_way == 2'h2 ? _GEN_3022 : _GEN_7514; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8028 = unuse_way == 2'h2 ? _GEN_3023 : _GEN_7515; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8029 = unuse_way == 2'h2 ? _GEN_3024 : _GEN_7516; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8030 = unuse_way == 2'h2 ? _GEN_3025 : _GEN_7517; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8031 = unuse_way == 2'h2 ? _GEN_3026 : _GEN_7518; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8032 = unuse_way == 2'h2 ? _GEN_3027 : _GEN_7519; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8033 = unuse_way == 2'h2 ? _GEN_3028 : _GEN_7520; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8034 = unuse_way == 2'h2 ? _GEN_3029 : _GEN_7521; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8035 = unuse_way == 2'h2 ? _GEN_3030 : _GEN_7522; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8036 = unuse_way == 2'h2 ? _GEN_3031 : _GEN_7523; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8037 = unuse_way == 2'h2 ? _GEN_3032 : _GEN_7524; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8038 = unuse_way == 2'h2 ? _GEN_3033 : _GEN_7525; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8039 = unuse_way == 2'h2 ? _GEN_3034 : _GEN_7526; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8040 = unuse_way == 2'h2 ? _GEN_3035 : _GEN_7527; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8041 = unuse_way == 2'h2 ? _GEN_3036 : _GEN_7528; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8042 = unuse_way == 2'h2 ? _GEN_3037 : _GEN_7529; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8043 = unuse_way == 2'h2 ? _GEN_3038 : _GEN_7530; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8044 = unuse_way == 2'h2 ? _GEN_3039 : _GEN_7531; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8045 = unuse_way == 2'h2 ? _GEN_3040 : _GEN_7532; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8046 = unuse_way == 2'h2 ? _GEN_3041 : _GEN_7533; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8047 = unuse_way == 2'h2 ? _GEN_3042 : _GEN_7534; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8048 = unuse_way == 2'h2 ? _GEN_3043 : _GEN_7535; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8049 = unuse_way == 2'h2 ? _GEN_3044 : _GEN_7536; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8050 = unuse_way == 2'h2 ? _GEN_3045 : _GEN_7537; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8051 = unuse_way == 2'h2 ? _GEN_3046 : _GEN_7538; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8052 = unuse_way == 2'h2 ? _GEN_3047 : _GEN_7539; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8053 = unuse_way == 2'h2 ? _GEN_3048 : _GEN_7540; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8054 = unuse_way == 2'h2 ? _GEN_3049 : _GEN_7541; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8055 = unuse_way == 2'h2 ? _GEN_3050 : _GEN_7542; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8056 = unuse_way == 2'h2 ? _GEN_3051 : _GEN_7543; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8057 = unuse_way == 2'h2 ? _GEN_3052 : _GEN_7544; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8058 = unuse_way == 2'h2 ? _GEN_3053 : _GEN_7545; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8059 = unuse_way == 2'h2 ? _GEN_3054 : _GEN_7546; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8060 = unuse_way == 2'h2 ? _GEN_3055 : _GEN_7547; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8061 = unuse_way == 2'h2 ? _GEN_3056 : _GEN_7548; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8062 = unuse_way == 2'h2 ? _GEN_3057 : _GEN_7549; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8063 = unuse_way == 2'h2 ? _GEN_3058 : _GEN_7550; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8064 = unuse_way == 2'h2 ? _GEN_3059 : _GEN_7551; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8065 = unuse_way == 2'h2 ? _GEN_3060 : _GEN_7552; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8066 = unuse_way == 2'h2 ? _GEN_3061 : _GEN_7553; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8067 = unuse_way == 2'h2 ? _GEN_3062 : _GEN_7554; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8068 = unuse_way == 2'h2 ? _GEN_3063 : _GEN_7555; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8069 = unuse_way == 2'h2 ? _GEN_3064 : _GEN_7556; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8070 = unuse_way == 2'h2 ? _GEN_3065 : _GEN_7557; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8071 = unuse_way == 2'h2 ? _GEN_3066 : _GEN_7558; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8072 = unuse_way == 2'h2 ? _GEN_3067 : _GEN_7559; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8073 = unuse_way == 2'h2 ? _GEN_3068 : _GEN_7560; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8074 = unuse_way == 2'h2 ? _GEN_3069 : _GEN_7561; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8075 = unuse_way == 2'h2 ? _GEN_3070 : _GEN_7562; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8076 = unuse_way == 2'h2 ? _GEN_3071 : _GEN_7563; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8077 = unuse_way == 2'h2 ? _GEN_3072 : _GEN_7564; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8078 = unuse_way == 2'h2 ? _GEN_3073 : _GEN_7565; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8079 = unuse_way == 2'h2 ? _GEN_3074 : _GEN_7566; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8080 = unuse_way == 2'h2 ? _GEN_3075 : _GEN_7567; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8081 = unuse_way == 2'h2 ? _GEN_3076 : _GEN_7568; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8082 = unuse_way == 2'h2 ? _GEN_3077 : _GEN_7569; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8083 = unuse_way == 2'h2 ? _GEN_3078 : _GEN_7570; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8084 = unuse_way == 2'h2 ? _GEN_3079 : _GEN_7571; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8085 = unuse_way == 2'h2 ? _GEN_3080 : _GEN_7572; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8086 = unuse_way == 2'h2 ? _GEN_3081 : _GEN_7573; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8087 = unuse_way == 2'h2 ? _GEN_3082 : _GEN_7574; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8088 = unuse_way == 2'h2 ? _GEN_3083 : _GEN_7575; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8089 = unuse_way == 2'h2 ? _GEN_3084 : _GEN_7576; // @[d_cache.scala 140:40]
  wire [63:0] _GEN_8090 = unuse_way == 2'h2 ? _GEN_3085 : _GEN_7577; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8091 = unuse_way == 2'h2 ? _GEN_3086 : _GEN_7578; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8092 = unuse_way == 2'h2 ? _GEN_3087 : _GEN_7579; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8093 = unuse_way == 2'h2 ? _GEN_3088 : _GEN_7580; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8094 = unuse_way == 2'h2 ? _GEN_3089 : _GEN_7581; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8095 = unuse_way == 2'h2 ? _GEN_3090 : _GEN_7582; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8096 = unuse_way == 2'h2 ? _GEN_3091 : _GEN_7583; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8097 = unuse_way == 2'h2 ? _GEN_3092 : _GEN_7584; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8098 = unuse_way == 2'h2 ? _GEN_3093 : _GEN_7585; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8099 = unuse_way == 2'h2 ? _GEN_3094 : _GEN_7586; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8100 = unuse_way == 2'h2 ? _GEN_3095 : _GEN_7587; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8101 = unuse_way == 2'h2 ? _GEN_3096 : _GEN_7588; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8102 = unuse_way == 2'h2 ? _GEN_3097 : _GEN_7589; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8103 = unuse_way == 2'h2 ? _GEN_3098 : _GEN_7590; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8104 = unuse_way == 2'h2 ? _GEN_3099 : _GEN_7591; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8105 = unuse_way == 2'h2 ? _GEN_3100 : _GEN_7592; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8106 = unuse_way == 2'h2 ? _GEN_3101 : _GEN_7593; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8107 = unuse_way == 2'h2 ? _GEN_3102 : _GEN_7594; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8108 = unuse_way == 2'h2 ? _GEN_3103 : _GEN_7595; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8109 = unuse_way == 2'h2 ? _GEN_3104 : _GEN_7596; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8110 = unuse_way == 2'h2 ? _GEN_3105 : _GEN_7597; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8111 = unuse_way == 2'h2 ? _GEN_3106 : _GEN_7598; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8112 = unuse_way == 2'h2 ? _GEN_3107 : _GEN_7599; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8113 = unuse_way == 2'h2 ? _GEN_3108 : _GEN_7600; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8114 = unuse_way == 2'h2 ? _GEN_3109 : _GEN_7601; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8115 = unuse_way == 2'h2 ? _GEN_3110 : _GEN_7602; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8116 = unuse_way == 2'h2 ? _GEN_3111 : _GEN_7603; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8117 = unuse_way == 2'h2 ? _GEN_3112 : _GEN_7604; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8118 = unuse_way == 2'h2 ? _GEN_3113 : _GEN_7605; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8119 = unuse_way == 2'h2 ? _GEN_3114 : _GEN_7606; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8120 = unuse_way == 2'h2 ? _GEN_3115 : _GEN_7607; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8121 = unuse_way == 2'h2 ? _GEN_3116 : _GEN_7608; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8122 = unuse_way == 2'h2 ? _GEN_3117 : _GEN_7609; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8123 = unuse_way == 2'h2 ? _GEN_3118 : _GEN_7610; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8124 = unuse_way == 2'h2 ? _GEN_3119 : _GEN_7611; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8125 = unuse_way == 2'h2 ? _GEN_3120 : _GEN_7612; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8126 = unuse_way == 2'h2 ? _GEN_3121 : _GEN_7613; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8127 = unuse_way == 2'h2 ? _GEN_3122 : _GEN_7614; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8128 = unuse_way == 2'h2 ? _GEN_3123 : _GEN_7615; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8129 = unuse_way == 2'h2 ? _GEN_3124 : _GEN_7616; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8130 = unuse_way == 2'h2 ? _GEN_3125 : _GEN_7617; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8131 = unuse_way == 2'h2 ? _GEN_3126 : _GEN_7618; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8132 = unuse_way == 2'h2 ? _GEN_3127 : _GEN_7619; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8133 = unuse_way == 2'h2 ? _GEN_3128 : _GEN_7620; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8134 = unuse_way == 2'h2 ? _GEN_3129 : _GEN_7621; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8135 = unuse_way == 2'h2 ? _GEN_3130 : _GEN_7622; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8136 = unuse_way == 2'h2 ? _GEN_3131 : _GEN_7623; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8137 = unuse_way == 2'h2 ? _GEN_3132 : _GEN_7624; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8138 = unuse_way == 2'h2 ? _GEN_3133 : _GEN_7625; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8139 = unuse_way == 2'h2 ? _GEN_3134 : _GEN_7626; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8140 = unuse_way == 2'h2 ? _GEN_3135 : _GEN_7627; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8141 = unuse_way == 2'h2 ? _GEN_3136 : _GEN_7628; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8142 = unuse_way == 2'h2 ? _GEN_3137 : _GEN_7629; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8143 = unuse_way == 2'h2 ? _GEN_3138 : _GEN_7630; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8144 = unuse_way == 2'h2 ? _GEN_3139 : _GEN_7631; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8145 = unuse_way == 2'h2 ? _GEN_3140 : _GEN_7632; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8146 = unuse_way == 2'h2 ? _GEN_3141 : _GEN_7633; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8147 = unuse_way == 2'h2 ? _GEN_3142 : _GEN_7634; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8148 = unuse_way == 2'h2 ? _GEN_3143 : _GEN_7635; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8149 = unuse_way == 2'h2 ? _GEN_3144 : _GEN_7636; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8150 = unuse_way == 2'h2 ? _GEN_3145 : _GEN_7637; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8151 = unuse_way == 2'h2 ? _GEN_3146 : _GEN_7638; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8152 = unuse_way == 2'h2 ? _GEN_3147 : _GEN_7639; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8153 = unuse_way == 2'h2 ? _GEN_3148 : _GEN_7640; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8154 = unuse_way == 2'h2 ? _GEN_3149 : _GEN_7641; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8155 = unuse_way == 2'h2 ? _GEN_3150 : _GEN_7642; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8156 = unuse_way == 2'h2 ? _GEN_3151 : _GEN_7643; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8157 = unuse_way == 2'h2 ? _GEN_3152 : _GEN_7644; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8158 = unuse_way == 2'h2 ? _GEN_3153 : _GEN_7645; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8159 = unuse_way == 2'h2 ? _GEN_3154 : _GEN_7646; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8160 = unuse_way == 2'h2 ? _GEN_3155 : _GEN_7647; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8161 = unuse_way == 2'h2 ? _GEN_3156 : _GEN_7648; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8162 = unuse_way == 2'h2 ? _GEN_3157 : _GEN_7649; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8163 = unuse_way == 2'h2 ? _GEN_3158 : _GEN_7650; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8164 = unuse_way == 2'h2 ? _GEN_3159 : _GEN_7651; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8165 = unuse_way == 2'h2 ? _GEN_3160 : _GEN_7652; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8166 = unuse_way == 2'h2 ? _GEN_3161 : _GEN_7653; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8167 = unuse_way == 2'h2 ? _GEN_3162 : _GEN_7654; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8168 = unuse_way == 2'h2 ? _GEN_3163 : _GEN_7655; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8169 = unuse_way == 2'h2 ? _GEN_3164 : _GEN_7656; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8170 = unuse_way == 2'h2 ? _GEN_3165 : _GEN_7657; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8171 = unuse_way == 2'h2 ? _GEN_3166 : _GEN_7658; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8172 = unuse_way == 2'h2 ? _GEN_3167 : _GEN_7659; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8173 = unuse_way == 2'h2 ? _GEN_3168 : _GEN_7660; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8174 = unuse_way == 2'h2 ? _GEN_3169 : _GEN_7661; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8175 = unuse_way == 2'h2 ? _GEN_3170 : _GEN_7662; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8176 = unuse_way == 2'h2 ? _GEN_3171 : _GEN_7663; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8177 = unuse_way == 2'h2 ? _GEN_3172 : _GEN_7664; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8178 = unuse_way == 2'h2 ? _GEN_3173 : _GEN_7665; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8179 = unuse_way == 2'h2 ? _GEN_3174 : _GEN_7666; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8180 = unuse_way == 2'h2 ? _GEN_3175 : _GEN_7667; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8181 = unuse_way == 2'h2 ? _GEN_3176 : _GEN_7668; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8182 = unuse_way == 2'h2 ? _GEN_3177 : _GEN_7669; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8183 = unuse_way == 2'h2 ? _GEN_3178 : _GEN_7670; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8184 = unuse_way == 2'h2 ? _GEN_3179 : _GEN_7671; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8185 = unuse_way == 2'h2 ? _GEN_3180 : _GEN_7672; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8186 = unuse_way == 2'h2 ? _GEN_3181 : _GEN_7673; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8187 = unuse_way == 2'h2 ? _GEN_3182 : _GEN_7674; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8188 = unuse_way == 2'h2 ? _GEN_3183 : _GEN_7675; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8189 = unuse_way == 2'h2 ? _GEN_3184 : _GEN_7676; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8190 = unuse_way == 2'h2 ? _GEN_3185 : _GEN_7677; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8191 = unuse_way == 2'h2 ? _GEN_3186 : _GEN_7678; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8192 = unuse_way == 2'h2 ? _GEN_3187 : _GEN_7679; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8193 = unuse_way == 2'h2 ? _GEN_3188 : _GEN_7680; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8194 = unuse_way == 2'h2 ? _GEN_3189 : _GEN_7681; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8195 = unuse_way == 2'h2 ? _GEN_3190 : _GEN_7682; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8196 = unuse_way == 2'h2 ? _GEN_3191 : _GEN_7683; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8197 = unuse_way == 2'h2 ? _GEN_3192 : _GEN_7684; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8198 = unuse_way == 2'h2 ? _GEN_3193 : _GEN_7685; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8199 = unuse_way == 2'h2 ? _GEN_3194 : _GEN_7686; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8200 = unuse_way == 2'h2 ? _GEN_3195 : _GEN_7687; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8201 = unuse_way == 2'h2 ? _GEN_3196 : _GEN_7688; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8202 = unuse_way == 2'h2 ? _GEN_3197 : _GEN_7689; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8203 = unuse_way == 2'h2 ? _GEN_3198 : _GEN_7690; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8204 = unuse_way == 2'h2 ? _GEN_3199 : _GEN_7691; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8205 = unuse_way == 2'h2 ? _GEN_3200 : _GEN_7692; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8206 = unuse_way == 2'h2 ? _GEN_3201 : _GEN_7693; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8207 = unuse_way == 2'h2 ? _GEN_3202 : _GEN_7694; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8208 = unuse_way == 2'h2 ? _GEN_3203 : _GEN_7695; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8209 = unuse_way == 2'h2 ? _GEN_3204 : _GEN_7696; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8210 = unuse_way == 2'h2 ? _GEN_3205 : _GEN_7697; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8211 = unuse_way == 2'h2 ? _GEN_3206 : _GEN_7698; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8212 = unuse_way == 2'h2 ? _GEN_3207 : _GEN_7699; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8213 = unuse_way == 2'h2 ? _GEN_3208 : _GEN_7700; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8214 = unuse_way == 2'h2 ? _GEN_3209 : _GEN_7701; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8215 = unuse_way == 2'h2 ? _GEN_3210 : _GEN_7702; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8216 = unuse_way == 2'h2 ? _GEN_3211 : _GEN_7703; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8217 = unuse_way == 2'h2 ? _GEN_3212 : _GEN_7704; // @[d_cache.scala 140:40]
  wire [31:0] _GEN_8218 = unuse_way == 2'h2 ? _GEN_3213 : _GEN_7705; // @[d_cache.scala 140:40]
  wire  _GEN_8219 = unuse_way == 2'h2 ? _GEN_3214 : _GEN_7834; // @[d_cache.scala 140:40]
  wire  _GEN_8220 = unuse_way == 2'h2 ? _GEN_3215 : _GEN_7835; // @[d_cache.scala 140:40]
  wire  _GEN_8221 = unuse_way == 2'h2 ? _GEN_3216 : _GEN_7836; // @[d_cache.scala 140:40]
  wire  _GEN_8222 = unuse_way == 2'h2 ? _GEN_3217 : _GEN_7837; // @[d_cache.scala 140:40]
  wire  _GEN_8223 = unuse_way == 2'h2 ? _GEN_3218 : _GEN_7838; // @[d_cache.scala 140:40]
  wire  _GEN_8224 = unuse_way == 2'h2 ? _GEN_3219 : _GEN_7839; // @[d_cache.scala 140:40]
  wire  _GEN_8225 = unuse_way == 2'h2 ? _GEN_3220 : _GEN_7840; // @[d_cache.scala 140:40]
  wire  _GEN_8226 = unuse_way == 2'h2 ? _GEN_3221 : _GEN_7841; // @[d_cache.scala 140:40]
  wire  _GEN_8227 = unuse_way == 2'h2 ? _GEN_3222 : _GEN_7842; // @[d_cache.scala 140:40]
  wire  _GEN_8228 = unuse_way == 2'h2 ? _GEN_3223 : _GEN_7843; // @[d_cache.scala 140:40]
  wire  _GEN_8229 = unuse_way == 2'h2 ? _GEN_3224 : _GEN_7844; // @[d_cache.scala 140:40]
  wire  _GEN_8230 = unuse_way == 2'h2 ? _GEN_3225 : _GEN_7845; // @[d_cache.scala 140:40]
  wire  _GEN_8231 = unuse_way == 2'h2 ? _GEN_3226 : _GEN_7846; // @[d_cache.scala 140:40]
  wire  _GEN_8232 = unuse_way == 2'h2 ? _GEN_3227 : _GEN_7847; // @[d_cache.scala 140:40]
  wire  _GEN_8233 = unuse_way == 2'h2 ? _GEN_3228 : _GEN_7848; // @[d_cache.scala 140:40]
  wire  _GEN_8234 = unuse_way == 2'h2 ? _GEN_3229 : _GEN_7849; // @[d_cache.scala 140:40]
  wire  _GEN_8235 = unuse_way == 2'h2 ? _GEN_3230 : _GEN_7850; // @[d_cache.scala 140:40]
  wire  _GEN_8236 = unuse_way == 2'h2 ? _GEN_3231 : _GEN_7851; // @[d_cache.scala 140:40]
  wire  _GEN_8237 = unuse_way == 2'h2 ? _GEN_3232 : _GEN_7852; // @[d_cache.scala 140:40]
  wire  _GEN_8238 = unuse_way == 2'h2 ? _GEN_3233 : _GEN_7853; // @[d_cache.scala 140:40]
  wire  _GEN_8239 = unuse_way == 2'h2 ? _GEN_3234 : _GEN_7854; // @[d_cache.scala 140:40]
  wire  _GEN_8240 = unuse_way == 2'h2 ? _GEN_3235 : _GEN_7855; // @[d_cache.scala 140:40]
  wire  _GEN_8241 = unuse_way == 2'h2 ? _GEN_3236 : _GEN_7856; // @[d_cache.scala 140:40]
  wire  _GEN_8242 = unuse_way == 2'h2 ? _GEN_3237 : _GEN_7857; // @[d_cache.scala 140:40]
  wire  _GEN_8243 = unuse_way == 2'h2 ? _GEN_3238 : _GEN_7858; // @[d_cache.scala 140:40]
  wire  _GEN_8244 = unuse_way == 2'h2 ? _GEN_3239 : _GEN_7859; // @[d_cache.scala 140:40]
  wire  _GEN_8245 = unuse_way == 2'h2 ? _GEN_3240 : _GEN_7860; // @[d_cache.scala 140:40]
  wire  _GEN_8246 = unuse_way == 2'h2 ? _GEN_3241 : _GEN_7861; // @[d_cache.scala 140:40]
  wire  _GEN_8247 = unuse_way == 2'h2 ? _GEN_3242 : _GEN_7862; // @[d_cache.scala 140:40]
  wire  _GEN_8248 = unuse_way == 2'h2 ? _GEN_3243 : _GEN_7863; // @[d_cache.scala 140:40]
  wire  _GEN_8249 = unuse_way == 2'h2 ? _GEN_3244 : _GEN_7864; // @[d_cache.scala 140:40]
  wire  _GEN_8250 = unuse_way == 2'h2 ? _GEN_3245 : _GEN_7865; // @[d_cache.scala 140:40]
  wire  _GEN_8251 = unuse_way == 2'h2 ? _GEN_3246 : _GEN_7866; // @[d_cache.scala 140:40]
  wire  _GEN_8252 = unuse_way == 2'h2 ? _GEN_3247 : _GEN_7867; // @[d_cache.scala 140:40]
  wire  _GEN_8253 = unuse_way == 2'h2 ? _GEN_3248 : _GEN_7868; // @[d_cache.scala 140:40]
  wire  _GEN_8254 = unuse_way == 2'h2 ? _GEN_3249 : _GEN_7869; // @[d_cache.scala 140:40]
  wire  _GEN_8255 = unuse_way == 2'h2 ? _GEN_3250 : _GEN_7870; // @[d_cache.scala 140:40]
  wire  _GEN_8256 = unuse_way == 2'h2 ? _GEN_3251 : _GEN_7871; // @[d_cache.scala 140:40]
  wire  _GEN_8257 = unuse_way == 2'h2 ? _GEN_3252 : _GEN_7872; // @[d_cache.scala 140:40]
  wire  _GEN_8258 = unuse_way == 2'h2 ? _GEN_3253 : _GEN_7873; // @[d_cache.scala 140:40]
  wire  _GEN_8259 = unuse_way == 2'h2 ? _GEN_3254 : _GEN_7874; // @[d_cache.scala 140:40]
  wire  _GEN_8260 = unuse_way == 2'h2 ? _GEN_3255 : _GEN_7875; // @[d_cache.scala 140:40]
  wire  _GEN_8261 = unuse_way == 2'h2 ? _GEN_3256 : _GEN_7876; // @[d_cache.scala 140:40]
  wire  _GEN_8262 = unuse_way == 2'h2 ? _GEN_3257 : _GEN_7877; // @[d_cache.scala 140:40]
  wire  _GEN_8263 = unuse_way == 2'h2 ? _GEN_3258 : _GEN_7878; // @[d_cache.scala 140:40]
  wire  _GEN_8264 = unuse_way == 2'h2 ? _GEN_3259 : _GEN_7879; // @[d_cache.scala 140:40]
  wire  _GEN_8265 = unuse_way == 2'h2 ? _GEN_3260 : _GEN_7880; // @[d_cache.scala 140:40]
  wire  _GEN_8266 = unuse_way == 2'h2 ? _GEN_3261 : _GEN_7881; // @[d_cache.scala 140:40]
  wire  _GEN_8267 = unuse_way == 2'h2 ? _GEN_3262 : _GEN_7882; // @[d_cache.scala 140:40]
  wire  _GEN_8268 = unuse_way == 2'h2 ? _GEN_3263 : _GEN_7883; // @[d_cache.scala 140:40]
  wire  _GEN_8269 = unuse_way == 2'h2 ? _GEN_3264 : _GEN_7884; // @[d_cache.scala 140:40]
  wire  _GEN_8270 = unuse_way == 2'h2 ? _GEN_3265 : _GEN_7885; // @[d_cache.scala 140:40]
  wire  _GEN_8271 = unuse_way == 2'h2 ? _GEN_3266 : _GEN_7886; // @[d_cache.scala 140:40]
  wire  _GEN_8272 = unuse_way == 2'h2 ? _GEN_3267 : _GEN_7887; // @[d_cache.scala 140:40]
  wire  _GEN_8273 = unuse_way == 2'h2 ? _GEN_3268 : _GEN_7888; // @[d_cache.scala 140:40]
  wire  _GEN_8274 = unuse_way == 2'h2 ? _GEN_3269 : _GEN_7889; // @[d_cache.scala 140:40]
  wire  _GEN_8275 = unuse_way == 2'h2 ? _GEN_3270 : _GEN_7890; // @[d_cache.scala 140:40]
  wire  _GEN_8276 = unuse_way == 2'h2 ? _GEN_3271 : _GEN_7891; // @[d_cache.scala 140:40]
  wire  _GEN_8277 = unuse_way == 2'h2 ? _GEN_3272 : _GEN_7892; // @[d_cache.scala 140:40]
  wire  _GEN_8278 = unuse_way == 2'h2 ? _GEN_3273 : _GEN_7893; // @[d_cache.scala 140:40]
  wire  _GEN_8279 = unuse_way == 2'h2 ? _GEN_3274 : _GEN_7894; // @[d_cache.scala 140:40]
  wire  _GEN_8280 = unuse_way == 2'h2 ? _GEN_3275 : _GEN_7895; // @[d_cache.scala 140:40]
  wire  _GEN_8281 = unuse_way == 2'h2 ? _GEN_3276 : _GEN_7896; // @[d_cache.scala 140:40]
  wire  _GEN_8282 = unuse_way == 2'h2 ? _GEN_3277 : _GEN_7897; // @[d_cache.scala 140:40]
  wire  _GEN_8283 = unuse_way == 2'h2 ? _GEN_3278 : _GEN_7898; // @[d_cache.scala 140:40]
  wire  _GEN_8284 = unuse_way == 2'h2 ? _GEN_3279 : _GEN_7899; // @[d_cache.scala 140:40]
  wire  _GEN_8285 = unuse_way == 2'h2 ? _GEN_3280 : _GEN_7900; // @[d_cache.scala 140:40]
  wire  _GEN_8286 = unuse_way == 2'h2 ? _GEN_3281 : _GEN_7901; // @[d_cache.scala 140:40]
  wire  _GEN_8287 = unuse_way == 2'h2 ? _GEN_3282 : _GEN_7902; // @[d_cache.scala 140:40]
  wire  _GEN_8288 = unuse_way == 2'h2 ? _GEN_3283 : _GEN_7903; // @[d_cache.scala 140:40]
  wire  _GEN_8289 = unuse_way == 2'h2 ? _GEN_3284 : _GEN_7904; // @[d_cache.scala 140:40]
  wire  _GEN_8290 = unuse_way == 2'h2 ? _GEN_3285 : _GEN_7905; // @[d_cache.scala 140:40]
  wire  _GEN_8291 = unuse_way == 2'h2 ? _GEN_3286 : _GEN_7906; // @[d_cache.scala 140:40]
  wire  _GEN_8292 = unuse_way == 2'h2 ? _GEN_3287 : _GEN_7907; // @[d_cache.scala 140:40]
  wire  _GEN_8293 = unuse_way == 2'h2 ? _GEN_3288 : _GEN_7908; // @[d_cache.scala 140:40]
  wire  _GEN_8294 = unuse_way == 2'h2 ? _GEN_3289 : _GEN_7909; // @[d_cache.scala 140:40]
  wire  _GEN_8295 = unuse_way == 2'h2 ? _GEN_3290 : _GEN_7910; // @[d_cache.scala 140:40]
  wire  _GEN_8296 = unuse_way == 2'h2 ? _GEN_3291 : _GEN_7911; // @[d_cache.scala 140:40]
  wire  _GEN_8297 = unuse_way == 2'h2 ? _GEN_3292 : _GEN_7912; // @[d_cache.scala 140:40]
  wire  _GEN_8298 = unuse_way == 2'h2 ? _GEN_3293 : _GEN_7913; // @[d_cache.scala 140:40]
  wire  _GEN_8299 = unuse_way == 2'h2 ? _GEN_3294 : _GEN_7914; // @[d_cache.scala 140:40]
  wire  _GEN_8300 = unuse_way == 2'h2 ? _GEN_3295 : _GEN_7915; // @[d_cache.scala 140:40]
  wire  _GEN_8301 = unuse_way == 2'h2 ? _GEN_3296 : _GEN_7916; // @[d_cache.scala 140:40]
  wire  _GEN_8302 = unuse_way == 2'h2 ? _GEN_3297 : _GEN_7917; // @[d_cache.scala 140:40]
  wire  _GEN_8303 = unuse_way == 2'h2 ? _GEN_3298 : _GEN_7918; // @[d_cache.scala 140:40]
  wire  _GEN_8304 = unuse_way == 2'h2 ? _GEN_3299 : _GEN_7919; // @[d_cache.scala 140:40]
  wire  _GEN_8305 = unuse_way == 2'h2 ? _GEN_3300 : _GEN_7920; // @[d_cache.scala 140:40]
  wire  _GEN_8306 = unuse_way == 2'h2 ? _GEN_3301 : _GEN_7921; // @[d_cache.scala 140:40]
  wire  _GEN_8307 = unuse_way == 2'h2 ? _GEN_3302 : _GEN_7922; // @[d_cache.scala 140:40]
  wire  _GEN_8308 = unuse_way == 2'h2 ? _GEN_3303 : _GEN_7923; // @[d_cache.scala 140:40]
  wire  _GEN_8309 = unuse_way == 2'h2 ? _GEN_3304 : _GEN_7924; // @[d_cache.scala 140:40]
  wire  _GEN_8310 = unuse_way == 2'h2 ? _GEN_3305 : _GEN_7925; // @[d_cache.scala 140:40]
  wire  _GEN_8311 = unuse_way == 2'h2 ? _GEN_3306 : _GEN_7926; // @[d_cache.scala 140:40]
  wire  _GEN_8312 = unuse_way == 2'h2 ? _GEN_3307 : _GEN_7927; // @[d_cache.scala 140:40]
  wire  _GEN_8313 = unuse_way == 2'h2 ? _GEN_3308 : _GEN_7928; // @[d_cache.scala 140:40]
  wire  _GEN_8314 = unuse_way == 2'h2 ? _GEN_3309 : _GEN_7929; // @[d_cache.scala 140:40]
  wire  _GEN_8315 = unuse_way == 2'h2 ? _GEN_3310 : _GEN_7930; // @[d_cache.scala 140:40]
  wire  _GEN_8316 = unuse_way == 2'h2 ? _GEN_3311 : _GEN_7931; // @[d_cache.scala 140:40]
  wire  _GEN_8317 = unuse_way == 2'h2 ? _GEN_3312 : _GEN_7932; // @[d_cache.scala 140:40]
  wire  _GEN_8318 = unuse_way == 2'h2 ? _GEN_3313 : _GEN_7933; // @[d_cache.scala 140:40]
  wire  _GEN_8319 = unuse_way == 2'h2 ? _GEN_3314 : _GEN_7934; // @[d_cache.scala 140:40]
  wire  _GEN_8320 = unuse_way == 2'h2 ? _GEN_3315 : _GEN_7935; // @[d_cache.scala 140:40]
  wire  _GEN_8321 = unuse_way == 2'h2 ? _GEN_3316 : _GEN_7936; // @[d_cache.scala 140:40]
  wire  _GEN_8322 = unuse_way == 2'h2 ? _GEN_3317 : _GEN_7937; // @[d_cache.scala 140:40]
  wire  _GEN_8323 = unuse_way == 2'h2 ? _GEN_3318 : _GEN_7938; // @[d_cache.scala 140:40]
  wire  _GEN_8324 = unuse_way == 2'h2 ? _GEN_3319 : _GEN_7939; // @[d_cache.scala 140:40]
  wire  _GEN_8325 = unuse_way == 2'h2 ? _GEN_3320 : _GEN_7940; // @[d_cache.scala 140:40]
  wire  _GEN_8326 = unuse_way == 2'h2 ? _GEN_3321 : _GEN_7941; // @[d_cache.scala 140:40]
  wire  _GEN_8327 = unuse_way == 2'h2 ? _GEN_3322 : _GEN_7942; // @[d_cache.scala 140:40]
  wire  _GEN_8328 = unuse_way == 2'h2 ? _GEN_3323 : _GEN_7943; // @[d_cache.scala 140:40]
  wire  _GEN_8329 = unuse_way == 2'h2 ? _GEN_3324 : _GEN_7944; // @[d_cache.scala 140:40]
  wire  _GEN_8330 = unuse_way == 2'h2 ? _GEN_3325 : _GEN_7945; // @[d_cache.scala 140:40]
  wire  _GEN_8331 = unuse_way == 2'h2 ? _GEN_3326 : _GEN_7946; // @[d_cache.scala 140:40]
  wire  _GEN_8332 = unuse_way == 2'h2 ? _GEN_3327 : _GEN_7947; // @[d_cache.scala 140:40]
  wire  _GEN_8333 = unuse_way == 2'h2 ? _GEN_3328 : _GEN_7948; // @[d_cache.scala 140:40]
  wire  _GEN_8334 = unuse_way == 2'h2 ? _GEN_3329 : _GEN_7949; // @[d_cache.scala 140:40]
  wire  _GEN_8335 = unuse_way == 2'h2 ? _GEN_3330 : _GEN_7950; // @[d_cache.scala 140:40]
  wire  _GEN_8336 = unuse_way == 2'h2 ? _GEN_3331 : _GEN_7951; // @[d_cache.scala 140:40]
  wire  _GEN_8337 = unuse_way == 2'h2 ? _GEN_3332 : _GEN_7952; // @[d_cache.scala 140:40]
  wire  _GEN_8338 = unuse_way == 2'h2 ? _GEN_3333 : _GEN_7953; // @[d_cache.scala 140:40]
  wire  _GEN_8339 = unuse_way == 2'h2 ? _GEN_3334 : _GEN_7954; // @[d_cache.scala 140:40]
  wire  _GEN_8340 = unuse_way == 2'h2 ? _GEN_3335 : _GEN_7955; // @[d_cache.scala 140:40]
  wire  _GEN_8341 = unuse_way == 2'h2 ? _GEN_3336 : _GEN_7956; // @[d_cache.scala 140:40]
  wire  _GEN_8342 = unuse_way == 2'h2 ? _GEN_3337 : _GEN_7957; // @[d_cache.scala 140:40]
  wire  _GEN_8343 = unuse_way == 2'h2 ? _GEN_3338 : _GEN_7958; // @[d_cache.scala 140:40]
  wire  _GEN_8344 = unuse_way == 2'h2 ? _GEN_3339 : _GEN_7959; // @[d_cache.scala 140:40]
  wire  _GEN_8345 = unuse_way == 2'h2 ? _GEN_3340 : _GEN_7960; // @[d_cache.scala 140:40]
  wire  _GEN_8346 = unuse_way == 2'h2 ? _GEN_3341 : _GEN_7961; // @[d_cache.scala 140:40]
  wire  _GEN_8347 = unuse_way == 2'h2 ? 1'h0 : _T_48; // @[d_cache.scala 140:40 145:23]
  wire [63:0] _GEN_8348 = unuse_way == 2'h2 ? write_back_data : _GEN_6934; // @[d_cache.scala 140:40 29:34]
  wire [41:0] _GEN_8349 = unuse_way == 2'h2 ? {{10'd0}, write_back_addr} : _GEN_6935; // @[d_cache.scala 140:40 30:34]
  wire [63:0] _GEN_8350 = unuse_way == 2'h2 ? ram_0_0 : _GEN_6936; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8351 = unuse_way == 2'h2 ? ram_0_1 : _GEN_6937; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8352 = unuse_way == 2'h2 ? ram_0_2 : _GEN_6938; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8353 = unuse_way == 2'h2 ? ram_0_3 : _GEN_6939; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8354 = unuse_way == 2'h2 ? ram_0_4 : _GEN_6940; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8355 = unuse_way == 2'h2 ? ram_0_5 : _GEN_6941; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8356 = unuse_way == 2'h2 ? ram_0_6 : _GEN_6942; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8357 = unuse_way == 2'h2 ? ram_0_7 : _GEN_6943; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8358 = unuse_way == 2'h2 ? ram_0_8 : _GEN_6944; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8359 = unuse_way == 2'h2 ? ram_0_9 : _GEN_6945; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8360 = unuse_way == 2'h2 ? ram_0_10 : _GEN_6946; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8361 = unuse_way == 2'h2 ? ram_0_11 : _GEN_6947; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8362 = unuse_way == 2'h2 ? ram_0_12 : _GEN_6948; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8363 = unuse_way == 2'h2 ? ram_0_13 : _GEN_6949; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8364 = unuse_way == 2'h2 ? ram_0_14 : _GEN_6950; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8365 = unuse_way == 2'h2 ? ram_0_15 : _GEN_6951; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8366 = unuse_way == 2'h2 ? ram_0_16 : _GEN_6952; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8367 = unuse_way == 2'h2 ? ram_0_17 : _GEN_6953; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8368 = unuse_way == 2'h2 ? ram_0_18 : _GEN_6954; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8369 = unuse_way == 2'h2 ? ram_0_19 : _GEN_6955; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8370 = unuse_way == 2'h2 ? ram_0_20 : _GEN_6956; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8371 = unuse_way == 2'h2 ? ram_0_21 : _GEN_6957; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8372 = unuse_way == 2'h2 ? ram_0_22 : _GEN_6958; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8373 = unuse_way == 2'h2 ? ram_0_23 : _GEN_6959; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8374 = unuse_way == 2'h2 ? ram_0_24 : _GEN_6960; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8375 = unuse_way == 2'h2 ? ram_0_25 : _GEN_6961; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8376 = unuse_way == 2'h2 ? ram_0_26 : _GEN_6962; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8377 = unuse_way == 2'h2 ? ram_0_27 : _GEN_6963; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8378 = unuse_way == 2'h2 ? ram_0_28 : _GEN_6964; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8379 = unuse_way == 2'h2 ? ram_0_29 : _GEN_6965; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8380 = unuse_way == 2'h2 ? ram_0_30 : _GEN_6966; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8381 = unuse_way == 2'h2 ? ram_0_31 : _GEN_6967; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8382 = unuse_way == 2'h2 ? ram_0_32 : _GEN_6968; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8383 = unuse_way == 2'h2 ? ram_0_33 : _GEN_6969; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8384 = unuse_way == 2'h2 ? ram_0_34 : _GEN_6970; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8385 = unuse_way == 2'h2 ? ram_0_35 : _GEN_6971; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8386 = unuse_way == 2'h2 ? ram_0_36 : _GEN_6972; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8387 = unuse_way == 2'h2 ? ram_0_37 : _GEN_6973; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8388 = unuse_way == 2'h2 ? ram_0_38 : _GEN_6974; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8389 = unuse_way == 2'h2 ? ram_0_39 : _GEN_6975; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8390 = unuse_way == 2'h2 ? ram_0_40 : _GEN_6976; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8391 = unuse_way == 2'h2 ? ram_0_41 : _GEN_6977; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8392 = unuse_way == 2'h2 ? ram_0_42 : _GEN_6978; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8393 = unuse_way == 2'h2 ? ram_0_43 : _GEN_6979; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8394 = unuse_way == 2'h2 ? ram_0_44 : _GEN_6980; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8395 = unuse_way == 2'h2 ? ram_0_45 : _GEN_6981; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8396 = unuse_way == 2'h2 ? ram_0_46 : _GEN_6982; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8397 = unuse_way == 2'h2 ? ram_0_47 : _GEN_6983; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8398 = unuse_way == 2'h2 ? ram_0_48 : _GEN_6984; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8399 = unuse_way == 2'h2 ? ram_0_49 : _GEN_6985; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8400 = unuse_way == 2'h2 ? ram_0_50 : _GEN_6986; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8401 = unuse_way == 2'h2 ? ram_0_51 : _GEN_6987; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8402 = unuse_way == 2'h2 ? ram_0_52 : _GEN_6988; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8403 = unuse_way == 2'h2 ? ram_0_53 : _GEN_6989; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8404 = unuse_way == 2'h2 ? ram_0_54 : _GEN_6990; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8405 = unuse_way == 2'h2 ? ram_0_55 : _GEN_6991; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8406 = unuse_way == 2'h2 ? ram_0_56 : _GEN_6992; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8407 = unuse_way == 2'h2 ? ram_0_57 : _GEN_6993; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8408 = unuse_way == 2'h2 ? ram_0_58 : _GEN_6994; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8409 = unuse_way == 2'h2 ? ram_0_59 : _GEN_6995; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8410 = unuse_way == 2'h2 ? ram_0_60 : _GEN_6996; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8411 = unuse_way == 2'h2 ? ram_0_61 : _GEN_6997; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8412 = unuse_way == 2'h2 ? ram_0_62 : _GEN_6998; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8413 = unuse_way == 2'h2 ? ram_0_63 : _GEN_6999; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8414 = unuse_way == 2'h2 ? ram_0_64 : _GEN_7000; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8415 = unuse_way == 2'h2 ? ram_0_65 : _GEN_7001; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8416 = unuse_way == 2'h2 ? ram_0_66 : _GEN_7002; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8417 = unuse_way == 2'h2 ? ram_0_67 : _GEN_7003; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8418 = unuse_way == 2'h2 ? ram_0_68 : _GEN_7004; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8419 = unuse_way == 2'h2 ? ram_0_69 : _GEN_7005; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8420 = unuse_way == 2'h2 ? ram_0_70 : _GEN_7006; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8421 = unuse_way == 2'h2 ? ram_0_71 : _GEN_7007; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8422 = unuse_way == 2'h2 ? ram_0_72 : _GEN_7008; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8423 = unuse_way == 2'h2 ? ram_0_73 : _GEN_7009; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8424 = unuse_way == 2'h2 ? ram_0_74 : _GEN_7010; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8425 = unuse_way == 2'h2 ? ram_0_75 : _GEN_7011; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8426 = unuse_way == 2'h2 ? ram_0_76 : _GEN_7012; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8427 = unuse_way == 2'h2 ? ram_0_77 : _GEN_7013; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8428 = unuse_way == 2'h2 ? ram_0_78 : _GEN_7014; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8429 = unuse_way == 2'h2 ? ram_0_79 : _GEN_7015; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8430 = unuse_way == 2'h2 ? ram_0_80 : _GEN_7016; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8431 = unuse_way == 2'h2 ? ram_0_81 : _GEN_7017; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8432 = unuse_way == 2'h2 ? ram_0_82 : _GEN_7018; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8433 = unuse_way == 2'h2 ? ram_0_83 : _GEN_7019; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8434 = unuse_way == 2'h2 ? ram_0_84 : _GEN_7020; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8435 = unuse_way == 2'h2 ? ram_0_85 : _GEN_7021; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8436 = unuse_way == 2'h2 ? ram_0_86 : _GEN_7022; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8437 = unuse_way == 2'h2 ? ram_0_87 : _GEN_7023; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8438 = unuse_way == 2'h2 ? ram_0_88 : _GEN_7024; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8439 = unuse_way == 2'h2 ? ram_0_89 : _GEN_7025; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8440 = unuse_way == 2'h2 ? ram_0_90 : _GEN_7026; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8441 = unuse_way == 2'h2 ? ram_0_91 : _GEN_7027; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8442 = unuse_way == 2'h2 ? ram_0_92 : _GEN_7028; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8443 = unuse_way == 2'h2 ? ram_0_93 : _GEN_7029; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8444 = unuse_way == 2'h2 ? ram_0_94 : _GEN_7030; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8445 = unuse_way == 2'h2 ? ram_0_95 : _GEN_7031; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8446 = unuse_way == 2'h2 ? ram_0_96 : _GEN_7032; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8447 = unuse_way == 2'h2 ? ram_0_97 : _GEN_7033; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8448 = unuse_way == 2'h2 ? ram_0_98 : _GEN_7034; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8449 = unuse_way == 2'h2 ? ram_0_99 : _GEN_7035; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8450 = unuse_way == 2'h2 ? ram_0_100 : _GEN_7036; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8451 = unuse_way == 2'h2 ? ram_0_101 : _GEN_7037; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8452 = unuse_way == 2'h2 ? ram_0_102 : _GEN_7038; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8453 = unuse_way == 2'h2 ? ram_0_103 : _GEN_7039; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8454 = unuse_way == 2'h2 ? ram_0_104 : _GEN_7040; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8455 = unuse_way == 2'h2 ? ram_0_105 : _GEN_7041; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8456 = unuse_way == 2'h2 ? ram_0_106 : _GEN_7042; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8457 = unuse_way == 2'h2 ? ram_0_107 : _GEN_7043; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8458 = unuse_way == 2'h2 ? ram_0_108 : _GEN_7044; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8459 = unuse_way == 2'h2 ? ram_0_109 : _GEN_7045; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8460 = unuse_way == 2'h2 ? ram_0_110 : _GEN_7046; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8461 = unuse_way == 2'h2 ? ram_0_111 : _GEN_7047; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8462 = unuse_way == 2'h2 ? ram_0_112 : _GEN_7048; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8463 = unuse_way == 2'h2 ? ram_0_113 : _GEN_7049; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8464 = unuse_way == 2'h2 ? ram_0_114 : _GEN_7050; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8465 = unuse_way == 2'h2 ? ram_0_115 : _GEN_7051; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8466 = unuse_way == 2'h2 ? ram_0_116 : _GEN_7052; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8467 = unuse_way == 2'h2 ? ram_0_117 : _GEN_7053; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8468 = unuse_way == 2'h2 ? ram_0_118 : _GEN_7054; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8469 = unuse_way == 2'h2 ? ram_0_119 : _GEN_7055; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8470 = unuse_way == 2'h2 ? ram_0_120 : _GEN_7056; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8471 = unuse_way == 2'h2 ? ram_0_121 : _GEN_7057; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8472 = unuse_way == 2'h2 ? ram_0_122 : _GEN_7058; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8473 = unuse_way == 2'h2 ? ram_0_123 : _GEN_7059; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8474 = unuse_way == 2'h2 ? ram_0_124 : _GEN_7060; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8475 = unuse_way == 2'h2 ? ram_0_125 : _GEN_7061; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8476 = unuse_way == 2'h2 ? ram_0_126 : _GEN_7062; // @[d_cache.scala 140:40 18:24]
  wire [63:0] _GEN_8477 = unuse_way == 2'h2 ? ram_0_127 : _GEN_7063; // @[d_cache.scala 140:40 18:24]
  wire [31:0] _GEN_8478 = unuse_way == 2'h2 ? tag_0_0 : _GEN_7064; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8479 = unuse_way == 2'h2 ? tag_0_1 : _GEN_7065; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8480 = unuse_way == 2'h2 ? tag_0_2 : _GEN_7066; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8481 = unuse_way == 2'h2 ? tag_0_3 : _GEN_7067; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8482 = unuse_way == 2'h2 ? tag_0_4 : _GEN_7068; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8483 = unuse_way == 2'h2 ? tag_0_5 : _GEN_7069; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8484 = unuse_way == 2'h2 ? tag_0_6 : _GEN_7070; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8485 = unuse_way == 2'h2 ? tag_0_7 : _GEN_7071; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8486 = unuse_way == 2'h2 ? tag_0_8 : _GEN_7072; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8487 = unuse_way == 2'h2 ? tag_0_9 : _GEN_7073; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8488 = unuse_way == 2'h2 ? tag_0_10 : _GEN_7074; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8489 = unuse_way == 2'h2 ? tag_0_11 : _GEN_7075; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8490 = unuse_way == 2'h2 ? tag_0_12 : _GEN_7076; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8491 = unuse_way == 2'h2 ? tag_0_13 : _GEN_7077; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8492 = unuse_way == 2'h2 ? tag_0_14 : _GEN_7078; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8493 = unuse_way == 2'h2 ? tag_0_15 : _GEN_7079; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8494 = unuse_way == 2'h2 ? tag_0_16 : _GEN_7080; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8495 = unuse_way == 2'h2 ? tag_0_17 : _GEN_7081; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8496 = unuse_way == 2'h2 ? tag_0_18 : _GEN_7082; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8497 = unuse_way == 2'h2 ? tag_0_19 : _GEN_7083; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8498 = unuse_way == 2'h2 ? tag_0_20 : _GEN_7084; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8499 = unuse_way == 2'h2 ? tag_0_21 : _GEN_7085; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8500 = unuse_way == 2'h2 ? tag_0_22 : _GEN_7086; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8501 = unuse_way == 2'h2 ? tag_0_23 : _GEN_7087; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8502 = unuse_way == 2'h2 ? tag_0_24 : _GEN_7088; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8503 = unuse_way == 2'h2 ? tag_0_25 : _GEN_7089; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8504 = unuse_way == 2'h2 ? tag_0_26 : _GEN_7090; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8505 = unuse_way == 2'h2 ? tag_0_27 : _GEN_7091; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8506 = unuse_way == 2'h2 ? tag_0_28 : _GEN_7092; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8507 = unuse_way == 2'h2 ? tag_0_29 : _GEN_7093; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8508 = unuse_way == 2'h2 ? tag_0_30 : _GEN_7094; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8509 = unuse_way == 2'h2 ? tag_0_31 : _GEN_7095; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8510 = unuse_way == 2'h2 ? tag_0_32 : _GEN_7096; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8511 = unuse_way == 2'h2 ? tag_0_33 : _GEN_7097; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8512 = unuse_way == 2'h2 ? tag_0_34 : _GEN_7098; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8513 = unuse_way == 2'h2 ? tag_0_35 : _GEN_7099; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8514 = unuse_way == 2'h2 ? tag_0_36 : _GEN_7100; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8515 = unuse_way == 2'h2 ? tag_0_37 : _GEN_7101; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8516 = unuse_way == 2'h2 ? tag_0_38 : _GEN_7102; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8517 = unuse_way == 2'h2 ? tag_0_39 : _GEN_7103; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8518 = unuse_way == 2'h2 ? tag_0_40 : _GEN_7104; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8519 = unuse_way == 2'h2 ? tag_0_41 : _GEN_7105; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8520 = unuse_way == 2'h2 ? tag_0_42 : _GEN_7106; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8521 = unuse_way == 2'h2 ? tag_0_43 : _GEN_7107; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8522 = unuse_way == 2'h2 ? tag_0_44 : _GEN_7108; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8523 = unuse_way == 2'h2 ? tag_0_45 : _GEN_7109; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8524 = unuse_way == 2'h2 ? tag_0_46 : _GEN_7110; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8525 = unuse_way == 2'h2 ? tag_0_47 : _GEN_7111; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8526 = unuse_way == 2'h2 ? tag_0_48 : _GEN_7112; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8527 = unuse_way == 2'h2 ? tag_0_49 : _GEN_7113; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8528 = unuse_way == 2'h2 ? tag_0_50 : _GEN_7114; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8529 = unuse_way == 2'h2 ? tag_0_51 : _GEN_7115; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8530 = unuse_way == 2'h2 ? tag_0_52 : _GEN_7116; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8531 = unuse_way == 2'h2 ? tag_0_53 : _GEN_7117; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8532 = unuse_way == 2'h2 ? tag_0_54 : _GEN_7118; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8533 = unuse_way == 2'h2 ? tag_0_55 : _GEN_7119; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8534 = unuse_way == 2'h2 ? tag_0_56 : _GEN_7120; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8535 = unuse_way == 2'h2 ? tag_0_57 : _GEN_7121; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8536 = unuse_way == 2'h2 ? tag_0_58 : _GEN_7122; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8537 = unuse_way == 2'h2 ? tag_0_59 : _GEN_7123; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8538 = unuse_way == 2'h2 ? tag_0_60 : _GEN_7124; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8539 = unuse_way == 2'h2 ? tag_0_61 : _GEN_7125; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8540 = unuse_way == 2'h2 ? tag_0_62 : _GEN_7126; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8541 = unuse_way == 2'h2 ? tag_0_63 : _GEN_7127; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8542 = unuse_way == 2'h2 ? tag_0_64 : _GEN_7128; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8543 = unuse_way == 2'h2 ? tag_0_65 : _GEN_7129; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8544 = unuse_way == 2'h2 ? tag_0_66 : _GEN_7130; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8545 = unuse_way == 2'h2 ? tag_0_67 : _GEN_7131; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8546 = unuse_way == 2'h2 ? tag_0_68 : _GEN_7132; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8547 = unuse_way == 2'h2 ? tag_0_69 : _GEN_7133; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8548 = unuse_way == 2'h2 ? tag_0_70 : _GEN_7134; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8549 = unuse_way == 2'h2 ? tag_0_71 : _GEN_7135; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8550 = unuse_way == 2'h2 ? tag_0_72 : _GEN_7136; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8551 = unuse_way == 2'h2 ? tag_0_73 : _GEN_7137; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8552 = unuse_way == 2'h2 ? tag_0_74 : _GEN_7138; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8553 = unuse_way == 2'h2 ? tag_0_75 : _GEN_7139; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8554 = unuse_way == 2'h2 ? tag_0_76 : _GEN_7140; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8555 = unuse_way == 2'h2 ? tag_0_77 : _GEN_7141; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8556 = unuse_way == 2'h2 ? tag_0_78 : _GEN_7142; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8557 = unuse_way == 2'h2 ? tag_0_79 : _GEN_7143; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8558 = unuse_way == 2'h2 ? tag_0_80 : _GEN_7144; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8559 = unuse_way == 2'h2 ? tag_0_81 : _GEN_7145; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8560 = unuse_way == 2'h2 ? tag_0_82 : _GEN_7146; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8561 = unuse_way == 2'h2 ? tag_0_83 : _GEN_7147; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8562 = unuse_way == 2'h2 ? tag_0_84 : _GEN_7148; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8563 = unuse_way == 2'h2 ? tag_0_85 : _GEN_7149; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8564 = unuse_way == 2'h2 ? tag_0_86 : _GEN_7150; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8565 = unuse_way == 2'h2 ? tag_0_87 : _GEN_7151; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8566 = unuse_way == 2'h2 ? tag_0_88 : _GEN_7152; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8567 = unuse_way == 2'h2 ? tag_0_89 : _GEN_7153; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8568 = unuse_way == 2'h2 ? tag_0_90 : _GEN_7154; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8569 = unuse_way == 2'h2 ? tag_0_91 : _GEN_7155; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8570 = unuse_way == 2'h2 ? tag_0_92 : _GEN_7156; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8571 = unuse_way == 2'h2 ? tag_0_93 : _GEN_7157; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8572 = unuse_way == 2'h2 ? tag_0_94 : _GEN_7158; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8573 = unuse_way == 2'h2 ? tag_0_95 : _GEN_7159; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8574 = unuse_way == 2'h2 ? tag_0_96 : _GEN_7160; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8575 = unuse_way == 2'h2 ? tag_0_97 : _GEN_7161; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8576 = unuse_way == 2'h2 ? tag_0_98 : _GEN_7162; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8577 = unuse_way == 2'h2 ? tag_0_99 : _GEN_7163; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8578 = unuse_way == 2'h2 ? tag_0_100 : _GEN_7164; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8579 = unuse_way == 2'h2 ? tag_0_101 : _GEN_7165; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8580 = unuse_way == 2'h2 ? tag_0_102 : _GEN_7166; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8581 = unuse_way == 2'h2 ? tag_0_103 : _GEN_7167; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8582 = unuse_way == 2'h2 ? tag_0_104 : _GEN_7168; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8583 = unuse_way == 2'h2 ? tag_0_105 : _GEN_7169; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8584 = unuse_way == 2'h2 ? tag_0_106 : _GEN_7170; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8585 = unuse_way == 2'h2 ? tag_0_107 : _GEN_7171; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8586 = unuse_way == 2'h2 ? tag_0_108 : _GEN_7172; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8587 = unuse_way == 2'h2 ? tag_0_109 : _GEN_7173; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8588 = unuse_way == 2'h2 ? tag_0_110 : _GEN_7174; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8589 = unuse_way == 2'h2 ? tag_0_111 : _GEN_7175; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8590 = unuse_way == 2'h2 ? tag_0_112 : _GEN_7176; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8591 = unuse_way == 2'h2 ? tag_0_113 : _GEN_7177; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8592 = unuse_way == 2'h2 ? tag_0_114 : _GEN_7178; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8593 = unuse_way == 2'h2 ? tag_0_115 : _GEN_7179; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8594 = unuse_way == 2'h2 ? tag_0_116 : _GEN_7180; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8595 = unuse_way == 2'h2 ? tag_0_117 : _GEN_7181; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8596 = unuse_way == 2'h2 ? tag_0_118 : _GEN_7182; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8597 = unuse_way == 2'h2 ? tag_0_119 : _GEN_7183; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8598 = unuse_way == 2'h2 ? tag_0_120 : _GEN_7184; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8599 = unuse_way == 2'h2 ? tag_0_121 : _GEN_7185; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8600 = unuse_way == 2'h2 ? tag_0_122 : _GEN_7186; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8601 = unuse_way == 2'h2 ? tag_0_123 : _GEN_7187; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8602 = unuse_way == 2'h2 ? tag_0_124 : _GEN_7188; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8603 = unuse_way == 2'h2 ? tag_0_125 : _GEN_7189; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8604 = unuse_way == 2'h2 ? tag_0_126 : _GEN_7190; // @[d_cache.scala 140:40 20:24]
  wire [31:0] _GEN_8605 = unuse_way == 2'h2 ? tag_0_127 : _GEN_7191; // @[d_cache.scala 140:40 20:24]
  wire  _GEN_8606 = unuse_way == 2'h2 ? dirty_0_0 : _GEN_7192; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8607 = unuse_way == 2'h2 ? dirty_0_1 : _GEN_7193; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8608 = unuse_way == 2'h2 ? dirty_0_2 : _GEN_7194; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8609 = unuse_way == 2'h2 ? dirty_0_3 : _GEN_7195; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8610 = unuse_way == 2'h2 ? dirty_0_4 : _GEN_7196; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8611 = unuse_way == 2'h2 ? dirty_0_5 : _GEN_7197; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8612 = unuse_way == 2'h2 ? dirty_0_6 : _GEN_7198; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8613 = unuse_way == 2'h2 ? dirty_0_7 : _GEN_7199; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8614 = unuse_way == 2'h2 ? dirty_0_8 : _GEN_7200; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8615 = unuse_way == 2'h2 ? dirty_0_9 : _GEN_7201; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8616 = unuse_way == 2'h2 ? dirty_0_10 : _GEN_7202; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8617 = unuse_way == 2'h2 ? dirty_0_11 : _GEN_7203; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8618 = unuse_way == 2'h2 ? dirty_0_12 : _GEN_7204; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8619 = unuse_way == 2'h2 ? dirty_0_13 : _GEN_7205; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8620 = unuse_way == 2'h2 ? dirty_0_14 : _GEN_7206; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8621 = unuse_way == 2'h2 ? dirty_0_15 : _GEN_7207; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8622 = unuse_way == 2'h2 ? dirty_0_16 : _GEN_7208; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8623 = unuse_way == 2'h2 ? dirty_0_17 : _GEN_7209; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8624 = unuse_way == 2'h2 ? dirty_0_18 : _GEN_7210; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8625 = unuse_way == 2'h2 ? dirty_0_19 : _GEN_7211; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8626 = unuse_way == 2'h2 ? dirty_0_20 : _GEN_7212; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8627 = unuse_way == 2'h2 ? dirty_0_21 : _GEN_7213; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8628 = unuse_way == 2'h2 ? dirty_0_22 : _GEN_7214; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8629 = unuse_way == 2'h2 ? dirty_0_23 : _GEN_7215; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8630 = unuse_way == 2'h2 ? dirty_0_24 : _GEN_7216; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8631 = unuse_way == 2'h2 ? dirty_0_25 : _GEN_7217; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8632 = unuse_way == 2'h2 ? dirty_0_26 : _GEN_7218; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8633 = unuse_way == 2'h2 ? dirty_0_27 : _GEN_7219; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8634 = unuse_way == 2'h2 ? dirty_0_28 : _GEN_7220; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8635 = unuse_way == 2'h2 ? dirty_0_29 : _GEN_7221; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8636 = unuse_way == 2'h2 ? dirty_0_30 : _GEN_7222; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8637 = unuse_way == 2'h2 ? dirty_0_31 : _GEN_7223; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8638 = unuse_way == 2'h2 ? dirty_0_32 : _GEN_7224; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8639 = unuse_way == 2'h2 ? dirty_0_33 : _GEN_7225; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8640 = unuse_way == 2'h2 ? dirty_0_34 : _GEN_7226; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8641 = unuse_way == 2'h2 ? dirty_0_35 : _GEN_7227; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8642 = unuse_way == 2'h2 ? dirty_0_36 : _GEN_7228; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8643 = unuse_way == 2'h2 ? dirty_0_37 : _GEN_7229; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8644 = unuse_way == 2'h2 ? dirty_0_38 : _GEN_7230; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8645 = unuse_way == 2'h2 ? dirty_0_39 : _GEN_7231; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8646 = unuse_way == 2'h2 ? dirty_0_40 : _GEN_7232; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8647 = unuse_way == 2'h2 ? dirty_0_41 : _GEN_7233; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8648 = unuse_way == 2'h2 ? dirty_0_42 : _GEN_7234; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8649 = unuse_way == 2'h2 ? dirty_0_43 : _GEN_7235; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8650 = unuse_way == 2'h2 ? dirty_0_44 : _GEN_7236; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8651 = unuse_way == 2'h2 ? dirty_0_45 : _GEN_7237; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8652 = unuse_way == 2'h2 ? dirty_0_46 : _GEN_7238; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8653 = unuse_way == 2'h2 ? dirty_0_47 : _GEN_7239; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8654 = unuse_way == 2'h2 ? dirty_0_48 : _GEN_7240; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8655 = unuse_way == 2'h2 ? dirty_0_49 : _GEN_7241; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8656 = unuse_way == 2'h2 ? dirty_0_50 : _GEN_7242; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8657 = unuse_way == 2'h2 ? dirty_0_51 : _GEN_7243; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8658 = unuse_way == 2'h2 ? dirty_0_52 : _GEN_7244; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8659 = unuse_way == 2'h2 ? dirty_0_53 : _GEN_7245; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8660 = unuse_way == 2'h2 ? dirty_0_54 : _GEN_7246; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8661 = unuse_way == 2'h2 ? dirty_0_55 : _GEN_7247; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8662 = unuse_way == 2'h2 ? dirty_0_56 : _GEN_7248; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8663 = unuse_way == 2'h2 ? dirty_0_57 : _GEN_7249; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8664 = unuse_way == 2'h2 ? dirty_0_58 : _GEN_7250; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8665 = unuse_way == 2'h2 ? dirty_0_59 : _GEN_7251; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8666 = unuse_way == 2'h2 ? dirty_0_60 : _GEN_7252; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8667 = unuse_way == 2'h2 ? dirty_0_61 : _GEN_7253; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8668 = unuse_way == 2'h2 ? dirty_0_62 : _GEN_7254; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8669 = unuse_way == 2'h2 ? dirty_0_63 : _GEN_7255; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8670 = unuse_way == 2'h2 ? dirty_0_64 : _GEN_7256; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8671 = unuse_way == 2'h2 ? dirty_0_65 : _GEN_7257; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8672 = unuse_way == 2'h2 ? dirty_0_66 : _GEN_7258; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8673 = unuse_way == 2'h2 ? dirty_0_67 : _GEN_7259; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8674 = unuse_way == 2'h2 ? dirty_0_68 : _GEN_7260; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8675 = unuse_way == 2'h2 ? dirty_0_69 : _GEN_7261; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8676 = unuse_way == 2'h2 ? dirty_0_70 : _GEN_7262; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8677 = unuse_way == 2'h2 ? dirty_0_71 : _GEN_7263; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8678 = unuse_way == 2'h2 ? dirty_0_72 : _GEN_7264; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8679 = unuse_way == 2'h2 ? dirty_0_73 : _GEN_7265; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8680 = unuse_way == 2'h2 ? dirty_0_74 : _GEN_7266; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8681 = unuse_way == 2'h2 ? dirty_0_75 : _GEN_7267; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8682 = unuse_way == 2'h2 ? dirty_0_76 : _GEN_7268; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8683 = unuse_way == 2'h2 ? dirty_0_77 : _GEN_7269; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8684 = unuse_way == 2'h2 ? dirty_0_78 : _GEN_7270; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8685 = unuse_way == 2'h2 ? dirty_0_79 : _GEN_7271; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8686 = unuse_way == 2'h2 ? dirty_0_80 : _GEN_7272; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8687 = unuse_way == 2'h2 ? dirty_0_81 : _GEN_7273; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8688 = unuse_way == 2'h2 ? dirty_0_82 : _GEN_7274; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8689 = unuse_way == 2'h2 ? dirty_0_83 : _GEN_7275; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8690 = unuse_way == 2'h2 ? dirty_0_84 : _GEN_7276; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8691 = unuse_way == 2'h2 ? dirty_0_85 : _GEN_7277; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8692 = unuse_way == 2'h2 ? dirty_0_86 : _GEN_7278; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8693 = unuse_way == 2'h2 ? dirty_0_87 : _GEN_7279; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8694 = unuse_way == 2'h2 ? dirty_0_88 : _GEN_7280; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8695 = unuse_way == 2'h2 ? dirty_0_89 : _GEN_7281; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8696 = unuse_way == 2'h2 ? dirty_0_90 : _GEN_7282; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8697 = unuse_way == 2'h2 ? dirty_0_91 : _GEN_7283; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8698 = unuse_way == 2'h2 ? dirty_0_92 : _GEN_7284; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8699 = unuse_way == 2'h2 ? dirty_0_93 : _GEN_7285; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8700 = unuse_way == 2'h2 ? dirty_0_94 : _GEN_7286; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8701 = unuse_way == 2'h2 ? dirty_0_95 : _GEN_7287; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8702 = unuse_way == 2'h2 ? dirty_0_96 : _GEN_7288; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8703 = unuse_way == 2'h2 ? dirty_0_97 : _GEN_7289; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8704 = unuse_way == 2'h2 ? dirty_0_98 : _GEN_7290; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8705 = unuse_way == 2'h2 ? dirty_0_99 : _GEN_7291; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8706 = unuse_way == 2'h2 ? dirty_0_100 : _GEN_7292; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8707 = unuse_way == 2'h2 ? dirty_0_101 : _GEN_7293; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8708 = unuse_way == 2'h2 ? dirty_0_102 : _GEN_7294; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8709 = unuse_way == 2'h2 ? dirty_0_103 : _GEN_7295; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8710 = unuse_way == 2'h2 ? dirty_0_104 : _GEN_7296; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8711 = unuse_way == 2'h2 ? dirty_0_105 : _GEN_7297; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8712 = unuse_way == 2'h2 ? dirty_0_106 : _GEN_7298; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8713 = unuse_way == 2'h2 ? dirty_0_107 : _GEN_7299; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8714 = unuse_way == 2'h2 ? dirty_0_108 : _GEN_7300; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8715 = unuse_way == 2'h2 ? dirty_0_109 : _GEN_7301; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8716 = unuse_way == 2'h2 ? dirty_0_110 : _GEN_7302; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8717 = unuse_way == 2'h2 ? dirty_0_111 : _GEN_7303; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8718 = unuse_way == 2'h2 ? dirty_0_112 : _GEN_7304; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8719 = unuse_way == 2'h2 ? dirty_0_113 : _GEN_7305; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8720 = unuse_way == 2'h2 ? dirty_0_114 : _GEN_7306; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8721 = unuse_way == 2'h2 ? dirty_0_115 : _GEN_7307; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8722 = unuse_way == 2'h2 ? dirty_0_116 : _GEN_7308; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8723 = unuse_way == 2'h2 ? dirty_0_117 : _GEN_7309; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8724 = unuse_way == 2'h2 ? dirty_0_118 : _GEN_7310; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8725 = unuse_way == 2'h2 ? dirty_0_119 : _GEN_7311; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8726 = unuse_way == 2'h2 ? dirty_0_120 : _GEN_7312; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8727 = unuse_way == 2'h2 ? dirty_0_121 : _GEN_7313; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8728 = unuse_way == 2'h2 ? dirty_0_122 : _GEN_7314; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8729 = unuse_way == 2'h2 ? dirty_0_123 : _GEN_7315; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8730 = unuse_way == 2'h2 ? dirty_0_124 : _GEN_7316; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8731 = unuse_way == 2'h2 ? dirty_0_125 : _GEN_7317; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8732 = unuse_way == 2'h2 ? dirty_0_126 : _GEN_7318; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8733 = unuse_way == 2'h2 ? dirty_0_127 : _GEN_7319; // @[d_cache.scala 140:40 24:26]
  wire  _GEN_8734 = unuse_way == 2'h2 ? valid_0_0 : _GEN_7320; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8735 = unuse_way == 2'h2 ? valid_0_1 : _GEN_7321; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8736 = unuse_way == 2'h2 ? valid_0_2 : _GEN_7322; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8737 = unuse_way == 2'h2 ? valid_0_3 : _GEN_7323; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8738 = unuse_way == 2'h2 ? valid_0_4 : _GEN_7324; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8739 = unuse_way == 2'h2 ? valid_0_5 : _GEN_7325; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8740 = unuse_way == 2'h2 ? valid_0_6 : _GEN_7326; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8741 = unuse_way == 2'h2 ? valid_0_7 : _GEN_7327; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8742 = unuse_way == 2'h2 ? valid_0_8 : _GEN_7328; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8743 = unuse_way == 2'h2 ? valid_0_9 : _GEN_7329; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8744 = unuse_way == 2'h2 ? valid_0_10 : _GEN_7330; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8745 = unuse_way == 2'h2 ? valid_0_11 : _GEN_7331; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8746 = unuse_way == 2'h2 ? valid_0_12 : _GEN_7332; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8747 = unuse_way == 2'h2 ? valid_0_13 : _GEN_7333; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8748 = unuse_way == 2'h2 ? valid_0_14 : _GEN_7334; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8749 = unuse_way == 2'h2 ? valid_0_15 : _GEN_7335; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8750 = unuse_way == 2'h2 ? valid_0_16 : _GEN_7336; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8751 = unuse_way == 2'h2 ? valid_0_17 : _GEN_7337; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8752 = unuse_way == 2'h2 ? valid_0_18 : _GEN_7338; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8753 = unuse_way == 2'h2 ? valid_0_19 : _GEN_7339; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8754 = unuse_way == 2'h2 ? valid_0_20 : _GEN_7340; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8755 = unuse_way == 2'h2 ? valid_0_21 : _GEN_7341; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8756 = unuse_way == 2'h2 ? valid_0_22 : _GEN_7342; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8757 = unuse_way == 2'h2 ? valid_0_23 : _GEN_7343; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8758 = unuse_way == 2'h2 ? valid_0_24 : _GEN_7344; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8759 = unuse_way == 2'h2 ? valid_0_25 : _GEN_7345; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8760 = unuse_way == 2'h2 ? valid_0_26 : _GEN_7346; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8761 = unuse_way == 2'h2 ? valid_0_27 : _GEN_7347; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8762 = unuse_way == 2'h2 ? valid_0_28 : _GEN_7348; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8763 = unuse_way == 2'h2 ? valid_0_29 : _GEN_7349; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8764 = unuse_way == 2'h2 ? valid_0_30 : _GEN_7350; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8765 = unuse_way == 2'h2 ? valid_0_31 : _GEN_7351; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8766 = unuse_way == 2'h2 ? valid_0_32 : _GEN_7352; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8767 = unuse_way == 2'h2 ? valid_0_33 : _GEN_7353; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8768 = unuse_way == 2'h2 ? valid_0_34 : _GEN_7354; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8769 = unuse_way == 2'h2 ? valid_0_35 : _GEN_7355; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8770 = unuse_way == 2'h2 ? valid_0_36 : _GEN_7356; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8771 = unuse_way == 2'h2 ? valid_0_37 : _GEN_7357; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8772 = unuse_way == 2'h2 ? valid_0_38 : _GEN_7358; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8773 = unuse_way == 2'h2 ? valid_0_39 : _GEN_7359; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8774 = unuse_way == 2'h2 ? valid_0_40 : _GEN_7360; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8775 = unuse_way == 2'h2 ? valid_0_41 : _GEN_7361; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8776 = unuse_way == 2'h2 ? valid_0_42 : _GEN_7362; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8777 = unuse_way == 2'h2 ? valid_0_43 : _GEN_7363; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8778 = unuse_way == 2'h2 ? valid_0_44 : _GEN_7364; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8779 = unuse_way == 2'h2 ? valid_0_45 : _GEN_7365; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8780 = unuse_way == 2'h2 ? valid_0_46 : _GEN_7366; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8781 = unuse_way == 2'h2 ? valid_0_47 : _GEN_7367; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8782 = unuse_way == 2'h2 ? valid_0_48 : _GEN_7368; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8783 = unuse_way == 2'h2 ? valid_0_49 : _GEN_7369; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8784 = unuse_way == 2'h2 ? valid_0_50 : _GEN_7370; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8785 = unuse_way == 2'h2 ? valid_0_51 : _GEN_7371; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8786 = unuse_way == 2'h2 ? valid_0_52 : _GEN_7372; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8787 = unuse_way == 2'h2 ? valid_0_53 : _GEN_7373; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8788 = unuse_way == 2'h2 ? valid_0_54 : _GEN_7374; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8789 = unuse_way == 2'h2 ? valid_0_55 : _GEN_7375; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8790 = unuse_way == 2'h2 ? valid_0_56 : _GEN_7376; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8791 = unuse_way == 2'h2 ? valid_0_57 : _GEN_7377; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8792 = unuse_way == 2'h2 ? valid_0_58 : _GEN_7378; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8793 = unuse_way == 2'h2 ? valid_0_59 : _GEN_7379; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8794 = unuse_way == 2'h2 ? valid_0_60 : _GEN_7380; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8795 = unuse_way == 2'h2 ? valid_0_61 : _GEN_7381; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8796 = unuse_way == 2'h2 ? valid_0_62 : _GEN_7382; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8797 = unuse_way == 2'h2 ? valid_0_63 : _GEN_7383; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8798 = unuse_way == 2'h2 ? valid_0_64 : _GEN_7384; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8799 = unuse_way == 2'h2 ? valid_0_65 : _GEN_7385; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8800 = unuse_way == 2'h2 ? valid_0_66 : _GEN_7386; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8801 = unuse_way == 2'h2 ? valid_0_67 : _GEN_7387; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8802 = unuse_way == 2'h2 ? valid_0_68 : _GEN_7388; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8803 = unuse_way == 2'h2 ? valid_0_69 : _GEN_7389; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8804 = unuse_way == 2'h2 ? valid_0_70 : _GEN_7390; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8805 = unuse_way == 2'h2 ? valid_0_71 : _GEN_7391; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8806 = unuse_way == 2'h2 ? valid_0_72 : _GEN_7392; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8807 = unuse_way == 2'h2 ? valid_0_73 : _GEN_7393; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8808 = unuse_way == 2'h2 ? valid_0_74 : _GEN_7394; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8809 = unuse_way == 2'h2 ? valid_0_75 : _GEN_7395; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8810 = unuse_way == 2'h2 ? valid_0_76 : _GEN_7396; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8811 = unuse_way == 2'h2 ? valid_0_77 : _GEN_7397; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8812 = unuse_way == 2'h2 ? valid_0_78 : _GEN_7398; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8813 = unuse_way == 2'h2 ? valid_0_79 : _GEN_7399; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8814 = unuse_way == 2'h2 ? valid_0_80 : _GEN_7400; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8815 = unuse_way == 2'h2 ? valid_0_81 : _GEN_7401; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8816 = unuse_way == 2'h2 ? valid_0_82 : _GEN_7402; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8817 = unuse_way == 2'h2 ? valid_0_83 : _GEN_7403; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8818 = unuse_way == 2'h2 ? valid_0_84 : _GEN_7404; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8819 = unuse_way == 2'h2 ? valid_0_85 : _GEN_7405; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8820 = unuse_way == 2'h2 ? valid_0_86 : _GEN_7406; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8821 = unuse_way == 2'h2 ? valid_0_87 : _GEN_7407; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8822 = unuse_way == 2'h2 ? valid_0_88 : _GEN_7408; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8823 = unuse_way == 2'h2 ? valid_0_89 : _GEN_7409; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8824 = unuse_way == 2'h2 ? valid_0_90 : _GEN_7410; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8825 = unuse_way == 2'h2 ? valid_0_91 : _GEN_7411; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8826 = unuse_way == 2'h2 ? valid_0_92 : _GEN_7412; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8827 = unuse_way == 2'h2 ? valid_0_93 : _GEN_7413; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8828 = unuse_way == 2'h2 ? valid_0_94 : _GEN_7414; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8829 = unuse_way == 2'h2 ? valid_0_95 : _GEN_7415; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8830 = unuse_way == 2'h2 ? valid_0_96 : _GEN_7416; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8831 = unuse_way == 2'h2 ? valid_0_97 : _GEN_7417; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8832 = unuse_way == 2'h2 ? valid_0_98 : _GEN_7418; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8833 = unuse_way == 2'h2 ? valid_0_99 : _GEN_7419; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8834 = unuse_way == 2'h2 ? valid_0_100 : _GEN_7420; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8835 = unuse_way == 2'h2 ? valid_0_101 : _GEN_7421; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8836 = unuse_way == 2'h2 ? valid_0_102 : _GEN_7422; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8837 = unuse_way == 2'h2 ? valid_0_103 : _GEN_7423; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8838 = unuse_way == 2'h2 ? valid_0_104 : _GEN_7424; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8839 = unuse_way == 2'h2 ? valid_0_105 : _GEN_7425; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8840 = unuse_way == 2'h2 ? valid_0_106 : _GEN_7426; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8841 = unuse_way == 2'h2 ? valid_0_107 : _GEN_7427; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8842 = unuse_way == 2'h2 ? valid_0_108 : _GEN_7428; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8843 = unuse_way == 2'h2 ? valid_0_109 : _GEN_7429; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8844 = unuse_way == 2'h2 ? valid_0_110 : _GEN_7430; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8845 = unuse_way == 2'h2 ? valid_0_111 : _GEN_7431; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8846 = unuse_way == 2'h2 ? valid_0_112 : _GEN_7432; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8847 = unuse_way == 2'h2 ? valid_0_113 : _GEN_7433; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8848 = unuse_way == 2'h2 ? valid_0_114 : _GEN_7434; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8849 = unuse_way == 2'h2 ? valid_0_115 : _GEN_7435; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8850 = unuse_way == 2'h2 ? valid_0_116 : _GEN_7436; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8851 = unuse_way == 2'h2 ? valid_0_117 : _GEN_7437; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8852 = unuse_way == 2'h2 ? valid_0_118 : _GEN_7438; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8853 = unuse_way == 2'h2 ? valid_0_119 : _GEN_7439; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8854 = unuse_way == 2'h2 ? valid_0_120 : _GEN_7440; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8855 = unuse_way == 2'h2 ? valid_0_121 : _GEN_7441; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8856 = unuse_way == 2'h2 ? valid_0_122 : _GEN_7442; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8857 = unuse_way == 2'h2 ? valid_0_123 : _GEN_7443; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8858 = unuse_way == 2'h2 ? valid_0_124 : _GEN_7444; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8859 = unuse_way == 2'h2 ? valid_0_125 : _GEN_7445; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8860 = unuse_way == 2'h2 ? valid_0_126 : _GEN_7446; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8861 = unuse_way == 2'h2 ? valid_0_127 : _GEN_7447; // @[d_cache.scala 140:40 22:26]
  wire  _GEN_8862 = unuse_way == 2'h2 ? dirty_1_0 : _GEN_7706; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8863 = unuse_way == 2'h2 ? dirty_1_1 : _GEN_7707; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8864 = unuse_way == 2'h2 ? dirty_1_2 : _GEN_7708; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8865 = unuse_way == 2'h2 ? dirty_1_3 : _GEN_7709; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8866 = unuse_way == 2'h2 ? dirty_1_4 : _GEN_7710; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8867 = unuse_way == 2'h2 ? dirty_1_5 : _GEN_7711; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8868 = unuse_way == 2'h2 ? dirty_1_6 : _GEN_7712; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8869 = unuse_way == 2'h2 ? dirty_1_7 : _GEN_7713; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8870 = unuse_way == 2'h2 ? dirty_1_8 : _GEN_7714; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8871 = unuse_way == 2'h2 ? dirty_1_9 : _GEN_7715; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8872 = unuse_way == 2'h2 ? dirty_1_10 : _GEN_7716; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8873 = unuse_way == 2'h2 ? dirty_1_11 : _GEN_7717; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8874 = unuse_way == 2'h2 ? dirty_1_12 : _GEN_7718; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8875 = unuse_way == 2'h2 ? dirty_1_13 : _GEN_7719; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8876 = unuse_way == 2'h2 ? dirty_1_14 : _GEN_7720; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8877 = unuse_way == 2'h2 ? dirty_1_15 : _GEN_7721; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8878 = unuse_way == 2'h2 ? dirty_1_16 : _GEN_7722; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8879 = unuse_way == 2'h2 ? dirty_1_17 : _GEN_7723; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8880 = unuse_way == 2'h2 ? dirty_1_18 : _GEN_7724; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8881 = unuse_way == 2'h2 ? dirty_1_19 : _GEN_7725; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8882 = unuse_way == 2'h2 ? dirty_1_20 : _GEN_7726; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8883 = unuse_way == 2'h2 ? dirty_1_21 : _GEN_7727; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8884 = unuse_way == 2'h2 ? dirty_1_22 : _GEN_7728; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8885 = unuse_way == 2'h2 ? dirty_1_23 : _GEN_7729; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8886 = unuse_way == 2'h2 ? dirty_1_24 : _GEN_7730; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8887 = unuse_way == 2'h2 ? dirty_1_25 : _GEN_7731; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8888 = unuse_way == 2'h2 ? dirty_1_26 : _GEN_7732; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8889 = unuse_way == 2'h2 ? dirty_1_27 : _GEN_7733; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8890 = unuse_way == 2'h2 ? dirty_1_28 : _GEN_7734; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8891 = unuse_way == 2'h2 ? dirty_1_29 : _GEN_7735; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8892 = unuse_way == 2'h2 ? dirty_1_30 : _GEN_7736; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8893 = unuse_way == 2'h2 ? dirty_1_31 : _GEN_7737; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8894 = unuse_way == 2'h2 ? dirty_1_32 : _GEN_7738; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8895 = unuse_way == 2'h2 ? dirty_1_33 : _GEN_7739; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8896 = unuse_way == 2'h2 ? dirty_1_34 : _GEN_7740; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8897 = unuse_way == 2'h2 ? dirty_1_35 : _GEN_7741; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8898 = unuse_way == 2'h2 ? dirty_1_36 : _GEN_7742; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8899 = unuse_way == 2'h2 ? dirty_1_37 : _GEN_7743; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8900 = unuse_way == 2'h2 ? dirty_1_38 : _GEN_7744; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8901 = unuse_way == 2'h2 ? dirty_1_39 : _GEN_7745; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8902 = unuse_way == 2'h2 ? dirty_1_40 : _GEN_7746; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8903 = unuse_way == 2'h2 ? dirty_1_41 : _GEN_7747; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8904 = unuse_way == 2'h2 ? dirty_1_42 : _GEN_7748; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8905 = unuse_way == 2'h2 ? dirty_1_43 : _GEN_7749; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8906 = unuse_way == 2'h2 ? dirty_1_44 : _GEN_7750; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8907 = unuse_way == 2'h2 ? dirty_1_45 : _GEN_7751; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8908 = unuse_way == 2'h2 ? dirty_1_46 : _GEN_7752; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8909 = unuse_way == 2'h2 ? dirty_1_47 : _GEN_7753; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8910 = unuse_way == 2'h2 ? dirty_1_48 : _GEN_7754; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8911 = unuse_way == 2'h2 ? dirty_1_49 : _GEN_7755; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8912 = unuse_way == 2'h2 ? dirty_1_50 : _GEN_7756; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8913 = unuse_way == 2'h2 ? dirty_1_51 : _GEN_7757; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8914 = unuse_way == 2'h2 ? dirty_1_52 : _GEN_7758; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8915 = unuse_way == 2'h2 ? dirty_1_53 : _GEN_7759; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8916 = unuse_way == 2'h2 ? dirty_1_54 : _GEN_7760; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8917 = unuse_way == 2'h2 ? dirty_1_55 : _GEN_7761; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8918 = unuse_way == 2'h2 ? dirty_1_56 : _GEN_7762; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8919 = unuse_way == 2'h2 ? dirty_1_57 : _GEN_7763; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8920 = unuse_way == 2'h2 ? dirty_1_58 : _GEN_7764; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8921 = unuse_way == 2'h2 ? dirty_1_59 : _GEN_7765; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8922 = unuse_way == 2'h2 ? dirty_1_60 : _GEN_7766; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8923 = unuse_way == 2'h2 ? dirty_1_61 : _GEN_7767; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8924 = unuse_way == 2'h2 ? dirty_1_62 : _GEN_7768; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8925 = unuse_way == 2'h2 ? dirty_1_63 : _GEN_7769; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8926 = unuse_way == 2'h2 ? dirty_1_64 : _GEN_7770; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8927 = unuse_way == 2'h2 ? dirty_1_65 : _GEN_7771; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8928 = unuse_way == 2'h2 ? dirty_1_66 : _GEN_7772; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8929 = unuse_way == 2'h2 ? dirty_1_67 : _GEN_7773; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8930 = unuse_way == 2'h2 ? dirty_1_68 : _GEN_7774; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8931 = unuse_way == 2'h2 ? dirty_1_69 : _GEN_7775; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8932 = unuse_way == 2'h2 ? dirty_1_70 : _GEN_7776; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8933 = unuse_way == 2'h2 ? dirty_1_71 : _GEN_7777; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8934 = unuse_way == 2'h2 ? dirty_1_72 : _GEN_7778; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8935 = unuse_way == 2'h2 ? dirty_1_73 : _GEN_7779; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8936 = unuse_way == 2'h2 ? dirty_1_74 : _GEN_7780; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8937 = unuse_way == 2'h2 ? dirty_1_75 : _GEN_7781; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8938 = unuse_way == 2'h2 ? dirty_1_76 : _GEN_7782; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8939 = unuse_way == 2'h2 ? dirty_1_77 : _GEN_7783; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8940 = unuse_way == 2'h2 ? dirty_1_78 : _GEN_7784; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8941 = unuse_way == 2'h2 ? dirty_1_79 : _GEN_7785; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8942 = unuse_way == 2'h2 ? dirty_1_80 : _GEN_7786; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8943 = unuse_way == 2'h2 ? dirty_1_81 : _GEN_7787; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8944 = unuse_way == 2'h2 ? dirty_1_82 : _GEN_7788; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8945 = unuse_way == 2'h2 ? dirty_1_83 : _GEN_7789; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8946 = unuse_way == 2'h2 ? dirty_1_84 : _GEN_7790; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8947 = unuse_way == 2'h2 ? dirty_1_85 : _GEN_7791; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8948 = unuse_way == 2'h2 ? dirty_1_86 : _GEN_7792; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8949 = unuse_way == 2'h2 ? dirty_1_87 : _GEN_7793; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8950 = unuse_way == 2'h2 ? dirty_1_88 : _GEN_7794; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8951 = unuse_way == 2'h2 ? dirty_1_89 : _GEN_7795; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8952 = unuse_way == 2'h2 ? dirty_1_90 : _GEN_7796; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8953 = unuse_way == 2'h2 ? dirty_1_91 : _GEN_7797; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8954 = unuse_way == 2'h2 ? dirty_1_92 : _GEN_7798; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8955 = unuse_way == 2'h2 ? dirty_1_93 : _GEN_7799; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8956 = unuse_way == 2'h2 ? dirty_1_94 : _GEN_7800; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8957 = unuse_way == 2'h2 ? dirty_1_95 : _GEN_7801; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8958 = unuse_way == 2'h2 ? dirty_1_96 : _GEN_7802; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8959 = unuse_way == 2'h2 ? dirty_1_97 : _GEN_7803; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8960 = unuse_way == 2'h2 ? dirty_1_98 : _GEN_7804; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8961 = unuse_way == 2'h2 ? dirty_1_99 : _GEN_7805; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8962 = unuse_way == 2'h2 ? dirty_1_100 : _GEN_7806; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8963 = unuse_way == 2'h2 ? dirty_1_101 : _GEN_7807; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8964 = unuse_way == 2'h2 ? dirty_1_102 : _GEN_7808; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8965 = unuse_way == 2'h2 ? dirty_1_103 : _GEN_7809; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8966 = unuse_way == 2'h2 ? dirty_1_104 : _GEN_7810; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8967 = unuse_way == 2'h2 ? dirty_1_105 : _GEN_7811; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8968 = unuse_way == 2'h2 ? dirty_1_106 : _GEN_7812; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8969 = unuse_way == 2'h2 ? dirty_1_107 : _GEN_7813; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8970 = unuse_way == 2'h2 ? dirty_1_108 : _GEN_7814; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8971 = unuse_way == 2'h2 ? dirty_1_109 : _GEN_7815; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8972 = unuse_way == 2'h2 ? dirty_1_110 : _GEN_7816; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8973 = unuse_way == 2'h2 ? dirty_1_111 : _GEN_7817; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8974 = unuse_way == 2'h2 ? dirty_1_112 : _GEN_7818; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8975 = unuse_way == 2'h2 ? dirty_1_113 : _GEN_7819; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8976 = unuse_way == 2'h2 ? dirty_1_114 : _GEN_7820; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8977 = unuse_way == 2'h2 ? dirty_1_115 : _GEN_7821; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8978 = unuse_way == 2'h2 ? dirty_1_116 : _GEN_7822; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8979 = unuse_way == 2'h2 ? dirty_1_117 : _GEN_7823; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8980 = unuse_way == 2'h2 ? dirty_1_118 : _GEN_7824; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8981 = unuse_way == 2'h2 ? dirty_1_119 : _GEN_7825; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8982 = unuse_way == 2'h2 ? dirty_1_120 : _GEN_7826; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8983 = unuse_way == 2'h2 ? dirty_1_121 : _GEN_7827; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8984 = unuse_way == 2'h2 ? dirty_1_122 : _GEN_7828; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8985 = unuse_way == 2'h2 ? dirty_1_123 : _GEN_7829; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8986 = unuse_way == 2'h2 ? dirty_1_124 : _GEN_7830; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8987 = unuse_way == 2'h2 ? dirty_1_125 : _GEN_7831; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8988 = unuse_way == 2'h2 ? dirty_1_126 : _GEN_7832; // @[d_cache.scala 140:40 25:26]
  wire  _GEN_8989 = unuse_way == 2'h2 ? dirty_1_127 : _GEN_7833; // @[d_cache.scala 140:40 25:26]
  wire [2:0] _GEN_8990 = unuse_way == 2'h1 ? 3'h7 : _GEN_7962; // @[d_cache.scala 134:34 135:23]
  wire [63:0] _GEN_8991 = unuse_way == 2'h1 ? _GEN_2574 : _GEN_8350; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_8992 = unuse_way == 2'h1 ? _GEN_2575 : _GEN_8351; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_8993 = unuse_way == 2'h1 ? _GEN_2576 : _GEN_8352; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_8994 = unuse_way == 2'h1 ? _GEN_2577 : _GEN_8353; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_8995 = unuse_way == 2'h1 ? _GEN_2578 : _GEN_8354; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_8996 = unuse_way == 2'h1 ? _GEN_2579 : _GEN_8355; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_8997 = unuse_way == 2'h1 ? _GEN_2580 : _GEN_8356; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_8998 = unuse_way == 2'h1 ? _GEN_2581 : _GEN_8357; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_8999 = unuse_way == 2'h1 ? _GEN_2582 : _GEN_8358; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9000 = unuse_way == 2'h1 ? _GEN_2583 : _GEN_8359; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9001 = unuse_way == 2'h1 ? _GEN_2584 : _GEN_8360; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9002 = unuse_way == 2'h1 ? _GEN_2585 : _GEN_8361; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9003 = unuse_way == 2'h1 ? _GEN_2586 : _GEN_8362; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9004 = unuse_way == 2'h1 ? _GEN_2587 : _GEN_8363; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9005 = unuse_way == 2'h1 ? _GEN_2588 : _GEN_8364; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9006 = unuse_way == 2'h1 ? _GEN_2589 : _GEN_8365; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9007 = unuse_way == 2'h1 ? _GEN_2590 : _GEN_8366; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9008 = unuse_way == 2'h1 ? _GEN_2591 : _GEN_8367; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9009 = unuse_way == 2'h1 ? _GEN_2592 : _GEN_8368; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9010 = unuse_way == 2'h1 ? _GEN_2593 : _GEN_8369; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9011 = unuse_way == 2'h1 ? _GEN_2594 : _GEN_8370; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9012 = unuse_way == 2'h1 ? _GEN_2595 : _GEN_8371; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9013 = unuse_way == 2'h1 ? _GEN_2596 : _GEN_8372; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9014 = unuse_way == 2'h1 ? _GEN_2597 : _GEN_8373; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9015 = unuse_way == 2'h1 ? _GEN_2598 : _GEN_8374; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9016 = unuse_way == 2'h1 ? _GEN_2599 : _GEN_8375; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9017 = unuse_way == 2'h1 ? _GEN_2600 : _GEN_8376; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9018 = unuse_way == 2'h1 ? _GEN_2601 : _GEN_8377; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9019 = unuse_way == 2'h1 ? _GEN_2602 : _GEN_8378; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9020 = unuse_way == 2'h1 ? _GEN_2603 : _GEN_8379; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9021 = unuse_way == 2'h1 ? _GEN_2604 : _GEN_8380; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9022 = unuse_way == 2'h1 ? _GEN_2605 : _GEN_8381; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9023 = unuse_way == 2'h1 ? _GEN_2606 : _GEN_8382; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9024 = unuse_way == 2'h1 ? _GEN_2607 : _GEN_8383; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9025 = unuse_way == 2'h1 ? _GEN_2608 : _GEN_8384; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9026 = unuse_way == 2'h1 ? _GEN_2609 : _GEN_8385; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9027 = unuse_way == 2'h1 ? _GEN_2610 : _GEN_8386; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9028 = unuse_way == 2'h1 ? _GEN_2611 : _GEN_8387; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9029 = unuse_way == 2'h1 ? _GEN_2612 : _GEN_8388; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9030 = unuse_way == 2'h1 ? _GEN_2613 : _GEN_8389; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9031 = unuse_way == 2'h1 ? _GEN_2614 : _GEN_8390; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9032 = unuse_way == 2'h1 ? _GEN_2615 : _GEN_8391; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9033 = unuse_way == 2'h1 ? _GEN_2616 : _GEN_8392; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9034 = unuse_way == 2'h1 ? _GEN_2617 : _GEN_8393; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9035 = unuse_way == 2'h1 ? _GEN_2618 : _GEN_8394; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9036 = unuse_way == 2'h1 ? _GEN_2619 : _GEN_8395; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9037 = unuse_way == 2'h1 ? _GEN_2620 : _GEN_8396; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9038 = unuse_way == 2'h1 ? _GEN_2621 : _GEN_8397; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9039 = unuse_way == 2'h1 ? _GEN_2622 : _GEN_8398; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9040 = unuse_way == 2'h1 ? _GEN_2623 : _GEN_8399; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9041 = unuse_way == 2'h1 ? _GEN_2624 : _GEN_8400; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9042 = unuse_way == 2'h1 ? _GEN_2625 : _GEN_8401; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9043 = unuse_way == 2'h1 ? _GEN_2626 : _GEN_8402; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9044 = unuse_way == 2'h1 ? _GEN_2627 : _GEN_8403; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9045 = unuse_way == 2'h1 ? _GEN_2628 : _GEN_8404; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9046 = unuse_way == 2'h1 ? _GEN_2629 : _GEN_8405; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9047 = unuse_way == 2'h1 ? _GEN_2630 : _GEN_8406; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9048 = unuse_way == 2'h1 ? _GEN_2631 : _GEN_8407; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9049 = unuse_way == 2'h1 ? _GEN_2632 : _GEN_8408; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9050 = unuse_way == 2'h1 ? _GEN_2633 : _GEN_8409; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9051 = unuse_way == 2'h1 ? _GEN_2634 : _GEN_8410; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9052 = unuse_way == 2'h1 ? _GEN_2635 : _GEN_8411; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9053 = unuse_way == 2'h1 ? _GEN_2636 : _GEN_8412; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9054 = unuse_way == 2'h1 ? _GEN_2637 : _GEN_8413; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9055 = unuse_way == 2'h1 ? _GEN_2638 : _GEN_8414; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9056 = unuse_way == 2'h1 ? _GEN_2639 : _GEN_8415; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9057 = unuse_way == 2'h1 ? _GEN_2640 : _GEN_8416; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9058 = unuse_way == 2'h1 ? _GEN_2641 : _GEN_8417; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9059 = unuse_way == 2'h1 ? _GEN_2642 : _GEN_8418; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9060 = unuse_way == 2'h1 ? _GEN_2643 : _GEN_8419; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9061 = unuse_way == 2'h1 ? _GEN_2644 : _GEN_8420; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9062 = unuse_way == 2'h1 ? _GEN_2645 : _GEN_8421; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9063 = unuse_way == 2'h1 ? _GEN_2646 : _GEN_8422; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9064 = unuse_way == 2'h1 ? _GEN_2647 : _GEN_8423; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9065 = unuse_way == 2'h1 ? _GEN_2648 : _GEN_8424; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9066 = unuse_way == 2'h1 ? _GEN_2649 : _GEN_8425; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9067 = unuse_way == 2'h1 ? _GEN_2650 : _GEN_8426; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9068 = unuse_way == 2'h1 ? _GEN_2651 : _GEN_8427; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9069 = unuse_way == 2'h1 ? _GEN_2652 : _GEN_8428; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9070 = unuse_way == 2'h1 ? _GEN_2653 : _GEN_8429; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9071 = unuse_way == 2'h1 ? _GEN_2654 : _GEN_8430; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9072 = unuse_way == 2'h1 ? _GEN_2655 : _GEN_8431; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9073 = unuse_way == 2'h1 ? _GEN_2656 : _GEN_8432; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9074 = unuse_way == 2'h1 ? _GEN_2657 : _GEN_8433; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9075 = unuse_way == 2'h1 ? _GEN_2658 : _GEN_8434; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9076 = unuse_way == 2'h1 ? _GEN_2659 : _GEN_8435; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9077 = unuse_way == 2'h1 ? _GEN_2660 : _GEN_8436; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9078 = unuse_way == 2'h1 ? _GEN_2661 : _GEN_8437; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9079 = unuse_way == 2'h1 ? _GEN_2662 : _GEN_8438; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9080 = unuse_way == 2'h1 ? _GEN_2663 : _GEN_8439; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9081 = unuse_way == 2'h1 ? _GEN_2664 : _GEN_8440; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9082 = unuse_way == 2'h1 ? _GEN_2665 : _GEN_8441; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9083 = unuse_way == 2'h1 ? _GEN_2666 : _GEN_8442; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9084 = unuse_way == 2'h1 ? _GEN_2667 : _GEN_8443; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9085 = unuse_way == 2'h1 ? _GEN_2668 : _GEN_8444; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9086 = unuse_way == 2'h1 ? _GEN_2669 : _GEN_8445; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9087 = unuse_way == 2'h1 ? _GEN_2670 : _GEN_8446; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9088 = unuse_way == 2'h1 ? _GEN_2671 : _GEN_8447; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9089 = unuse_way == 2'h1 ? _GEN_2672 : _GEN_8448; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9090 = unuse_way == 2'h1 ? _GEN_2673 : _GEN_8449; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9091 = unuse_way == 2'h1 ? _GEN_2674 : _GEN_8450; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9092 = unuse_way == 2'h1 ? _GEN_2675 : _GEN_8451; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9093 = unuse_way == 2'h1 ? _GEN_2676 : _GEN_8452; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9094 = unuse_way == 2'h1 ? _GEN_2677 : _GEN_8453; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9095 = unuse_way == 2'h1 ? _GEN_2678 : _GEN_8454; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9096 = unuse_way == 2'h1 ? _GEN_2679 : _GEN_8455; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9097 = unuse_way == 2'h1 ? _GEN_2680 : _GEN_8456; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9098 = unuse_way == 2'h1 ? _GEN_2681 : _GEN_8457; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9099 = unuse_way == 2'h1 ? _GEN_2682 : _GEN_8458; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9100 = unuse_way == 2'h1 ? _GEN_2683 : _GEN_8459; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9101 = unuse_way == 2'h1 ? _GEN_2684 : _GEN_8460; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9102 = unuse_way == 2'h1 ? _GEN_2685 : _GEN_8461; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9103 = unuse_way == 2'h1 ? _GEN_2686 : _GEN_8462; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9104 = unuse_way == 2'h1 ? _GEN_2687 : _GEN_8463; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9105 = unuse_way == 2'h1 ? _GEN_2688 : _GEN_8464; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9106 = unuse_way == 2'h1 ? _GEN_2689 : _GEN_8465; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9107 = unuse_way == 2'h1 ? _GEN_2690 : _GEN_8466; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9108 = unuse_way == 2'h1 ? _GEN_2691 : _GEN_8467; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9109 = unuse_way == 2'h1 ? _GEN_2692 : _GEN_8468; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9110 = unuse_way == 2'h1 ? _GEN_2693 : _GEN_8469; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9111 = unuse_way == 2'h1 ? _GEN_2694 : _GEN_8470; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9112 = unuse_way == 2'h1 ? _GEN_2695 : _GEN_8471; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9113 = unuse_way == 2'h1 ? _GEN_2696 : _GEN_8472; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9114 = unuse_way == 2'h1 ? _GEN_2697 : _GEN_8473; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9115 = unuse_way == 2'h1 ? _GEN_2698 : _GEN_8474; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9116 = unuse_way == 2'h1 ? _GEN_2699 : _GEN_8475; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9117 = unuse_way == 2'h1 ? _GEN_2700 : _GEN_8476; // @[d_cache.scala 134:34]
  wire [63:0] _GEN_9118 = unuse_way == 2'h1 ? _GEN_2701 : _GEN_8477; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9119 = unuse_way == 2'h1 ? _GEN_2702 : _GEN_8478; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9120 = unuse_way == 2'h1 ? _GEN_2703 : _GEN_8479; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9121 = unuse_way == 2'h1 ? _GEN_2704 : _GEN_8480; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9122 = unuse_way == 2'h1 ? _GEN_2705 : _GEN_8481; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9123 = unuse_way == 2'h1 ? _GEN_2706 : _GEN_8482; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9124 = unuse_way == 2'h1 ? _GEN_2707 : _GEN_8483; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9125 = unuse_way == 2'h1 ? _GEN_2708 : _GEN_8484; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9126 = unuse_way == 2'h1 ? _GEN_2709 : _GEN_8485; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9127 = unuse_way == 2'h1 ? _GEN_2710 : _GEN_8486; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9128 = unuse_way == 2'h1 ? _GEN_2711 : _GEN_8487; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9129 = unuse_way == 2'h1 ? _GEN_2712 : _GEN_8488; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9130 = unuse_way == 2'h1 ? _GEN_2713 : _GEN_8489; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9131 = unuse_way == 2'h1 ? _GEN_2714 : _GEN_8490; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9132 = unuse_way == 2'h1 ? _GEN_2715 : _GEN_8491; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9133 = unuse_way == 2'h1 ? _GEN_2716 : _GEN_8492; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9134 = unuse_way == 2'h1 ? _GEN_2717 : _GEN_8493; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9135 = unuse_way == 2'h1 ? _GEN_2718 : _GEN_8494; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9136 = unuse_way == 2'h1 ? _GEN_2719 : _GEN_8495; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9137 = unuse_way == 2'h1 ? _GEN_2720 : _GEN_8496; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9138 = unuse_way == 2'h1 ? _GEN_2721 : _GEN_8497; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9139 = unuse_way == 2'h1 ? _GEN_2722 : _GEN_8498; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9140 = unuse_way == 2'h1 ? _GEN_2723 : _GEN_8499; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9141 = unuse_way == 2'h1 ? _GEN_2724 : _GEN_8500; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9142 = unuse_way == 2'h1 ? _GEN_2725 : _GEN_8501; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9143 = unuse_way == 2'h1 ? _GEN_2726 : _GEN_8502; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9144 = unuse_way == 2'h1 ? _GEN_2727 : _GEN_8503; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9145 = unuse_way == 2'h1 ? _GEN_2728 : _GEN_8504; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9146 = unuse_way == 2'h1 ? _GEN_2729 : _GEN_8505; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9147 = unuse_way == 2'h1 ? _GEN_2730 : _GEN_8506; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9148 = unuse_way == 2'h1 ? _GEN_2731 : _GEN_8507; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9149 = unuse_way == 2'h1 ? _GEN_2732 : _GEN_8508; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9150 = unuse_way == 2'h1 ? _GEN_2733 : _GEN_8509; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9151 = unuse_way == 2'h1 ? _GEN_2734 : _GEN_8510; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9152 = unuse_way == 2'h1 ? _GEN_2735 : _GEN_8511; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9153 = unuse_way == 2'h1 ? _GEN_2736 : _GEN_8512; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9154 = unuse_way == 2'h1 ? _GEN_2737 : _GEN_8513; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9155 = unuse_way == 2'h1 ? _GEN_2738 : _GEN_8514; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9156 = unuse_way == 2'h1 ? _GEN_2739 : _GEN_8515; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9157 = unuse_way == 2'h1 ? _GEN_2740 : _GEN_8516; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9158 = unuse_way == 2'h1 ? _GEN_2741 : _GEN_8517; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9159 = unuse_way == 2'h1 ? _GEN_2742 : _GEN_8518; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9160 = unuse_way == 2'h1 ? _GEN_2743 : _GEN_8519; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9161 = unuse_way == 2'h1 ? _GEN_2744 : _GEN_8520; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9162 = unuse_way == 2'h1 ? _GEN_2745 : _GEN_8521; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9163 = unuse_way == 2'h1 ? _GEN_2746 : _GEN_8522; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9164 = unuse_way == 2'h1 ? _GEN_2747 : _GEN_8523; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9165 = unuse_way == 2'h1 ? _GEN_2748 : _GEN_8524; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9166 = unuse_way == 2'h1 ? _GEN_2749 : _GEN_8525; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9167 = unuse_way == 2'h1 ? _GEN_2750 : _GEN_8526; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9168 = unuse_way == 2'h1 ? _GEN_2751 : _GEN_8527; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9169 = unuse_way == 2'h1 ? _GEN_2752 : _GEN_8528; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9170 = unuse_way == 2'h1 ? _GEN_2753 : _GEN_8529; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9171 = unuse_way == 2'h1 ? _GEN_2754 : _GEN_8530; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9172 = unuse_way == 2'h1 ? _GEN_2755 : _GEN_8531; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9173 = unuse_way == 2'h1 ? _GEN_2756 : _GEN_8532; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9174 = unuse_way == 2'h1 ? _GEN_2757 : _GEN_8533; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9175 = unuse_way == 2'h1 ? _GEN_2758 : _GEN_8534; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9176 = unuse_way == 2'h1 ? _GEN_2759 : _GEN_8535; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9177 = unuse_way == 2'h1 ? _GEN_2760 : _GEN_8536; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9178 = unuse_way == 2'h1 ? _GEN_2761 : _GEN_8537; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9179 = unuse_way == 2'h1 ? _GEN_2762 : _GEN_8538; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9180 = unuse_way == 2'h1 ? _GEN_2763 : _GEN_8539; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9181 = unuse_way == 2'h1 ? _GEN_2764 : _GEN_8540; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9182 = unuse_way == 2'h1 ? _GEN_2765 : _GEN_8541; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9183 = unuse_way == 2'h1 ? _GEN_2766 : _GEN_8542; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9184 = unuse_way == 2'h1 ? _GEN_2767 : _GEN_8543; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9185 = unuse_way == 2'h1 ? _GEN_2768 : _GEN_8544; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9186 = unuse_way == 2'h1 ? _GEN_2769 : _GEN_8545; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9187 = unuse_way == 2'h1 ? _GEN_2770 : _GEN_8546; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9188 = unuse_way == 2'h1 ? _GEN_2771 : _GEN_8547; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9189 = unuse_way == 2'h1 ? _GEN_2772 : _GEN_8548; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9190 = unuse_way == 2'h1 ? _GEN_2773 : _GEN_8549; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9191 = unuse_way == 2'h1 ? _GEN_2774 : _GEN_8550; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9192 = unuse_way == 2'h1 ? _GEN_2775 : _GEN_8551; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9193 = unuse_way == 2'h1 ? _GEN_2776 : _GEN_8552; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9194 = unuse_way == 2'h1 ? _GEN_2777 : _GEN_8553; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9195 = unuse_way == 2'h1 ? _GEN_2778 : _GEN_8554; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9196 = unuse_way == 2'h1 ? _GEN_2779 : _GEN_8555; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9197 = unuse_way == 2'h1 ? _GEN_2780 : _GEN_8556; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9198 = unuse_way == 2'h1 ? _GEN_2781 : _GEN_8557; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9199 = unuse_way == 2'h1 ? _GEN_2782 : _GEN_8558; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9200 = unuse_way == 2'h1 ? _GEN_2783 : _GEN_8559; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9201 = unuse_way == 2'h1 ? _GEN_2784 : _GEN_8560; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9202 = unuse_way == 2'h1 ? _GEN_2785 : _GEN_8561; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9203 = unuse_way == 2'h1 ? _GEN_2786 : _GEN_8562; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9204 = unuse_way == 2'h1 ? _GEN_2787 : _GEN_8563; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9205 = unuse_way == 2'h1 ? _GEN_2788 : _GEN_8564; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9206 = unuse_way == 2'h1 ? _GEN_2789 : _GEN_8565; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9207 = unuse_way == 2'h1 ? _GEN_2790 : _GEN_8566; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9208 = unuse_way == 2'h1 ? _GEN_2791 : _GEN_8567; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9209 = unuse_way == 2'h1 ? _GEN_2792 : _GEN_8568; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9210 = unuse_way == 2'h1 ? _GEN_2793 : _GEN_8569; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9211 = unuse_way == 2'h1 ? _GEN_2794 : _GEN_8570; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9212 = unuse_way == 2'h1 ? _GEN_2795 : _GEN_8571; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9213 = unuse_way == 2'h1 ? _GEN_2796 : _GEN_8572; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9214 = unuse_way == 2'h1 ? _GEN_2797 : _GEN_8573; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9215 = unuse_way == 2'h1 ? _GEN_2798 : _GEN_8574; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9216 = unuse_way == 2'h1 ? _GEN_2799 : _GEN_8575; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9217 = unuse_way == 2'h1 ? _GEN_2800 : _GEN_8576; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9218 = unuse_way == 2'h1 ? _GEN_2801 : _GEN_8577; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9219 = unuse_way == 2'h1 ? _GEN_2802 : _GEN_8578; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9220 = unuse_way == 2'h1 ? _GEN_2803 : _GEN_8579; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9221 = unuse_way == 2'h1 ? _GEN_2804 : _GEN_8580; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9222 = unuse_way == 2'h1 ? _GEN_2805 : _GEN_8581; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9223 = unuse_way == 2'h1 ? _GEN_2806 : _GEN_8582; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9224 = unuse_way == 2'h1 ? _GEN_2807 : _GEN_8583; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9225 = unuse_way == 2'h1 ? _GEN_2808 : _GEN_8584; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9226 = unuse_way == 2'h1 ? _GEN_2809 : _GEN_8585; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9227 = unuse_way == 2'h1 ? _GEN_2810 : _GEN_8586; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9228 = unuse_way == 2'h1 ? _GEN_2811 : _GEN_8587; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9229 = unuse_way == 2'h1 ? _GEN_2812 : _GEN_8588; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9230 = unuse_way == 2'h1 ? _GEN_2813 : _GEN_8589; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9231 = unuse_way == 2'h1 ? _GEN_2814 : _GEN_8590; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9232 = unuse_way == 2'h1 ? _GEN_2815 : _GEN_8591; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9233 = unuse_way == 2'h1 ? _GEN_2816 : _GEN_8592; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9234 = unuse_way == 2'h1 ? _GEN_2817 : _GEN_8593; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9235 = unuse_way == 2'h1 ? _GEN_2818 : _GEN_8594; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9236 = unuse_way == 2'h1 ? _GEN_2819 : _GEN_8595; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9237 = unuse_way == 2'h1 ? _GEN_2820 : _GEN_8596; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9238 = unuse_way == 2'h1 ? _GEN_2821 : _GEN_8597; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9239 = unuse_way == 2'h1 ? _GEN_2822 : _GEN_8598; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9240 = unuse_way == 2'h1 ? _GEN_2823 : _GEN_8599; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9241 = unuse_way == 2'h1 ? _GEN_2824 : _GEN_8600; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9242 = unuse_way == 2'h1 ? _GEN_2825 : _GEN_8601; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9243 = unuse_way == 2'h1 ? _GEN_2826 : _GEN_8602; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9244 = unuse_way == 2'h1 ? _GEN_2827 : _GEN_8603; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9245 = unuse_way == 2'h1 ? _GEN_2828 : _GEN_8604; // @[d_cache.scala 134:34]
  wire [31:0] _GEN_9246 = unuse_way == 2'h1 ? _GEN_2829 : _GEN_8605; // @[d_cache.scala 134:34]
  wire  _GEN_9247 = unuse_way == 2'h1 ? _GEN_2830 : _GEN_8734; // @[d_cache.scala 134:34]
  wire  _GEN_9248 = unuse_way == 2'h1 ? _GEN_2831 : _GEN_8735; // @[d_cache.scala 134:34]
  wire  _GEN_9249 = unuse_way == 2'h1 ? _GEN_2832 : _GEN_8736; // @[d_cache.scala 134:34]
  wire  _GEN_9250 = unuse_way == 2'h1 ? _GEN_2833 : _GEN_8737; // @[d_cache.scala 134:34]
  wire  _GEN_9251 = unuse_way == 2'h1 ? _GEN_2834 : _GEN_8738; // @[d_cache.scala 134:34]
  wire  _GEN_9252 = unuse_way == 2'h1 ? _GEN_2835 : _GEN_8739; // @[d_cache.scala 134:34]
  wire  _GEN_9253 = unuse_way == 2'h1 ? _GEN_2836 : _GEN_8740; // @[d_cache.scala 134:34]
  wire  _GEN_9254 = unuse_way == 2'h1 ? _GEN_2837 : _GEN_8741; // @[d_cache.scala 134:34]
  wire  _GEN_9255 = unuse_way == 2'h1 ? _GEN_2838 : _GEN_8742; // @[d_cache.scala 134:34]
  wire  _GEN_9256 = unuse_way == 2'h1 ? _GEN_2839 : _GEN_8743; // @[d_cache.scala 134:34]
  wire  _GEN_9257 = unuse_way == 2'h1 ? _GEN_2840 : _GEN_8744; // @[d_cache.scala 134:34]
  wire  _GEN_9258 = unuse_way == 2'h1 ? _GEN_2841 : _GEN_8745; // @[d_cache.scala 134:34]
  wire  _GEN_9259 = unuse_way == 2'h1 ? _GEN_2842 : _GEN_8746; // @[d_cache.scala 134:34]
  wire  _GEN_9260 = unuse_way == 2'h1 ? _GEN_2843 : _GEN_8747; // @[d_cache.scala 134:34]
  wire  _GEN_9261 = unuse_way == 2'h1 ? _GEN_2844 : _GEN_8748; // @[d_cache.scala 134:34]
  wire  _GEN_9262 = unuse_way == 2'h1 ? _GEN_2845 : _GEN_8749; // @[d_cache.scala 134:34]
  wire  _GEN_9263 = unuse_way == 2'h1 ? _GEN_2846 : _GEN_8750; // @[d_cache.scala 134:34]
  wire  _GEN_9264 = unuse_way == 2'h1 ? _GEN_2847 : _GEN_8751; // @[d_cache.scala 134:34]
  wire  _GEN_9265 = unuse_way == 2'h1 ? _GEN_2848 : _GEN_8752; // @[d_cache.scala 134:34]
  wire  _GEN_9266 = unuse_way == 2'h1 ? _GEN_2849 : _GEN_8753; // @[d_cache.scala 134:34]
  wire  _GEN_9267 = unuse_way == 2'h1 ? _GEN_2850 : _GEN_8754; // @[d_cache.scala 134:34]
  wire  _GEN_9268 = unuse_way == 2'h1 ? _GEN_2851 : _GEN_8755; // @[d_cache.scala 134:34]
  wire  _GEN_9269 = unuse_way == 2'h1 ? _GEN_2852 : _GEN_8756; // @[d_cache.scala 134:34]
  wire  _GEN_9270 = unuse_way == 2'h1 ? _GEN_2853 : _GEN_8757; // @[d_cache.scala 134:34]
  wire  _GEN_9271 = unuse_way == 2'h1 ? _GEN_2854 : _GEN_8758; // @[d_cache.scala 134:34]
  wire  _GEN_9272 = unuse_way == 2'h1 ? _GEN_2855 : _GEN_8759; // @[d_cache.scala 134:34]
  wire  _GEN_9273 = unuse_way == 2'h1 ? _GEN_2856 : _GEN_8760; // @[d_cache.scala 134:34]
  wire  _GEN_9274 = unuse_way == 2'h1 ? _GEN_2857 : _GEN_8761; // @[d_cache.scala 134:34]
  wire  _GEN_9275 = unuse_way == 2'h1 ? _GEN_2858 : _GEN_8762; // @[d_cache.scala 134:34]
  wire  _GEN_9276 = unuse_way == 2'h1 ? _GEN_2859 : _GEN_8763; // @[d_cache.scala 134:34]
  wire  _GEN_9277 = unuse_way == 2'h1 ? _GEN_2860 : _GEN_8764; // @[d_cache.scala 134:34]
  wire  _GEN_9278 = unuse_way == 2'h1 ? _GEN_2861 : _GEN_8765; // @[d_cache.scala 134:34]
  wire  _GEN_9279 = unuse_way == 2'h1 ? _GEN_2862 : _GEN_8766; // @[d_cache.scala 134:34]
  wire  _GEN_9280 = unuse_way == 2'h1 ? _GEN_2863 : _GEN_8767; // @[d_cache.scala 134:34]
  wire  _GEN_9281 = unuse_way == 2'h1 ? _GEN_2864 : _GEN_8768; // @[d_cache.scala 134:34]
  wire  _GEN_9282 = unuse_way == 2'h1 ? _GEN_2865 : _GEN_8769; // @[d_cache.scala 134:34]
  wire  _GEN_9283 = unuse_way == 2'h1 ? _GEN_2866 : _GEN_8770; // @[d_cache.scala 134:34]
  wire  _GEN_9284 = unuse_way == 2'h1 ? _GEN_2867 : _GEN_8771; // @[d_cache.scala 134:34]
  wire  _GEN_9285 = unuse_way == 2'h1 ? _GEN_2868 : _GEN_8772; // @[d_cache.scala 134:34]
  wire  _GEN_9286 = unuse_way == 2'h1 ? _GEN_2869 : _GEN_8773; // @[d_cache.scala 134:34]
  wire  _GEN_9287 = unuse_way == 2'h1 ? _GEN_2870 : _GEN_8774; // @[d_cache.scala 134:34]
  wire  _GEN_9288 = unuse_way == 2'h1 ? _GEN_2871 : _GEN_8775; // @[d_cache.scala 134:34]
  wire  _GEN_9289 = unuse_way == 2'h1 ? _GEN_2872 : _GEN_8776; // @[d_cache.scala 134:34]
  wire  _GEN_9290 = unuse_way == 2'h1 ? _GEN_2873 : _GEN_8777; // @[d_cache.scala 134:34]
  wire  _GEN_9291 = unuse_way == 2'h1 ? _GEN_2874 : _GEN_8778; // @[d_cache.scala 134:34]
  wire  _GEN_9292 = unuse_way == 2'h1 ? _GEN_2875 : _GEN_8779; // @[d_cache.scala 134:34]
  wire  _GEN_9293 = unuse_way == 2'h1 ? _GEN_2876 : _GEN_8780; // @[d_cache.scala 134:34]
  wire  _GEN_9294 = unuse_way == 2'h1 ? _GEN_2877 : _GEN_8781; // @[d_cache.scala 134:34]
  wire  _GEN_9295 = unuse_way == 2'h1 ? _GEN_2878 : _GEN_8782; // @[d_cache.scala 134:34]
  wire  _GEN_9296 = unuse_way == 2'h1 ? _GEN_2879 : _GEN_8783; // @[d_cache.scala 134:34]
  wire  _GEN_9297 = unuse_way == 2'h1 ? _GEN_2880 : _GEN_8784; // @[d_cache.scala 134:34]
  wire  _GEN_9298 = unuse_way == 2'h1 ? _GEN_2881 : _GEN_8785; // @[d_cache.scala 134:34]
  wire  _GEN_9299 = unuse_way == 2'h1 ? _GEN_2882 : _GEN_8786; // @[d_cache.scala 134:34]
  wire  _GEN_9300 = unuse_way == 2'h1 ? _GEN_2883 : _GEN_8787; // @[d_cache.scala 134:34]
  wire  _GEN_9301 = unuse_way == 2'h1 ? _GEN_2884 : _GEN_8788; // @[d_cache.scala 134:34]
  wire  _GEN_9302 = unuse_way == 2'h1 ? _GEN_2885 : _GEN_8789; // @[d_cache.scala 134:34]
  wire  _GEN_9303 = unuse_way == 2'h1 ? _GEN_2886 : _GEN_8790; // @[d_cache.scala 134:34]
  wire  _GEN_9304 = unuse_way == 2'h1 ? _GEN_2887 : _GEN_8791; // @[d_cache.scala 134:34]
  wire  _GEN_9305 = unuse_way == 2'h1 ? _GEN_2888 : _GEN_8792; // @[d_cache.scala 134:34]
  wire  _GEN_9306 = unuse_way == 2'h1 ? _GEN_2889 : _GEN_8793; // @[d_cache.scala 134:34]
  wire  _GEN_9307 = unuse_way == 2'h1 ? _GEN_2890 : _GEN_8794; // @[d_cache.scala 134:34]
  wire  _GEN_9308 = unuse_way == 2'h1 ? _GEN_2891 : _GEN_8795; // @[d_cache.scala 134:34]
  wire  _GEN_9309 = unuse_way == 2'h1 ? _GEN_2892 : _GEN_8796; // @[d_cache.scala 134:34]
  wire  _GEN_9310 = unuse_way == 2'h1 ? _GEN_2893 : _GEN_8797; // @[d_cache.scala 134:34]
  wire  _GEN_9311 = unuse_way == 2'h1 ? _GEN_2894 : _GEN_8798; // @[d_cache.scala 134:34]
  wire  _GEN_9312 = unuse_way == 2'h1 ? _GEN_2895 : _GEN_8799; // @[d_cache.scala 134:34]
  wire  _GEN_9313 = unuse_way == 2'h1 ? _GEN_2896 : _GEN_8800; // @[d_cache.scala 134:34]
  wire  _GEN_9314 = unuse_way == 2'h1 ? _GEN_2897 : _GEN_8801; // @[d_cache.scala 134:34]
  wire  _GEN_9315 = unuse_way == 2'h1 ? _GEN_2898 : _GEN_8802; // @[d_cache.scala 134:34]
  wire  _GEN_9316 = unuse_way == 2'h1 ? _GEN_2899 : _GEN_8803; // @[d_cache.scala 134:34]
  wire  _GEN_9317 = unuse_way == 2'h1 ? _GEN_2900 : _GEN_8804; // @[d_cache.scala 134:34]
  wire  _GEN_9318 = unuse_way == 2'h1 ? _GEN_2901 : _GEN_8805; // @[d_cache.scala 134:34]
  wire  _GEN_9319 = unuse_way == 2'h1 ? _GEN_2902 : _GEN_8806; // @[d_cache.scala 134:34]
  wire  _GEN_9320 = unuse_way == 2'h1 ? _GEN_2903 : _GEN_8807; // @[d_cache.scala 134:34]
  wire  _GEN_9321 = unuse_way == 2'h1 ? _GEN_2904 : _GEN_8808; // @[d_cache.scala 134:34]
  wire  _GEN_9322 = unuse_way == 2'h1 ? _GEN_2905 : _GEN_8809; // @[d_cache.scala 134:34]
  wire  _GEN_9323 = unuse_way == 2'h1 ? _GEN_2906 : _GEN_8810; // @[d_cache.scala 134:34]
  wire  _GEN_9324 = unuse_way == 2'h1 ? _GEN_2907 : _GEN_8811; // @[d_cache.scala 134:34]
  wire  _GEN_9325 = unuse_way == 2'h1 ? _GEN_2908 : _GEN_8812; // @[d_cache.scala 134:34]
  wire  _GEN_9326 = unuse_way == 2'h1 ? _GEN_2909 : _GEN_8813; // @[d_cache.scala 134:34]
  wire  _GEN_9327 = unuse_way == 2'h1 ? _GEN_2910 : _GEN_8814; // @[d_cache.scala 134:34]
  wire  _GEN_9328 = unuse_way == 2'h1 ? _GEN_2911 : _GEN_8815; // @[d_cache.scala 134:34]
  wire  _GEN_9329 = unuse_way == 2'h1 ? _GEN_2912 : _GEN_8816; // @[d_cache.scala 134:34]
  wire  _GEN_9330 = unuse_way == 2'h1 ? _GEN_2913 : _GEN_8817; // @[d_cache.scala 134:34]
  wire  _GEN_9331 = unuse_way == 2'h1 ? _GEN_2914 : _GEN_8818; // @[d_cache.scala 134:34]
  wire  _GEN_9332 = unuse_way == 2'h1 ? _GEN_2915 : _GEN_8819; // @[d_cache.scala 134:34]
  wire  _GEN_9333 = unuse_way == 2'h1 ? _GEN_2916 : _GEN_8820; // @[d_cache.scala 134:34]
  wire  _GEN_9334 = unuse_way == 2'h1 ? _GEN_2917 : _GEN_8821; // @[d_cache.scala 134:34]
  wire  _GEN_9335 = unuse_way == 2'h1 ? _GEN_2918 : _GEN_8822; // @[d_cache.scala 134:34]
  wire  _GEN_9336 = unuse_way == 2'h1 ? _GEN_2919 : _GEN_8823; // @[d_cache.scala 134:34]
  wire  _GEN_9337 = unuse_way == 2'h1 ? _GEN_2920 : _GEN_8824; // @[d_cache.scala 134:34]
  wire  _GEN_9338 = unuse_way == 2'h1 ? _GEN_2921 : _GEN_8825; // @[d_cache.scala 134:34]
  wire  _GEN_9339 = unuse_way == 2'h1 ? _GEN_2922 : _GEN_8826; // @[d_cache.scala 134:34]
  wire  _GEN_9340 = unuse_way == 2'h1 ? _GEN_2923 : _GEN_8827; // @[d_cache.scala 134:34]
  wire  _GEN_9341 = unuse_way == 2'h1 ? _GEN_2924 : _GEN_8828; // @[d_cache.scala 134:34]
  wire  _GEN_9342 = unuse_way == 2'h1 ? _GEN_2925 : _GEN_8829; // @[d_cache.scala 134:34]
  wire  _GEN_9343 = unuse_way == 2'h1 ? _GEN_2926 : _GEN_8830; // @[d_cache.scala 134:34]
  wire  _GEN_9344 = unuse_way == 2'h1 ? _GEN_2927 : _GEN_8831; // @[d_cache.scala 134:34]
  wire  _GEN_9345 = unuse_way == 2'h1 ? _GEN_2928 : _GEN_8832; // @[d_cache.scala 134:34]
  wire  _GEN_9346 = unuse_way == 2'h1 ? _GEN_2929 : _GEN_8833; // @[d_cache.scala 134:34]
  wire  _GEN_9347 = unuse_way == 2'h1 ? _GEN_2930 : _GEN_8834; // @[d_cache.scala 134:34]
  wire  _GEN_9348 = unuse_way == 2'h1 ? _GEN_2931 : _GEN_8835; // @[d_cache.scala 134:34]
  wire  _GEN_9349 = unuse_way == 2'h1 ? _GEN_2932 : _GEN_8836; // @[d_cache.scala 134:34]
  wire  _GEN_9350 = unuse_way == 2'h1 ? _GEN_2933 : _GEN_8837; // @[d_cache.scala 134:34]
  wire  _GEN_9351 = unuse_way == 2'h1 ? _GEN_2934 : _GEN_8838; // @[d_cache.scala 134:34]
  wire  _GEN_9352 = unuse_way == 2'h1 ? _GEN_2935 : _GEN_8839; // @[d_cache.scala 134:34]
  wire  _GEN_9353 = unuse_way == 2'h1 ? _GEN_2936 : _GEN_8840; // @[d_cache.scala 134:34]
  wire  _GEN_9354 = unuse_way == 2'h1 ? _GEN_2937 : _GEN_8841; // @[d_cache.scala 134:34]
  wire  _GEN_9355 = unuse_way == 2'h1 ? _GEN_2938 : _GEN_8842; // @[d_cache.scala 134:34]
  wire  _GEN_9356 = unuse_way == 2'h1 ? _GEN_2939 : _GEN_8843; // @[d_cache.scala 134:34]
  wire  _GEN_9357 = unuse_way == 2'h1 ? _GEN_2940 : _GEN_8844; // @[d_cache.scala 134:34]
  wire  _GEN_9358 = unuse_way == 2'h1 ? _GEN_2941 : _GEN_8845; // @[d_cache.scala 134:34]
  wire  _GEN_9359 = unuse_way == 2'h1 ? _GEN_2942 : _GEN_8846; // @[d_cache.scala 134:34]
  wire  _GEN_9360 = unuse_way == 2'h1 ? _GEN_2943 : _GEN_8847; // @[d_cache.scala 134:34]
  wire  _GEN_9361 = unuse_way == 2'h1 ? _GEN_2944 : _GEN_8848; // @[d_cache.scala 134:34]
  wire  _GEN_9362 = unuse_way == 2'h1 ? _GEN_2945 : _GEN_8849; // @[d_cache.scala 134:34]
  wire  _GEN_9363 = unuse_way == 2'h1 ? _GEN_2946 : _GEN_8850; // @[d_cache.scala 134:34]
  wire  _GEN_9364 = unuse_way == 2'h1 ? _GEN_2947 : _GEN_8851; // @[d_cache.scala 134:34]
  wire  _GEN_9365 = unuse_way == 2'h1 ? _GEN_2948 : _GEN_8852; // @[d_cache.scala 134:34]
  wire  _GEN_9366 = unuse_way == 2'h1 ? _GEN_2949 : _GEN_8853; // @[d_cache.scala 134:34]
  wire  _GEN_9367 = unuse_way == 2'h1 ? _GEN_2950 : _GEN_8854; // @[d_cache.scala 134:34]
  wire  _GEN_9368 = unuse_way == 2'h1 ? _GEN_2951 : _GEN_8855; // @[d_cache.scala 134:34]
  wire  _GEN_9369 = unuse_way == 2'h1 ? _GEN_2952 : _GEN_8856; // @[d_cache.scala 134:34]
  wire  _GEN_9370 = unuse_way == 2'h1 ? _GEN_2953 : _GEN_8857; // @[d_cache.scala 134:34]
  wire  _GEN_9371 = unuse_way == 2'h1 ? _GEN_2954 : _GEN_8858; // @[d_cache.scala 134:34]
  wire  _GEN_9372 = unuse_way == 2'h1 ? _GEN_2955 : _GEN_8859; // @[d_cache.scala 134:34]
  wire  _GEN_9373 = unuse_way == 2'h1 ? _GEN_2956 : _GEN_8860; // @[d_cache.scala 134:34]
  wire  _GEN_9374 = unuse_way == 2'h1 ? _GEN_2957 : _GEN_8861; // @[d_cache.scala 134:34]
  wire  _GEN_9375 = unuse_way == 2'h1 | _GEN_8347; // @[d_cache.scala 134:34 139:23]
  wire [63:0] _GEN_9376 = unuse_way == 2'h1 ? ram_1_0 : _GEN_7963; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9377 = unuse_way == 2'h1 ? ram_1_1 : _GEN_7964; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9378 = unuse_way == 2'h1 ? ram_1_2 : _GEN_7965; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9379 = unuse_way == 2'h1 ? ram_1_3 : _GEN_7966; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9380 = unuse_way == 2'h1 ? ram_1_4 : _GEN_7967; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9381 = unuse_way == 2'h1 ? ram_1_5 : _GEN_7968; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9382 = unuse_way == 2'h1 ? ram_1_6 : _GEN_7969; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9383 = unuse_way == 2'h1 ? ram_1_7 : _GEN_7970; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9384 = unuse_way == 2'h1 ? ram_1_8 : _GEN_7971; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9385 = unuse_way == 2'h1 ? ram_1_9 : _GEN_7972; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9386 = unuse_way == 2'h1 ? ram_1_10 : _GEN_7973; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9387 = unuse_way == 2'h1 ? ram_1_11 : _GEN_7974; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9388 = unuse_way == 2'h1 ? ram_1_12 : _GEN_7975; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9389 = unuse_way == 2'h1 ? ram_1_13 : _GEN_7976; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9390 = unuse_way == 2'h1 ? ram_1_14 : _GEN_7977; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9391 = unuse_way == 2'h1 ? ram_1_15 : _GEN_7978; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9392 = unuse_way == 2'h1 ? ram_1_16 : _GEN_7979; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9393 = unuse_way == 2'h1 ? ram_1_17 : _GEN_7980; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9394 = unuse_way == 2'h1 ? ram_1_18 : _GEN_7981; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9395 = unuse_way == 2'h1 ? ram_1_19 : _GEN_7982; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9396 = unuse_way == 2'h1 ? ram_1_20 : _GEN_7983; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9397 = unuse_way == 2'h1 ? ram_1_21 : _GEN_7984; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9398 = unuse_way == 2'h1 ? ram_1_22 : _GEN_7985; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9399 = unuse_way == 2'h1 ? ram_1_23 : _GEN_7986; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9400 = unuse_way == 2'h1 ? ram_1_24 : _GEN_7987; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9401 = unuse_way == 2'h1 ? ram_1_25 : _GEN_7988; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9402 = unuse_way == 2'h1 ? ram_1_26 : _GEN_7989; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9403 = unuse_way == 2'h1 ? ram_1_27 : _GEN_7990; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9404 = unuse_way == 2'h1 ? ram_1_28 : _GEN_7991; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9405 = unuse_way == 2'h1 ? ram_1_29 : _GEN_7992; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9406 = unuse_way == 2'h1 ? ram_1_30 : _GEN_7993; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9407 = unuse_way == 2'h1 ? ram_1_31 : _GEN_7994; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9408 = unuse_way == 2'h1 ? ram_1_32 : _GEN_7995; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9409 = unuse_way == 2'h1 ? ram_1_33 : _GEN_7996; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9410 = unuse_way == 2'h1 ? ram_1_34 : _GEN_7997; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9411 = unuse_way == 2'h1 ? ram_1_35 : _GEN_7998; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9412 = unuse_way == 2'h1 ? ram_1_36 : _GEN_7999; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9413 = unuse_way == 2'h1 ? ram_1_37 : _GEN_8000; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9414 = unuse_way == 2'h1 ? ram_1_38 : _GEN_8001; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9415 = unuse_way == 2'h1 ? ram_1_39 : _GEN_8002; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9416 = unuse_way == 2'h1 ? ram_1_40 : _GEN_8003; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9417 = unuse_way == 2'h1 ? ram_1_41 : _GEN_8004; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9418 = unuse_way == 2'h1 ? ram_1_42 : _GEN_8005; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9419 = unuse_way == 2'h1 ? ram_1_43 : _GEN_8006; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9420 = unuse_way == 2'h1 ? ram_1_44 : _GEN_8007; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9421 = unuse_way == 2'h1 ? ram_1_45 : _GEN_8008; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9422 = unuse_way == 2'h1 ? ram_1_46 : _GEN_8009; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9423 = unuse_way == 2'h1 ? ram_1_47 : _GEN_8010; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9424 = unuse_way == 2'h1 ? ram_1_48 : _GEN_8011; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9425 = unuse_way == 2'h1 ? ram_1_49 : _GEN_8012; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9426 = unuse_way == 2'h1 ? ram_1_50 : _GEN_8013; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9427 = unuse_way == 2'h1 ? ram_1_51 : _GEN_8014; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9428 = unuse_way == 2'h1 ? ram_1_52 : _GEN_8015; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9429 = unuse_way == 2'h1 ? ram_1_53 : _GEN_8016; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9430 = unuse_way == 2'h1 ? ram_1_54 : _GEN_8017; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9431 = unuse_way == 2'h1 ? ram_1_55 : _GEN_8018; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9432 = unuse_way == 2'h1 ? ram_1_56 : _GEN_8019; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9433 = unuse_way == 2'h1 ? ram_1_57 : _GEN_8020; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9434 = unuse_way == 2'h1 ? ram_1_58 : _GEN_8021; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9435 = unuse_way == 2'h1 ? ram_1_59 : _GEN_8022; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9436 = unuse_way == 2'h1 ? ram_1_60 : _GEN_8023; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9437 = unuse_way == 2'h1 ? ram_1_61 : _GEN_8024; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9438 = unuse_way == 2'h1 ? ram_1_62 : _GEN_8025; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9439 = unuse_way == 2'h1 ? ram_1_63 : _GEN_8026; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9440 = unuse_way == 2'h1 ? ram_1_64 : _GEN_8027; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9441 = unuse_way == 2'h1 ? ram_1_65 : _GEN_8028; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9442 = unuse_way == 2'h1 ? ram_1_66 : _GEN_8029; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9443 = unuse_way == 2'h1 ? ram_1_67 : _GEN_8030; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9444 = unuse_way == 2'h1 ? ram_1_68 : _GEN_8031; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9445 = unuse_way == 2'h1 ? ram_1_69 : _GEN_8032; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9446 = unuse_way == 2'h1 ? ram_1_70 : _GEN_8033; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9447 = unuse_way == 2'h1 ? ram_1_71 : _GEN_8034; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9448 = unuse_way == 2'h1 ? ram_1_72 : _GEN_8035; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9449 = unuse_way == 2'h1 ? ram_1_73 : _GEN_8036; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9450 = unuse_way == 2'h1 ? ram_1_74 : _GEN_8037; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9451 = unuse_way == 2'h1 ? ram_1_75 : _GEN_8038; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9452 = unuse_way == 2'h1 ? ram_1_76 : _GEN_8039; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9453 = unuse_way == 2'h1 ? ram_1_77 : _GEN_8040; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9454 = unuse_way == 2'h1 ? ram_1_78 : _GEN_8041; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9455 = unuse_way == 2'h1 ? ram_1_79 : _GEN_8042; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9456 = unuse_way == 2'h1 ? ram_1_80 : _GEN_8043; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9457 = unuse_way == 2'h1 ? ram_1_81 : _GEN_8044; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9458 = unuse_way == 2'h1 ? ram_1_82 : _GEN_8045; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9459 = unuse_way == 2'h1 ? ram_1_83 : _GEN_8046; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9460 = unuse_way == 2'h1 ? ram_1_84 : _GEN_8047; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9461 = unuse_way == 2'h1 ? ram_1_85 : _GEN_8048; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9462 = unuse_way == 2'h1 ? ram_1_86 : _GEN_8049; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9463 = unuse_way == 2'h1 ? ram_1_87 : _GEN_8050; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9464 = unuse_way == 2'h1 ? ram_1_88 : _GEN_8051; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9465 = unuse_way == 2'h1 ? ram_1_89 : _GEN_8052; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9466 = unuse_way == 2'h1 ? ram_1_90 : _GEN_8053; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9467 = unuse_way == 2'h1 ? ram_1_91 : _GEN_8054; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9468 = unuse_way == 2'h1 ? ram_1_92 : _GEN_8055; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9469 = unuse_way == 2'h1 ? ram_1_93 : _GEN_8056; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9470 = unuse_way == 2'h1 ? ram_1_94 : _GEN_8057; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9471 = unuse_way == 2'h1 ? ram_1_95 : _GEN_8058; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9472 = unuse_way == 2'h1 ? ram_1_96 : _GEN_8059; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9473 = unuse_way == 2'h1 ? ram_1_97 : _GEN_8060; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9474 = unuse_way == 2'h1 ? ram_1_98 : _GEN_8061; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9475 = unuse_way == 2'h1 ? ram_1_99 : _GEN_8062; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9476 = unuse_way == 2'h1 ? ram_1_100 : _GEN_8063; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9477 = unuse_way == 2'h1 ? ram_1_101 : _GEN_8064; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9478 = unuse_way == 2'h1 ? ram_1_102 : _GEN_8065; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9479 = unuse_way == 2'h1 ? ram_1_103 : _GEN_8066; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9480 = unuse_way == 2'h1 ? ram_1_104 : _GEN_8067; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9481 = unuse_way == 2'h1 ? ram_1_105 : _GEN_8068; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9482 = unuse_way == 2'h1 ? ram_1_106 : _GEN_8069; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9483 = unuse_way == 2'h1 ? ram_1_107 : _GEN_8070; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9484 = unuse_way == 2'h1 ? ram_1_108 : _GEN_8071; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9485 = unuse_way == 2'h1 ? ram_1_109 : _GEN_8072; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9486 = unuse_way == 2'h1 ? ram_1_110 : _GEN_8073; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9487 = unuse_way == 2'h1 ? ram_1_111 : _GEN_8074; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9488 = unuse_way == 2'h1 ? ram_1_112 : _GEN_8075; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9489 = unuse_way == 2'h1 ? ram_1_113 : _GEN_8076; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9490 = unuse_way == 2'h1 ? ram_1_114 : _GEN_8077; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9491 = unuse_way == 2'h1 ? ram_1_115 : _GEN_8078; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9492 = unuse_way == 2'h1 ? ram_1_116 : _GEN_8079; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9493 = unuse_way == 2'h1 ? ram_1_117 : _GEN_8080; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9494 = unuse_way == 2'h1 ? ram_1_118 : _GEN_8081; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9495 = unuse_way == 2'h1 ? ram_1_119 : _GEN_8082; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9496 = unuse_way == 2'h1 ? ram_1_120 : _GEN_8083; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9497 = unuse_way == 2'h1 ? ram_1_121 : _GEN_8084; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9498 = unuse_way == 2'h1 ? ram_1_122 : _GEN_8085; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9499 = unuse_way == 2'h1 ? ram_1_123 : _GEN_8086; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9500 = unuse_way == 2'h1 ? ram_1_124 : _GEN_8087; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9501 = unuse_way == 2'h1 ? ram_1_125 : _GEN_8088; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9502 = unuse_way == 2'h1 ? ram_1_126 : _GEN_8089; // @[d_cache.scala 134:34 19:24]
  wire [63:0] _GEN_9503 = unuse_way == 2'h1 ? ram_1_127 : _GEN_8090; // @[d_cache.scala 134:34 19:24]
  wire [31:0] _GEN_9504 = unuse_way == 2'h1 ? tag_1_0 : _GEN_8091; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9505 = unuse_way == 2'h1 ? tag_1_1 : _GEN_8092; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9506 = unuse_way == 2'h1 ? tag_1_2 : _GEN_8093; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9507 = unuse_way == 2'h1 ? tag_1_3 : _GEN_8094; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9508 = unuse_way == 2'h1 ? tag_1_4 : _GEN_8095; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9509 = unuse_way == 2'h1 ? tag_1_5 : _GEN_8096; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9510 = unuse_way == 2'h1 ? tag_1_6 : _GEN_8097; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9511 = unuse_way == 2'h1 ? tag_1_7 : _GEN_8098; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9512 = unuse_way == 2'h1 ? tag_1_8 : _GEN_8099; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9513 = unuse_way == 2'h1 ? tag_1_9 : _GEN_8100; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9514 = unuse_way == 2'h1 ? tag_1_10 : _GEN_8101; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9515 = unuse_way == 2'h1 ? tag_1_11 : _GEN_8102; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9516 = unuse_way == 2'h1 ? tag_1_12 : _GEN_8103; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9517 = unuse_way == 2'h1 ? tag_1_13 : _GEN_8104; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9518 = unuse_way == 2'h1 ? tag_1_14 : _GEN_8105; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9519 = unuse_way == 2'h1 ? tag_1_15 : _GEN_8106; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9520 = unuse_way == 2'h1 ? tag_1_16 : _GEN_8107; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9521 = unuse_way == 2'h1 ? tag_1_17 : _GEN_8108; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9522 = unuse_way == 2'h1 ? tag_1_18 : _GEN_8109; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9523 = unuse_way == 2'h1 ? tag_1_19 : _GEN_8110; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9524 = unuse_way == 2'h1 ? tag_1_20 : _GEN_8111; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9525 = unuse_way == 2'h1 ? tag_1_21 : _GEN_8112; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9526 = unuse_way == 2'h1 ? tag_1_22 : _GEN_8113; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9527 = unuse_way == 2'h1 ? tag_1_23 : _GEN_8114; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9528 = unuse_way == 2'h1 ? tag_1_24 : _GEN_8115; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9529 = unuse_way == 2'h1 ? tag_1_25 : _GEN_8116; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9530 = unuse_way == 2'h1 ? tag_1_26 : _GEN_8117; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9531 = unuse_way == 2'h1 ? tag_1_27 : _GEN_8118; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9532 = unuse_way == 2'h1 ? tag_1_28 : _GEN_8119; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9533 = unuse_way == 2'h1 ? tag_1_29 : _GEN_8120; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9534 = unuse_way == 2'h1 ? tag_1_30 : _GEN_8121; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9535 = unuse_way == 2'h1 ? tag_1_31 : _GEN_8122; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9536 = unuse_way == 2'h1 ? tag_1_32 : _GEN_8123; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9537 = unuse_way == 2'h1 ? tag_1_33 : _GEN_8124; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9538 = unuse_way == 2'h1 ? tag_1_34 : _GEN_8125; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9539 = unuse_way == 2'h1 ? tag_1_35 : _GEN_8126; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9540 = unuse_way == 2'h1 ? tag_1_36 : _GEN_8127; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9541 = unuse_way == 2'h1 ? tag_1_37 : _GEN_8128; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9542 = unuse_way == 2'h1 ? tag_1_38 : _GEN_8129; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9543 = unuse_way == 2'h1 ? tag_1_39 : _GEN_8130; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9544 = unuse_way == 2'h1 ? tag_1_40 : _GEN_8131; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9545 = unuse_way == 2'h1 ? tag_1_41 : _GEN_8132; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9546 = unuse_way == 2'h1 ? tag_1_42 : _GEN_8133; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9547 = unuse_way == 2'h1 ? tag_1_43 : _GEN_8134; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9548 = unuse_way == 2'h1 ? tag_1_44 : _GEN_8135; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9549 = unuse_way == 2'h1 ? tag_1_45 : _GEN_8136; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9550 = unuse_way == 2'h1 ? tag_1_46 : _GEN_8137; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9551 = unuse_way == 2'h1 ? tag_1_47 : _GEN_8138; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9552 = unuse_way == 2'h1 ? tag_1_48 : _GEN_8139; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9553 = unuse_way == 2'h1 ? tag_1_49 : _GEN_8140; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9554 = unuse_way == 2'h1 ? tag_1_50 : _GEN_8141; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9555 = unuse_way == 2'h1 ? tag_1_51 : _GEN_8142; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9556 = unuse_way == 2'h1 ? tag_1_52 : _GEN_8143; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9557 = unuse_way == 2'h1 ? tag_1_53 : _GEN_8144; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9558 = unuse_way == 2'h1 ? tag_1_54 : _GEN_8145; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9559 = unuse_way == 2'h1 ? tag_1_55 : _GEN_8146; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9560 = unuse_way == 2'h1 ? tag_1_56 : _GEN_8147; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9561 = unuse_way == 2'h1 ? tag_1_57 : _GEN_8148; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9562 = unuse_way == 2'h1 ? tag_1_58 : _GEN_8149; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9563 = unuse_way == 2'h1 ? tag_1_59 : _GEN_8150; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9564 = unuse_way == 2'h1 ? tag_1_60 : _GEN_8151; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9565 = unuse_way == 2'h1 ? tag_1_61 : _GEN_8152; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9566 = unuse_way == 2'h1 ? tag_1_62 : _GEN_8153; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9567 = unuse_way == 2'h1 ? tag_1_63 : _GEN_8154; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9568 = unuse_way == 2'h1 ? tag_1_64 : _GEN_8155; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9569 = unuse_way == 2'h1 ? tag_1_65 : _GEN_8156; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9570 = unuse_way == 2'h1 ? tag_1_66 : _GEN_8157; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9571 = unuse_way == 2'h1 ? tag_1_67 : _GEN_8158; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9572 = unuse_way == 2'h1 ? tag_1_68 : _GEN_8159; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9573 = unuse_way == 2'h1 ? tag_1_69 : _GEN_8160; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9574 = unuse_way == 2'h1 ? tag_1_70 : _GEN_8161; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9575 = unuse_way == 2'h1 ? tag_1_71 : _GEN_8162; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9576 = unuse_way == 2'h1 ? tag_1_72 : _GEN_8163; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9577 = unuse_way == 2'h1 ? tag_1_73 : _GEN_8164; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9578 = unuse_way == 2'h1 ? tag_1_74 : _GEN_8165; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9579 = unuse_way == 2'h1 ? tag_1_75 : _GEN_8166; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9580 = unuse_way == 2'h1 ? tag_1_76 : _GEN_8167; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9581 = unuse_way == 2'h1 ? tag_1_77 : _GEN_8168; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9582 = unuse_way == 2'h1 ? tag_1_78 : _GEN_8169; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9583 = unuse_way == 2'h1 ? tag_1_79 : _GEN_8170; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9584 = unuse_way == 2'h1 ? tag_1_80 : _GEN_8171; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9585 = unuse_way == 2'h1 ? tag_1_81 : _GEN_8172; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9586 = unuse_way == 2'h1 ? tag_1_82 : _GEN_8173; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9587 = unuse_way == 2'h1 ? tag_1_83 : _GEN_8174; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9588 = unuse_way == 2'h1 ? tag_1_84 : _GEN_8175; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9589 = unuse_way == 2'h1 ? tag_1_85 : _GEN_8176; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9590 = unuse_way == 2'h1 ? tag_1_86 : _GEN_8177; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9591 = unuse_way == 2'h1 ? tag_1_87 : _GEN_8178; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9592 = unuse_way == 2'h1 ? tag_1_88 : _GEN_8179; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9593 = unuse_way == 2'h1 ? tag_1_89 : _GEN_8180; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9594 = unuse_way == 2'h1 ? tag_1_90 : _GEN_8181; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9595 = unuse_way == 2'h1 ? tag_1_91 : _GEN_8182; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9596 = unuse_way == 2'h1 ? tag_1_92 : _GEN_8183; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9597 = unuse_way == 2'h1 ? tag_1_93 : _GEN_8184; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9598 = unuse_way == 2'h1 ? tag_1_94 : _GEN_8185; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9599 = unuse_way == 2'h1 ? tag_1_95 : _GEN_8186; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9600 = unuse_way == 2'h1 ? tag_1_96 : _GEN_8187; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9601 = unuse_way == 2'h1 ? tag_1_97 : _GEN_8188; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9602 = unuse_way == 2'h1 ? tag_1_98 : _GEN_8189; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9603 = unuse_way == 2'h1 ? tag_1_99 : _GEN_8190; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9604 = unuse_way == 2'h1 ? tag_1_100 : _GEN_8191; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9605 = unuse_way == 2'h1 ? tag_1_101 : _GEN_8192; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9606 = unuse_way == 2'h1 ? tag_1_102 : _GEN_8193; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9607 = unuse_way == 2'h1 ? tag_1_103 : _GEN_8194; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9608 = unuse_way == 2'h1 ? tag_1_104 : _GEN_8195; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9609 = unuse_way == 2'h1 ? tag_1_105 : _GEN_8196; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9610 = unuse_way == 2'h1 ? tag_1_106 : _GEN_8197; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9611 = unuse_way == 2'h1 ? tag_1_107 : _GEN_8198; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9612 = unuse_way == 2'h1 ? tag_1_108 : _GEN_8199; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9613 = unuse_way == 2'h1 ? tag_1_109 : _GEN_8200; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9614 = unuse_way == 2'h1 ? tag_1_110 : _GEN_8201; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9615 = unuse_way == 2'h1 ? tag_1_111 : _GEN_8202; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9616 = unuse_way == 2'h1 ? tag_1_112 : _GEN_8203; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9617 = unuse_way == 2'h1 ? tag_1_113 : _GEN_8204; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9618 = unuse_way == 2'h1 ? tag_1_114 : _GEN_8205; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9619 = unuse_way == 2'h1 ? tag_1_115 : _GEN_8206; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9620 = unuse_way == 2'h1 ? tag_1_116 : _GEN_8207; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9621 = unuse_way == 2'h1 ? tag_1_117 : _GEN_8208; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9622 = unuse_way == 2'h1 ? tag_1_118 : _GEN_8209; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9623 = unuse_way == 2'h1 ? tag_1_119 : _GEN_8210; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9624 = unuse_way == 2'h1 ? tag_1_120 : _GEN_8211; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9625 = unuse_way == 2'h1 ? tag_1_121 : _GEN_8212; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9626 = unuse_way == 2'h1 ? tag_1_122 : _GEN_8213; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9627 = unuse_way == 2'h1 ? tag_1_123 : _GEN_8214; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9628 = unuse_way == 2'h1 ? tag_1_124 : _GEN_8215; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9629 = unuse_way == 2'h1 ? tag_1_125 : _GEN_8216; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9630 = unuse_way == 2'h1 ? tag_1_126 : _GEN_8217; // @[d_cache.scala 134:34 21:24]
  wire [31:0] _GEN_9631 = unuse_way == 2'h1 ? tag_1_127 : _GEN_8218; // @[d_cache.scala 134:34 21:24]
  wire  _GEN_9632 = unuse_way == 2'h1 ? valid_1_0 : _GEN_8219; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9633 = unuse_way == 2'h1 ? valid_1_1 : _GEN_8220; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9634 = unuse_way == 2'h1 ? valid_1_2 : _GEN_8221; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9635 = unuse_way == 2'h1 ? valid_1_3 : _GEN_8222; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9636 = unuse_way == 2'h1 ? valid_1_4 : _GEN_8223; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9637 = unuse_way == 2'h1 ? valid_1_5 : _GEN_8224; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9638 = unuse_way == 2'h1 ? valid_1_6 : _GEN_8225; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9639 = unuse_way == 2'h1 ? valid_1_7 : _GEN_8226; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9640 = unuse_way == 2'h1 ? valid_1_8 : _GEN_8227; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9641 = unuse_way == 2'h1 ? valid_1_9 : _GEN_8228; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9642 = unuse_way == 2'h1 ? valid_1_10 : _GEN_8229; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9643 = unuse_way == 2'h1 ? valid_1_11 : _GEN_8230; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9644 = unuse_way == 2'h1 ? valid_1_12 : _GEN_8231; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9645 = unuse_way == 2'h1 ? valid_1_13 : _GEN_8232; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9646 = unuse_way == 2'h1 ? valid_1_14 : _GEN_8233; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9647 = unuse_way == 2'h1 ? valid_1_15 : _GEN_8234; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9648 = unuse_way == 2'h1 ? valid_1_16 : _GEN_8235; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9649 = unuse_way == 2'h1 ? valid_1_17 : _GEN_8236; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9650 = unuse_way == 2'h1 ? valid_1_18 : _GEN_8237; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9651 = unuse_way == 2'h1 ? valid_1_19 : _GEN_8238; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9652 = unuse_way == 2'h1 ? valid_1_20 : _GEN_8239; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9653 = unuse_way == 2'h1 ? valid_1_21 : _GEN_8240; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9654 = unuse_way == 2'h1 ? valid_1_22 : _GEN_8241; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9655 = unuse_way == 2'h1 ? valid_1_23 : _GEN_8242; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9656 = unuse_way == 2'h1 ? valid_1_24 : _GEN_8243; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9657 = unuse_way == 2'h1 ? valid_1_25 : _GEN_8244; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9658 = unuse_way == 2'h1 ? valid_1_26 : _GEN_8245; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9659 = unuse_way == 2'h1 ? valid_1_27 : _GEN_8246; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9660 = unuse_way == 2'h1 ? valid_1_28 : _GEN_8247; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9661 = unuse_way == 2'h1 ? valid_1_29 : _GEN_8248; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9662 = unuse_way == 2'h1 ? valid_1_30 : _GEN_8249; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9663 = unuse_way == 2'h1 ? valid_1_31 : _GEN_8250; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9664 = unuse_way == 2'h1 ? valid_1_32 : _GEN_8251; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9665 = unuse_way == 2'h1 ? valid_1_33 : _GEN_8252; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9666 = unuse_way == 2'h1 ? valid_1_34 : _GEN_8253; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9667 = unuse_way == 2'h1 ? valid_1_35 : _GEN_8254; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9668 = unuse_way == 2'h1 ? valid_1_36 : _GEN_8255; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9669 = unuse_way == 2'h1 ? valid_1_37 : _GEN_8256; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9670 = unuse_way == 2'h1 ? valid_1_38 : _GEN_8257; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9671 = unuse_way == 2'h1 ? valid_1_39 : _GEN_8258; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9672 = unuse_way == 2'h1 ? valid_1_40 : _GEN_8259; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9673 = unuse_way == 2'h1 ? valid_1_41 : _GEN_8260; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9674 = unuse_way == 2'h1 ? valid_1_42 : _GEN_8261; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9675 = unuse_way == 2'h1 ? valid_1_43 : _GEN_8262; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9676 = unuse_way == 2'h1 ? valid_1_44 : _GEN_8263; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9677 = unuse_way == 2'h1 ? valid_1_45 : _GEN_8264; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9678 = unuse_way == 2'h1 ? valid_1_46 : _GEN_8265; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9679 = unuse_way == 2'h1 ? valid_1_47 : _GEN_8266; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9680 = unuse_way == 2'h1 ? valid_1_48 : _GEN_8267; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9681 = unuse_way == 2'h1 ? valid_1_49 : _GEN_8268; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9682 = unuse_way == 2'h1 ? valid_1_50 : _GEN_8269; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9683 = unuse_way == 2'h1 ? valid_1_51 : _GEN_8270; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9684 = unuse_way == 2'h1 ? valid_1_52 : _GEN_8271; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9685 = unuse_way == 2'h1 ? valid_1_53 : _GEN_8272; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9686 = unuse_way == 2'h1 ? valid_1_54 : _GEN_8273; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9687 = unuse_way == 2'h1 ? valid_1_55 : _GEN_8274; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9688 = unuse_way == 2'h1 ? valid_1_56 : _GEN_8275; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9689 = unuse_way == 2'h1 ? valid_1_57 : _GEN_8276; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9690 = unuse_way == 2'h1 ? valid_1_58 : _GEN_8277; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9691 = unuse_way == 2'h1 ? valid_1_59 : _GEN_8278; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9692 = unuse_way == 2'h1 ? valid_1_60 : _GEN_8279; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9693 = unuse_way == 2'h1 ? valid_1_61 : _GEN_8280; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9694 = unuse_way == 2'h1 ? valid_1_62 : _GEN_8281; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9695 = unuse_way == 2'h1 ? valid_1_63 : _GEN_8282; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9696 = unuse_way == 2'h1 ? valid_1_64 : _GEN_8283; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9697 = unuse_way == 2'h1 ? valid_1_65 : _GEN_8284; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9698 = unuse_way == 2'h1 ? valid_1_66 : _GEN_8285; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9699 = unuse_way == 2'h1 ? valid_1_67 : _GEN_8286; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9700 = unuse_way == 2'h1 ? valid_1_68 : _GEN_8287; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9701 = unuse_way == 2'h1 ? valid_1_69 : _GEN_8288; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9702 = unuse_way == 2'h1 ? valid_1_70 : _GEN_8289; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9703 = unuse_way == 2'h1 ? valid_1_71 : _GEN_8290; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9704 = unuse_way == 2'h1 ? valid_1_72 : _GEN_8291; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9705 = unuse_way == 2'h1 ? valid_1_73 : _GEN_8292; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9706 = unuse_way == 2'h1 ? valid_1_74 : _GEN_8293; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9707 = unuse_way == 2'h1 ? valid_1_75 : _GEN_8294; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9708 = unuse_way == 2'h1 ? valid_1_76 : _GEN_8295; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9709 = unuse_way == 2'h1 ? valid_1_77 : _GEN_8296; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9710 = unuse_way == 2'h1 ? valid_1_78 : _GEN_8297; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9711 = unuse_way == 2'h1 ? valid_1_79 : _GEN_8298; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9712 = unuse_way == 2'h1 ? valid_1_80 : _GEN_8299; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9713 = unuse_way == 2'h1 ? valid_1_81 : _GEN_8300; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9714 = unuse_way == 2'h1 ? valid_1_82 : _GEN_8301; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9715 = unuse_way == 2'h1 ? valid_1_83 : _GEN_8302; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9716 = unuse_way == 2'h1 ? valid_1_84 : _GEN_8303; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9717 = unuse_way == 2'h1 ? valid_1_85 : _GEN_8304; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9718 = unuse_way == 2'h1 ? valid_1_86 : _GEN_8305; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9719 = unuse_way == 2'h1 ? valid_1_87 : _GEN_8306; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9720 = unuse_way == 2'h1 ? valid_1_88 : _GEN_8307; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9721 = unuse_way == 2'h1 ? valid_1_89 : _GEN_8308; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9722 = unuse_way == 2'h1 ? valid_1_90 : _GEN_8309; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9723 = unuse_way == 2'h1 ? valid_1_91 : _GEN_8310; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9724 = unuse_way == 2'h1 ? valid_1_92 : _GEN_8311; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9725 = unuse_way == 2'h1 ? valid_1_93 : _GEN_8312; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9726 = unuse_way == 2'h1 ? valid_1_94 : _GEN_8313; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9727 = unuse_way == 2'h1 ? valid_1_95 : _GEN_8314; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9728 = unuse_way == 2'h1 ? valid_1_96 : _GEN_8315; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9729 = unuse_way == 2'h1 ? valid_1_97 : _GEN_8316; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9730 = unuse_way == 2'h1 ? valid_1_98 : _GEN_8317; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9731 = unuse_way == 2'h1 ? valid_1_99 : _GEN_8318; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9732 = unuse_way == 2'h1 ? valid_1_100 : _GEN_8319; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9733 = unuse_way == 2'h1 ? valid_1_101 : _GEN_8320; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9734 = unuse_way == 2'h1 ? valid_1_102 : _GEN_8321; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9735 = unuse_way == 2'h1 ? valid_1_103 : _GEN_8322; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9736 = unuse_way == 2'h1 ? valid_1_104 : _GEN_8323; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9737 = unuse_way == 2'h1 ? valid_1_105 : _GEN_8324; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9738 = unuse_way == 2'h1 ? valid_1_106 : _GEN_8325; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9739 = unuse_way == 2'h1 ? valid_1_107 : _GEN_8326; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9740 = unuse_way == 2'h1 ? valid_1_108 : _GEN_8327; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9741 = unuse_way == 2'h1 ? valid_1_109 : _GEN_8328; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9742 = unuse_way == 2'h1 ? valid_1_110 : _GEN_8329; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9743 = unuse_way == 2'h1 ? valid_1_111 : _GEN_8330; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9744 = unuse_way == 2'h1 ? valid_1_112 : _GEN_8331; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9745 = unuse_way == 2'h1 ? valid_1_113 : _GEN_8332; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9746 = unuse_way == 2'h1 ? valid_1_114 : _GEN_8333; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9747 = unuse_way == 2'h1 ? valid_1_115 : _GEN_8334; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9748 = unuse_way == 2'h1 ? valid_1_116 : _GEN_8335; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9749 = unuse_way == 2'h1 ? valid_1_117 : _GEN_8336; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9750 = unuse_way == 2'h1 ? valid_1_118 : _GEN_8337; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9751 = unuse_way == 2'h1 ? valid_1_119 : _GEN_8338; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9752 = unuse_way == 2'h1 ? valid_1_120 : _GEN_8339; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9753 = unuse_way == 2'h1 ? valid_1_121 : _GEN_8340; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9754 = unuse_way == 2'h1 ? valid_1_122 : _GEN_8341; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9755 = unuse_way == 2'h1 ? valid_1_123 : _GEN_8342; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9756 = unuse_way == 2'h1 ? valid_1_124 : _GEN_8343; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9757 = unuse_way == 2'h1 ? valid_1_125 : _GEN_8344; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9758 = unuse_way == 2'h1 ? valid_1_126 : _GEN_8345; // @[d_cache.scala 134:34 23:26]
  wire  _GEN_9759 = unuse_way == 2'h1 ? valid_1_127 : _GEN_8346; // @[d_cache.scala 134:34 23:26]
  wire [63:0] _GEN_9760 = unuse_way == 2'h1 ? write_back_data : _GEN_8348; // @[d_cache.scala 134:34 29:34]
  wire [41:0] _GEN_9761 = unuse_way == 2'h1 ? {{10'd0}, write_back_addr} : _GEN_8349; // @[d_cache.scala 134:34 30:34]
  wire  _GEN_9762 = unuse_way == 2'h1 ? dirty_0_0 : _GEN_8606; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9763 = unuse_way == 2'h1 ? dirty_0_1 : _GEN_8607; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9764 = unuse_way == 2'h1 ? dirty_0_2 : _GEN_8608; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9765 = unuse_way == 2'h1 ? dirty_0_3 : _GEN_8609; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9766 = unuse_way == 2'h1 ? dirty_0_4 : _GEN_8610; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9767 = unuse_way == 2'h1 ? dirty_0_5 : _GEN_8611; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9768 = unuse_way == 2'h1 ? dirty_0_6 : _GEN_8612; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9769 = unuse_way == 2'h1 ? dirty_0_7 : _GEN_8613; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9770 = unuse_way == 2'h1 ? dirty_0_8 : _GEN_8614; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9771 = unuse_way == 2'h1 ? dirty_0_9 : _GEN_8615; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9772 = unuse_way == 2'h1 ? dirty_0_10 : _GEN_8616; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9773 = unuse_way == 2'h1 ? dirty_0_11 : _GEN_8617; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9774 = unuse_way == 2'h1 ? dirty_0_12 : _GEN_8618; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9775 = unuse_way == 2'h1 ? dirty_0_13 : _GEN_8619; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9776 = unuse_way == 2'h1 ? dirty_0_14 : _GEN_8620; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9777 = unuse_way == 2'h1 ? dirty_0_15 : _GEN_8621; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9778 = unuse_way == 2'h1 ? dirty_0_16 : _GEN_8622; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9779 = unuse_way == 2'h1 ? dirty_0_17 : _GEN_8623; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9780 = unuse_way == 2'h1 ? dirty_0_18 : _GEN_8624; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9781 = unuse_way == 2'h1 ? dirty_0_19 : _GEN_8625; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9782 = unuse_way == 2'h1 ? dirty_0_20 : _GEN_8626; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9783 = unuse_way == 2'h1 ? dirty_0_21 : _GEN_8627; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9784 = unuse_way == 2'h1 ? dirty_0_22 : _GEN_8628; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9785 = unuse_way == 2'h1 ? dirty_0_23 : _GEN_8629; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9786 = unuse_way == 2'h1 ? dirty_0_24 : _GEN_8630; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9787 = unuse_way == 2'h1 ? dirty_0_25 : _GEN_8631; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9788 = unuse_way == 2'h1 ? dirty_0_26 : _GEN_8632; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9789 = unuse_way == 2'h1 ? dirty_0_27 : _GEN_8633; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9790 = unuse_way == 2'h1 ? dirty_0_28 : _GEN_8634; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9791 = unuse_way == 2'h1 ? dirty_0_29 : _GEN_8635; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9792 = unuse_way == 2'h1 ? dirty_0_30 : _GEN_8636; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9793 = unuse_way == 2'h1 ? dirty_0_31 : _GEN_8637; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9794 = unuse_way == 2'h1 ? dirty_0_32 : _GEN_8638; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9795 = unuse_way == 2'h1 ? dirty_0_33 : _GEN_8639; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9796 = unuse_way == 2'h1 ? dirty_0_34 : _GEN_8640; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9797 = unuse_way == 2'h1 ? dirty_0_35 : _GEN_8641; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9798 = unuse_way == 2'h1 ? dirty_0_36 : _GEN_8642; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9799 = unuse_way == 2'h1 ? dirty_0_37 : _GEN_8643; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9800 = unuse_way == 2'h1 ? dirty_0_38 : _GEN_8644; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9801 = unuse_way == 2'h1 ? dirty_0_39 : _GEN_8645; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9802 = unuse_way == 2'h1 ? dirty_0_40 : _GEN_8646; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9803 = unuse_way == 2'h1 ? dirty_0_41 : _GEN_8647; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9804 = unuse_way == 2'h1 ? dirty_0_42 : _GEN_8648; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9805 = unuse_way == 2'h1 ? dirty_0_43 : _GEN_8649; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9806 = unuse_way == 2'h1 ? dirty_0_44 : _GEN_8650; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9807 = unuse_way == 2'h1 ? dirty_0_45 : _GEN_8651; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9808 = unuse_way == 2'h1 ? dirty_0_46 : _GEN_8652; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9809 = unuse_way == 2'h1 ? dirty_0_47 : _GEN_8653; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9810 = unuse_way == 2'h1 ? dirty_0_48 : _GEN_8654; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9811 = unuse_way == 2'h1 ? dirty_0_49 : _GEN_8655; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9812 = unuse_way == 2'h1 ? dirty_0_50 : _GEN_8656; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9813 = unuse_way == 2'h1 ? dirty_0_51 : _GEN_8657; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9814 = unuse_way == 2'h1 ? dirty_0_52 : _GEN_8658; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9815 = unuse_way == 2'h1 ? dirty_0_53 : _GEN_8659; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9816 = unuse_way == 2'h1 ? dirty_0_54 : _GEN_8660; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9817 = unuse_way == 2'h1 ? dirty_0_55 : _GEN_8661; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9818 = unuse_way == 2'h1 ? dirty_0_56 : _GEN_8662; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9819 = unuse_way == 2'h1 ? dirty_0_57 : _GEN_8663; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9820 = unuse_way == 2'h1 ? dirty_0_58 : _GEN_8664; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9821 = unuse_way == 2'h1 ? dirty_0_59 : _GEN_8665; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9822 = unuse_way == 2'h1 ? dirty_0_60 : _GEN_8666; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9823 = unuse_way == 2'h1 ? dirty_0_61 : _GEN_8667; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9824 = unuse_way == 2'h1 ? dirty_0_62 : _GEN_8668; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9825 = unuse_way == 2'h1 ? dirty_0_63 : _GEN_8669; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9826 = unuse_way == 2'h1 ? dirty_0_64 : _GEN_8670; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9827 = unuse_way == 2'h1 ? dirty_0_65 : _GEN_8671; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9828 = unuse_way == 2'h1 ? dirty_0_66 : _GEN_8672; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9829 = unuse_way == 2'h1 ? dirty_0_67 : _GEN_8673; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9830 = unuse_way == 2'h1 ? dirty_0_68 : _GEN_8674; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9831 = unuse_way == 2'h1 ? dirty_0_69 : _GEN_8675; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9832 = unuse_way == 2'h1 ? dirty_0_70 : _GEN_8676; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9833 = unuse_way == 2'h1 ? dirty_0_71 : _GEN_8677; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9834 = unuse_way == 2'h1 ? dirty_0_72 : _GEN_8678; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9835 = unuse_way == 2'h1 ? dirty_0_73 : _GEN_8679; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9836 = unuse_way == 2'h1 ? dirty_0_74 : _GEN_8680; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9837 = unuse_way == 2'h1 ? dirty_0_75 : _GEN_8681; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9838 = unuse_way == 2'h1 ? dirty_0_76 : _GEN_8682; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9839 = unuse_way == 2'h1 ? dirty_0_77 : _GEN_8683; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9840 = unuse_way == 2'h1 ? dirty_0_78 : _GEN_8684; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9841 = unuse_way == 2'h1 ? dirty_0_79 : _GEN_8685; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9842 = unuse_way == 2'h1 ? dirty_0_80 : _GEN_8686; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9843 = unuse_way == 2'h1 ? dirty_0_81 : _GEN_8687; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9844 = unuse_way == 2'h1 ? dirty_0_82 : _GEN_8688; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9845 = unuse_way == 2'h1 ? dirty_0_83 : _GEN_8689; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9846 = unuse_way == 2'h1 ? dirty_0_84 : _GEN_8690; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9847 = unuse_way == 2'h1 ? dirty_0_85 : _GEN_8691; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9848 = unuse_way == 2'h1 ? dirty_0_86 : _GEN_8692; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9849 = unuse_way == 2'h1 ? dirty_0_87 : _GEN_8693; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9850 = unuse_way == 2'h1 ? dirty_0_88 : _GEN_8694; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9851 = unuse_way == 2'h1 ? dirty_0_89 : _GEN_8695; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9852 = unuse_way == 2'h1 ? dirty_0_90 : _GEN_8696; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9853 = unuse_way == 2'h1 ? dirty_0_91 : _GEN_8697; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9854 = unuse_way == 2'h1 ? dirty_0_92 : _GEN_8698; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9855 = unuse_way == 2'h1 ? dirty_0_93 : _GEN_8699; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9856 = unuse_way == 2'h1 ? dirty_0_94 : _GEN_8700; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9857 = unuse_way == 2'h1 ? dirty_0_95 : _GEN_8701; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9858 = unuse_way == 2'h1 ? dirty_0_96 : _GEN_8702; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9859 = unuse_way == 2'h1 ? dirty_0_97 : _GEN_8703; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9860 = unuse_way == 2'h1 ? dirty_0_98 : _GEN_8704; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9861 = unuse_way == 2'h1 ? dirty_0_99 : _GEN_8705; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9862 = unuse_way == 2'h1 ? dirty_0_100 : _GEN_8706; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9863 = unuse_way == 2'h1 ? dirty_0_101 : _GEN_8707; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9864 = unuse_way == 2'h1 ? dirty_0_102 : _GEN_8708; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9865 = unuse_way == 2'h1 ? dirty_0_103 : _GEN_8709; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9866 = unuse_way == 2'h1 ? dirty_0_104 : _GEN_8710; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9867 = unuse_way == 2'h1 ? dirty_0_105 : _GEN_8711; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9868 = unuse_way == 2'h1 ? dirty_0_106 : _GEN_8712; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9869 = unuse_way == 2'h1 ? dirty_0_107 : _GEN_8713; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9870 = unuse_way == 2'h1 ? dirty_0_108 : _GEN_8714; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9871 = unuse_way == 2'h1 ? dirty_0_109 : _GEN_8715; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9872 = unuse_way == 2'h1 ? dirty_0_110 : _GEN_8716; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9873 = unuse_way == 2'h1 ? dirty_0_111 : _GEN_8717; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9874 = unuse_way == 2'h1 ? dirty_0_112 : _GEN_8718; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9875 = unuse_way == 2'h1 ? dirty_0_113 : _GEN_8719; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9876 = unuse_way == 2'h1 ? dirty_0_114 : _GEN_8720; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9877 = unuse_way == 2'h1 ? dirty_0_115 : _GEN_8721; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9878 = unuse_way == 2'h1 ? dirty_0_116 : _GEN_8722; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9879 = unuse_way == 2'h1 ? dirty_0_117 : _GEN_8723; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9880 = unuse_way == 2'h1 ? dirty_0_118 : _GEN_8724; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9881 = unuse_way == 2'h1 ? dirty_0_119 : _GEN_8725; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9882 = unuse_way == 2'h1 ? dirty_0_120 : _GEN_8726; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9883 = unuse_way == 2'h1 ? dirty_0_121 : _GEN_8727; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9884 = unuse_way == 2'h1 ? dirty_0_122 : _GEN_8728; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9885 = unuse_way == 2'h1 ? dirty_0_123 : _GEN_8729; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9886 = unuse_way == 2'h1 ? dirty_0_124 : _GEN_8730; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9887 = unuse_way == 2'h1 ? dirty_0_125 : _GEN_8731; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9888 = unuse_way == 2'h1 ? dirty_0_126 : _GEN_8732; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9889 = unuse_way == 2'h1 ? dirty_0_127 : _GEN_8733; // @[d_cache.scala 134:34 24:26]
  wire  _GEN_9890 = unuse_way == 2'h1 ? dirty_1_0 : _GEN_8862; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9891 = unuse_way == 2'h1 ? dirty_1_1 : _GEN_8863; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9892 = unuse_way == 2'h1 ? dirty_1_2 : _GEN_8864; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9893 = unuse_way == 2'h1 ? dirty_1_3 : _GEN_8865; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9894 = unuse_way == 2'h1 ? dirty_1_4 : _GEN_8866; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9895 = unuse_way == 2'h1 ? dirty_1_5 : _GEN_8867; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9896 = unuse_way == 2'h1 ? dirty_1_6 : _GEN_8868; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9897 = unuse_way == 2'h1 ? dirty_1_7 : _GEN_8869; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9898 = unuse_way == 2'h1 ? dirty_1_8 : _GEN_8870; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9899 = unuse_way == 2'h1 ? dirty_1_9 : _GEN_8871; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9900 = unuse_way == 2'h1 ? dirty_1_10 : _GEN_8872; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9901 = unuse_way == 2'h1 ? dirty_1_11 : _GEN_8873; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9902 = unuse_way == 2'h1 ? dirty_1_12 : _GEN_8874; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9903 = unuse_way == 2'h1 ? dirty_1_13 : _GEN_8875; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9904 = unuse_way == 2'h1 ? dirty_1_14 : _GEN_8876; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9905 = unuse_way == 2'h1 ? dirty_1_15 : _GEN_8877; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9906 = unuse_way == 2'h1 ? dirty_1_16 : _GEN_8878; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9907 = unuse_way == 2'h1 ? dirty_1_17 : _GEN_8879; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9908 = unuse_way == 2'h1 ? dirty_1_18 : _GEN_8880; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9909 = unuse_way == 2'h1 ? dirty_1_19 : _GEN_8881; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9910 = unuse_way == 2'h1 ? dirty_1_20 : _GEN_8882; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9911 = unuse_way == 2'h1 ? dirty_1_21 : _GEN_8883; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9912 = unuse_way == 2'h1 ? dirty_1_22 : _GEN_8884; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9913 = unuse_way == 2'h1 ? dirty_1_23 : _GEN_8885; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9914 = unuse_way == 2'h1 ? dirty_1_24 : _GEN_8886; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9915 = unuse_way == 2'h1 ? dirty_1_25 : _GEN_8887; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9916 = unuse_way == 2'h1 ? dirty_1_26 : _GEN_8888; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9917 = unuse_way == 2'h1 ? dirty_1_27 : _GEN_8889; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9918 = unuse_way == 2'h1 ? dirty_1_28 : _GEN_8890; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9919 = unuse_way == 2'h1 ? dirty_1_29 : _GEN_8891; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9920 = unuse_way == 2'h1 ? dirty_1_30 : _GEN_8892; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9921 = unuse_way == 2'h1 ? dirty_1_31 : _GEN_8893; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9922 = unuse_way == 2'h1 ? dirty_1_32 : _GEN_8894; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9923 = unuse_way == 2'h1 ? dirty_1_33 : _GEN_8895; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9924 = unuse_way == 2'h1 ? dirty_1_34 : _GEN_8896; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9925 = unuse_way == 2'h1 ? dirty_1_35 : _GEN_8897; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9926 = unuse_way == 2'h1 ? dirty_1_36 : _GEN_8898; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9927 = unuse_way == 2'h1 ? dirty_1_37 : _GEN_8899; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9928 = unuse_way == 2'h1 ? dirty_1_38 : _GEN_8900; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9929 = unuse_way == 2'h1 ? dirty_1_39 : _GEN_8901; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9930 = unuse_way == 2'h1 ? dirty_1_40 : _GEN_8902; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9931 = unuse_way == 2'h1 ? dirty_1_41 : _GEN_8903; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9932 = unuse_way == 2'h1 ? dirty_1_42 : _GEN_8904; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9933 = unuse_way == 2'h1 ? dirty_1_43 : _GEN_8905; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9934 = unuse_way == 2'h1 ? dirty_1_44 : _GEN_8906; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9935 = unuse_way == 2'h1 ? dirty_1_45 : _GEN_8907; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9936 = unuse_way == 2'h1 ? dirty_1_46 : _GEN_8908; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9937 = unuse_way == 2'h1 ? dirty_1_47 : _GEN_8909; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9938 = unuse_way == 2'h1 ? dirty_1_48 : _GEN_8910; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9939 = unuse_way == 2'h1 ? dirty_1_49 : _GEN_8911; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9940 = unuse_way == 2'h1 ? dirty_1_50 : _GEN_8912; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9941 = unuse_way == 2'h1 ? dirty_1_51 : _GEN_8913; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9942 = unuse_way == 2'h1 ? dirty_1_52 : _GEN_8914; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9943 = unuse_way == 2'h1 ? dirty_1_53 : _GEN_8915; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9944 = unuse_way == 2'h1 ? dirty_1_54 : _GEN_8916; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9945 = unuse_way == 2'h1 ? dirty_1_55 : _GEN_8917; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9946 = unuse_way == 2'h1 ? dirty_1_56 : _GEN_8918; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9947 = unuse_way == 2'h1 ? dirty_1_57 : _GEN_8919; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9948 = unuse_way == 2'h1 ? dirty_1_58 : _GEN_8920; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9949 = unuse_way == 2'h1 ? dirty_1_59 : _GEN_8921; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9950 = unuse_way == 2'h1 ? dirty_1_60 : _GEN_8922; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9951 = unuse_way == 2'h1 ? dirty_1_61 : _GEN_8923; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9952 = unuse_way == 2'h1 ? dirty_1_62 : _GEN_8924; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9953 = unuse_way == 2'h1 ? dirty_1_63 : _GEN_8925; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9954 = unuse_way == 2'h1 ? dirty_1_64 : _GEN_8926; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9955 = unuse_way == 2'h1 ? dirty_1_65 : _GEN_8927; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9956 = unuse_way == 2'h1 ? dirty_1_66 : _GEN_8928; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9957 = unuse_way == 2'h1 ? dirty_1_67 : _GEN_8929; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9958 = unuse_way == 2'h1 ? dirty_1_68 : _GEN_8930; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9959 = unuse_way == 2'h1 ? dirty_1_69 : _GEN_8931; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9960 = unuse_way == 2'h1 ? dirty_1_70 : _GEN_8932; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9961 = unuse_way == 2'h1 ? dirty_1_71 : _GEN_8933; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9962 = unuse_way == 2'h1 ? dirty_1_72 : _GEN_8934; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9963 = unuse_way == 2'h1 ? dirty_1_73 : _GEN_8935; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9964 = unuse_way == 2'h1 ? dirty_1_74 : _GEN_8936; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9965 = unuse_way == 2'h1 ? dirty_1_75 : _GEN_8937; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9966 = unuse_way == 2'h1 ? dirty_1_76 : _GEN_8938; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9967 = unuse_way == 2'h1 ? dirty_1_77 : _GEN_8939; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9968 = unuse_way == 2'h1 ? dirty_1_78 : _GEN_8940; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9969 = unuse_way == 2'h1 ? dirty_1_79 : _GEN_8941; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9970 = unuse_way == 2'h1 ? dirty_1_80 : _GEN_8942; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9971 = unuse_way == 2'h1 ? dirty_1_81 : _GEN_8943; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9972 = unuse_way == 2'h1 ? dirty_1_82 : _GEN_8944; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9973 = unuse_way == 2'h1 ? dirty_1_83 : _GEN_8945; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9974 = unuse_way == 2'h1 ? dirty_1_84 : _GEN_8946; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9975 = unuse_way == 2'h1 ? dirty_1_85 : _GEN_8947; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9976 = unuse_way == 2'h1 ? dirty_1_86 : _GEN_8948; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9977 = unuse_way == 2'h1 ? dirty_1_87 : _GEN_8949; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9978 = unuse_way == 2'h1 ? dirty_1_88 : _GEN_8950; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9979 = unuse_way == 2'h1 ? dirty_1_89 : _GEN_8951; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9980 = unuse_way == 2'h1 ? dirty_1_90 : _GEN_8952; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9981 = unuse_way == 2'h1 ? dirty_1_91 : _GEN_8953; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9982 = unuse_way == 2'h1 ? dirty_1_92 : _GEN_8954; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9983 = unuse_way == 2'h1 ? dirty_1_93 : _GEN_8955; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9984 = unuse_way == 2'h1 ? dirty_1_94 : _GEN_8956; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9985 = unuse_way == 2'h1 ? dirty_1_95 : _GEN_8957; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9986 = unuse_way == 2'h1 ? dirty_1_96 : _GEN_8958; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9987 = unuse_way == 2'h1 ? dirty_1_97 : _GEN_8959; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9988 = unuse_way == 2'h1 ? dirty_1_98 : _GEN_8960; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9989 = unuse_way == 2'h1 ? dirty_1_99 : _GEN_8961; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9990 = unuse_way == 2'h1 ? dirty_1_100 : _GEN_8962; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9991 = unuse_way == 2'h1 ? dirty_1_101 : _GEN_8963; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9992 = unuse_way == 2'h1 ? dirty_1_102 : _GEN_8964; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9993 = unuse_way == 2'h1 ? dirty_1_103 : _GEN_8965; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9994 = unuse_way == 2'h1 ? dirty_1_104 : _GEN_8966; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9995 = unuse_way == 2'h1 ? dirty_1_105 : _GEN_8967; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9996 = unuse_way == 2'h1 ? dirty_1_106 : _GEN_8968; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9997 = unuse_way == 2'h1 ? dirty_1_107 : _GEN_8969; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9998 = unuse_way == 2'h1 ? dirty_1_108 : _GEN_8970; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_9999 = unuse_way == 2'h1 ? dirty_1_109 : _GEN_8971; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10000 = unuse_way == 2'h1 ? dirty_1_110 : _GEN_8972; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10001 = unuse_way == 2'h1 ? dirty_1_111 : _GEN_8973; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10002 = unuse_way == 2'h1 ? dirty_1_112 : _GEN_8974; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10003 = unuse_way == 2'h1 ? dirty_1_113 : _GEN_8975; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10004 = unuse_way == 2'h1 ? dirty_1_114 : _GEN_8976; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10005 = unuse_way == 2'h1 ? dirty_1_115 : _GEN_8977; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10006 = unuse_way == 2'h1 ? dirty_1_116 : _GEN_8978; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10007 = unuse_way == 2'h1 ? dirty_1_117 : _GEN_8979; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10008 = unuse_way == 2'h1 ? dirty_1_118 : _GEN_8980; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10009 = unuse_way == 2'h1 ? dirty_1_119 : _GEN_8981; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10010 = unuse_way == 2'h1 ? dirty_1_120 : _GEN_8982; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10011 = unuse_way == 2'h1 ? dirty_1_121 : _GEN_8983; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10012 = unuse_way == 2'h1 ? dirty_1_122 : _GEN_8984; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10013 = unuse_way == 2'h1 ? dirty_1_123 : _GEN_8985; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10014 = unuse_way == 2'h1 ? dirty_1_124 : _GEN_8986; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10015 = unuse_way == 2'h1 ? dirty_1_125 : _GEN_8987; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10016 = unuse_way == 2'h1 ? dirty_1_126 : _GEN_8988; // @[d_cache.scala 134:34 25:26]
  wire  _GEN_10017 = unuse_way == 2'h1 ? dirty_1_127 : _GEN_8989; // @[d_cache.scala 134:34 25:26]
  wire [2:0] _GEN_10018 = io_from_axi_bvalid ? 3'h5 : state; // @[d_cache.scala 186:37 187:23 73:24]
  wire [2:0] _GEN_10019 = 3'h7 == state ? 3'h1 : state; // @[d_cache.scala 78:18 191:19 73:24]
  wire [2:0] _GEN_10020 = 3'h6 == state ? _GEN_10018 : _GEN_10019; // @[d_cache.scala 78:18]
  wire [2:0] _GEN_10021 = 3'h5 == state ? _GEN_8990 : _GEN_10020; // @[d_cache.scala 78:18]
  wire [63:0] _GEN_10022 = 3'h5 == state ? _GEN_8991 : ram_0_0; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10023 = 3'h5 == state ? _GEN_8992 : ram_0_1; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10024 = 3'h5 == state ? _GEN_8993 : ram_0_2; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10025 = 3'h5 == state ? _GEN_8994 : ram_0_3; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10026 = 3'h5 == state ? _GEN_8995 : ram_0_4; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10027 = 3'h5 == state ? _GEN_8996 : ram_0_5; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10028 = 3'h5 == state ? _GEN_8997 : ram_0_6; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10029 = 3'h5 == state ? _GEN_8998 : ram_0_7; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10030 = 3'h5 == state ? _GEN_8999 : ram_0_8; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10031 = 3'h5 == state ? _GEN_9000 : ram_0_9; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10032 = 3'h5 == state ? _GEN_9001 : ram_0_10; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10033 = 3'h5 == state ? _GEN_9002 : ram_0_11; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10034 = 3'h5 == state ? _GEN_9003 : ram_0_12; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10035 = 3'h5 == state ? _GEN_9004 : ram_0_13; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10036 = 3'h5 == state ? _GEN_9005 : ram_0_14; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10037 = 3'h5 == state ? _GEN_9006 : ram_0_15; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10038 = 3'h5 == state ? _GEN_9007 : ram_0_16; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10039 = 3'h5 == state ? _GEN_9008 : ram_0_17; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10040 = 3'h5 == state ? _GEN_9009 : ram_0_18; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10041 = 3'h5 == state ? _GEN_9010 : ram_0_19; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10042 = 3'h5 == state ? _GEN_9011 : ram_0_20; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10043 = 3'h5 == state ? _GEN_9012 : ram_0_21; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10044 = 3'h5 == state ? _GEN_9013 : ram_0_22; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10045 = 3'h5 == state ? _GEN_9014 : ram_0_23; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10046 = 3'h5 == state ? _GEN_9015 : ram_0_24; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10047 = 3'h5 == state ? _GEN_9016 : ram_0_25; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10048 = 3'h5 == state ? _GEN_9017 : ram_0_26; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10049 = 3'h5 == state ? _GEN_9018 : ram_0_27; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10050 = 3'h5 == state ? _GEN_9019 : ram_0_28; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10051 = 3'h5 == state ? _GEN_9020 : ram_0_29; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10052 = 3'h5 == state ? _GEN_9021 : ram_0_30; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10053 = 3'h5 == state ? _GEN_9022 : ram_0_31; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10054 = 3'h5 == state ? _GEN_9023 : ram_0_32; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10055 = 3'h5 == state ? _GEN_9024 : ram_0_33; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10056 = 3'h5 == state ? _GEN_9025 : ram_0_34; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10057 = 3'h5 == state ? _GEN_9026 : ram_0_35; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10058 = 3'h5 == state ? _GEN_9027 : ram_0_36; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10059 = 3'h5 == state ? _GEN_9028 : ram_0_37; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10060 = 3'h5 == state ? _GEN_9029 : ram_0_38; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10061 = 3'h5 == state ? _GEN_9030 : ram_0_39; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10062 = 3'h5 == state ? _GEN_9031 : ram_0_40; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10063 = 3'h5 == state ? _GEN_9032 : ram_0_41; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10064 = 3'h5 == state ? _GEN_9033 : ram_0_42; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10065 = 3'h5 == state ? _GEN_9034 : ram_0_43; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10066 = 3'h5 == state ? _GEN_9035 : ram_0_44; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10067 = 3'h5 == state ? _GEN_9036 : ram_0_45; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10068 = 3'h5 == state ? _GEN_9037 : ram_0_46; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10069 = 3'h5 == state ? _GEN_9038 : ram_0_47; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10070 = 3'h5 == state ? _GEN_9039 : ram_0_48; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10071 = 3'h5 == state ? _GEN_9040 : ram_0_49; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10072 = 3'h5 == state ? _GEN_9041 : ram_0_50; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10073 = 3'h5 == state ? _GEN_9042 : ram_0_51; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10074 = 3'h5 == state ? _GEN_9043 : ram_0_52; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10075 = 3'h5 == state ? _GEN_9044 : ram_0_53; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10076 = 3'h5 == state ? _GEN_9045 : ram_0_54; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10077 = 3'h5 == state ? _GEN_9046 : ram_0_55; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10078 = 3'h5 == state ? _GEN_9047 : ram_0_56; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10079 = 3'h5 == state ? _GEN_9048 : ram_0_57; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10080 = 3'h5 == state ? _GEN_9049 : ram_0_58; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10081 = 3'h5 == state ? _GEN_9050 : ram_0_59; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10082 = 3'h5 == state ? _GEN_9051 : ram_0_60; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10083 = 3'h5 == state ? _GEN_9052 : ram_0_61; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10084 = 3'h5 == state ? _GEN_9053 : ram_0_62; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10085 = 3'h5 == state ? _GEN_9054 : ram_0_63; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10086 = 3'h5 == state ? _GEN_9055 : ram_0_64; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10087 = 3'h5 == state ? _GEN_9056 : ram_0_65; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10088 = 3'h5 == state ? _GEN_9057 : ram_0_66; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10089 = 3'h5 == state ? _GEN_9058 : ram_0_67; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10090 = 3'h5 == state ? _GEN_9059 : ram_0_68; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10091 = 3'h5 == state ? _GEN_9060 : ram_0_69; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10092 = 3'h5 == state ? _GEN_9061 : ram_0_70; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10093 = 3'h5 == state ? _GEN_9062 : ram_0_71; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10094 = 3'h5 == state ? _GEN_9063 : ram_0_72; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10095 = 3'h5 == state ? _GEN_9064 : ram_0_73; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10096 = 3'h5 == state ? _GEN_9065 : ram_0_74; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10097 = 3'h5 == state ? _GEN_9066 : ram_0_75; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10098 = 3'h5 == state ? _GEN_9067 : ram_0_76; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10099 = 3'h5 == state ? _GEN_9068 : ram_0_77; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10100 = 3'h5 == state ? _GEN_9069 : ram_0_78; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10101 = 3'h5 == state ? _GEN_9070 : ram_0_79; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10102 = 3'h5 == state ? _GEN_9071 : ram_0_80; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10103 = 3'h5 == state ? _GEN_9072 : ram_0_81; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10104 = 3'h5 == state ? _GEN_9073 : ram_0_82; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10105 = 3'h5 == state ? _GEN_9074 : ram_0_83; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10106 = 3'h5 == state ? _GEN_9075 : ram_0_84; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10107 = 3'h5 == state ? _GEN_9076 : ram_0_85; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10108 = 3'h5 == state ? _GEN_9077 : ram_0_86; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10109 = 3'h5 == state ? _GEN_9078 : ram_0_87; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10110 = 3'h5 == state ? _GEN_9079 : ram_0_88; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10111 = 3'h5 == state ? _GEN_9080 : ram_0_89; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10112 = 3'h5 == state ? _GEN_9081 : ram_0_90; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10113 = 3'h5 == state ? _GEN_9082 : ram_0_91; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10114 = 3'h5 == state ? _GEN_9083 : ram_0_92; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10115 = 3'h5 == state ? _GEN_9084 : ram_0_93; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10116 = 3'h5 == state ? _GEN_9085 : ram_0_94; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10117 = 3'h5 == state ? _GEN_9086 : ram_0_95; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10118 = 3'h5 == state ? _GEN_9087 : ram_0_96; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10119 = 3'h5 == state ? _GEN_9088 : ram_0_97; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10120 = 3'h5 == state ? _GEN_9089 : ram_0_98; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10121 = 3'h5 == state ? _GEN_9090 : ram_0_99; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10122 = 3'h5 == state ? _GEN_9091 : ram_0_100; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10123 = 3'h5 == state ? _GEN_9092 : ram_0_101; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10124 = 3'h5 == state ? _GEN_9093 : ram_0_102; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10125 = 3'h5 == state ? _GEN_9094 : ram_0_103; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10126 = 3'h5 == state ? _GEN_9095 : ram_0_104; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10127 = 3'h5 == state ? _GEN_9096 : ram_0_105; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10128 = 3'h5 == state ? _GEN_9097 : ram_0_106; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10129 = 3'h5 == state ? _GEN_9098 : ram_0_107; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10130 = 3'h5 == state ? _GEN_9099 : ram_0_108; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10131 = 3'h5 == state ? _GEN_9100 : ram_0_109; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10132 = 3'h5 == state ? _GEN_9101 : ram_0_110; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10133 = 3'h5 == state ? _GEN_9102 : ram_0_111; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10134 = 3'h5 == state ? _GEN_9103 : ram_0_112; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10135 = 3'h5 == state ? _GEN_9104 : ram_0_113; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10136 = 3'h5 == state ? _GEN_9105 : ram_0_114; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10137 = 3'h5 == state ? _GEN_9106 : ram_0_115; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10138 = 3'h5 == state ? _GEN_9107 : ram_0_116; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10139 = 3'h5 == state ? _GEN_9108 : ram_0_117; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10140 = 3'h5 == state ? _GEN_9109 : ram_0_118; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10141 = 3'h5 == state ? _GEN_9110 : ram_0_119; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10142 = 3'h5 == state ? _GEN_9111 : ram_0_120; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10143 = 3'h5 == state ? _GEN_9112 : ram_0_121; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10144 = 3'h5 == state ? _GEN_9113 : ram_0_122; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10145 = 3'h5 == state ? _GEN_9114 : ram_0_123; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10146 = 3'h5 == state ? _GEN_9115 : ram_0_124; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10147 = 3'h5 == state ? _GEN_9116 : ram_0_125; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10148 = 3'h5 == state ? _GEN_9117 : ram_0_126; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_10149 = 3'h5 == state ? _GEN_9118 : ram_0_127; // @[d_cache.scala 78:18 18:24]
  wire [31:0] _GEN_10150 = 3'h5 == state ? _GEN_9119 : tag_0_0; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10151 = 3'h5 == state ? _GEN_9120 : tag_0_1; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10152 = 3'h5 == state ? _GEN_9121 : tag_0_2; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10153 = 3'h5 == state ? _GEN_9122 : tag_0_3; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10154 = 3'h5 == state ? _GEN_9123 : tag_0_4; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10155 = 3'h5 == state ? _GEN_9124 : tag_0_5; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10156 = 3'h5 == state ? _GEN_9125 : tag_0_6; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10157 = 3'h5 == state ? _GEN_9126 : tag_0_7; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10158 = 3'h5 == state ? _GEN_9127 : tag_0_8; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10159 = 3'h5 == state ? _GEN_9128 : tag_0_9; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10160 = 3'h5 == state ? _GEN_9129 : tag_0_10; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10161 = 3'h5 == state ? _GEN_9130 : tag_0_11; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10162 = 3'h5 == state ? _GEN_9131 : tag_0_12; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10163 = 3'h5 == state ? _GEN_9132 : tag_0_13; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10164 = 3'h5 == state ? _GEN_9133 : tag_0_14; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10165 = 3'h5 == state ? _GEN_9134 : tag_0_15; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10166 = 3'h5 == state ? _GEN_9135 : tag_0_16; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10167 = 3'h5 == state ? _GEN_9136 : tag_0_17; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10168 = 3'h5 == state ? _GEN_9137 : tag_0_18; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10169 = 3'h5 == state ? _GEN_9138 : tag_0_19; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10170 = 3'h5 == state ? _GEN_9139 : tag_0_20; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10171 = 3'h5 == state ? _GEN_9140 : tag_0_21; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10172 = 3'h5 == state ? _GEN_9141 : tag_0_22; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10173 = 3'h5 == state ? _GEN_9142 : tag_0_23; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10174 = 3'h5 == state ? _GEN_9143 : tag_0_24; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10175 = 3'h5 == state ? _GEN_9144 : tag_0_25; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10176 = 3'h5 == state ? _GEN_9145 : tag_0_26; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10177 = 3'h5 == state ? _GEN_9146 : tag_0_27; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10178 = 3'h5 == state ? _GEN_9147 : tag_0_28; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10179 = 3'h5 == state ? _GEN_9148 : tag_0_29; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10180 = 3'h5 == state ? _GEN_9149 : tag_0_30; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10181 = 3'h5 == state ? _GEN_9150 : tag_0_31; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10182 = 3'h5 == state ? _GEN_9151 : tag_0_32; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10183 = 3'h5 == state ? _GEN_9152 : tag_0_33; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10184 = 3'h5 == state ? _GEN_9153 : tag_0_34; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10185 = 3'h5 == state ? _GEN_9154 : tag_0_35; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10186 = 3'h5 == state ? _GEN_9155 : tag_0_36; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10187 = 3'h5 == state ? _GEN_9156 : tag_0_37; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10188 = 3'h5 == state ? _GEN_9157 : tag_0_38; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10189 = 3'h5 == state ? _GEN_9158 : tag_0_39; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10190 = 3'h5 == state ? _GEN_9159 : tag_0_40; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10191 = 3'h5 == state ? _GEN_9160 : tag_0_41; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10192 = 3'h5 == state ? _GEN_9161 : tag_0_42; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10193 = 3'h5 == state ? _GEN_9162 : tag_0_43; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10194 = 3'h5 == state ? _GEN_9163 : tag_0_44; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10195 = 3'h5 == state ? _GEN_9164 : tag_0_45; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10196 = 3'h5 == state ? _GEN_9165 : tag_0_46; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10197 = 3'h5 == state ? _GEN_9166 : tag_0_47; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10198 = 3'h5 == state ? _GEN_9167 : tag_0_48; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10199 = 3'h5 == state ? _GEN_9168 : tag_0_49; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10200 = 3'h5 == state ? _GEN_9169 : tag_0_50; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10201 = 3'h5 == state ? _GEN_9170 : tag_0_51; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10202 = 3'h5 == state ? _GEN_9171 : tag_0_52; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10203 = 3'h5 == state ? _GEN_9172 : tag_0_53; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10204 = 3'h5 == state ? _GEN_9173 : tag_0_54; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10205 = 3'h5 == state ? _GEN_9174 : tag_0_55; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10206 = 3'h5 == state ? _GEN_9175 : tag_0_56; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10207 = 3'h5 == state ? _GEN_9176 : tag_0_57; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10208 = 3'h5 == state ? _GEN_9177 : tag_0_58; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10209 = 3'h5 == state ? _GEN_9178 : tag_0_59; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10210 = 3'h5 == state ? _GEN_9179 : tag_0_60; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10211 = 3'h5 == state ? _GEN_9180 : tag_0_61; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10212 = 3'h5 == state ? _GEN_9181 : tag_0_62; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10213 = 3'h5 == state ? _GEN_9182 : tag_0_63; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10214 = 3'h5 == state ? _GEN_9183 : tag_0_64; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10215 = 3'h5 == state ? _GEN_9184 : tag_0_65; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10216 = 3'h5 == state ? _GEN_9185 : tag_0_66; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10217 = 3'h5 == state ? _GEN_9186 : tag_0_67; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10218 = 3'h5 == state ? _GEN_9187 : tag_0_68; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10219 = 3'h5 == state ? _GEN_9188 : tag_0_69; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10220 = 3'h5 == state ? _GEN_9189 : tag_0_70; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10221 = 3'h5 == state ? _GEN_9190 : tag_0_71; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10222 = 3'h5 == state ? _GEN_9191 : tag_0_72; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10223 = 3'h5 == state ? _GEN_9192 : tag_0_73; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10224 = 3'h5 == state ? _GEN_9193 : tag_0_74; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10225 = 3'h5 == state ? _GEN_9194 : tag_0_75; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10226 = 3'h5 == state ? _GEN_9195 : tag_0_76; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10227 = 3'h5 == state ? _GEN_9196 : tag_0_77; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10228 = 3'h5 == state ? _GEN_9197 : tag_0_78; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10229 = 3'h5 == state ? _GEN_9198 : tag_0_79; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10230 = 3'h5 == state ? _GEN_9199 : tag_0_80; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10231 = 3'h5 == state ? _GEN_9200 : tag_0_81; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10232 = 3'h5 == state ? _GEN_9201 : tag_0_82; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10233 = 3'h5 == state ? _GEN_9202 : tag_0_83; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10234 = 3'h5 == state ? _GEN_9203 : tag_0_84; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10235 = 3'h5 == state ? _GEN_9204 : tag_0_85; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10236 = 3'h5 == state ? _GEN_9205 : tag_0_86; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10237 = 3'h5 == state ? _GEN_9206 : tag_0_87; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10238 = 3'h5 == state ? _GEN_9207 : tag_0_88; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10239 = 3'h5 == state ? _GEN_9208 : tag_0_89; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10240 = 3'h5 == state ? _GEN_9209 : tag_0_90; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10241 = 3'h5 == state ? _GEN_9210 : tag_0_91; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10242 = 3'h5 == state ? _GEN_9211 : tag_0_92; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10243 = 3'h5 == state ? _GEN_9212 : tag_0_93; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10244 = 3'h5 == state ? _GEN_9213 : tag_0_94; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10245 = 3'h5 == state ? _GEN_9214 : tag_0_95; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10246 = 3'h5 == state ? _GEN_9215 : tag_0_96; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10247 = 3'h5 == state ? _GEN_9216 : tag_0_97; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10248 = 3'h5 == state ? _GEN_9217 : tag_0_98; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10249 = 3'h5 == state ? _GEN_9218 : tag_0_99; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10250 = 3'h5 == state ? _GEN_9219 : tag_0_100; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10251 = 3'h5 == state ? _GEN_9220 : tag_0_101; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10252 = 3'h5 == state ? _GEN_9221 : tag_0_102; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10253 = 3'h5 == state ? _GEN_9222 : tag_0_103; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10254 = 3'h5 == state ? _GEN_9223 : tag_0_104; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10255 = 3'h5 == state ? _GEN_9224 : tag_0_105; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10256 = 3'h5 == state ? _GEN_9225 : tag_0_106; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10257 = 3'h5 == state ? _GEN_9226 : tag_0_107; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10258 = 3'h5 == state ? _GEN_9227 : tag_0_108; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10259 = 3'h5 == state ? _GEN_9228 : tag_0_109; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10260 = 3'h5 == state ? _GEN_9229 : tag_0_110; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10261 = 3'h5 == state ? _GEN_9230 : tag_0_111; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10262 = 3'h5 == state ? _GEN_9231 : tag_0_112; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10263 = 3'h5 == state ? _GEN_9232 : tag_0_113; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10264 = 3'h5 == state ? _GEN_9233 : tag_0_114; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10265 = 3'h5 == state ? _GEN_9234 : tag_0_115; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10266 = 3'h5 == state ? _GEN_9235 : tag_0_116; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10267 = 3'h5 == state ? _GEN_9236 : tag_0_117; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10268 = 3'h5 == state ? _GEN_9237 : tag_0_118; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10269 = 3'h5 == state ? _GEN_9238 : tag_0_119; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10270 = 3'h5 == state ? _GEN_9239 : tag_0_120; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10271 = 3'h5 == state ? _GEN_9240 : tag_0_121; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10272 = 3'h5 == state ? _GEN_9241 : tag_0_122; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10273 = 3'h5 == state ? _GEN_9242 : tag_0_123; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10274 = 3'h5 == state ? _GEN_9243 : tag_0_124; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10275 = 3'h5 == state ? _GEN_9244 : tag_0_125; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10276 = 3'h5 == state ? _GEN_9245 : tag_0_126; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_10277 = 3'h5 == state ? _GEN_9246 : tag_0_127; // @[d_cache.scala 78:18 20:24]
  wire  _GEN_10278 = 3'h5 == state ? _GEN_9247 : valid_0_0; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10279 = 3'h5 == state ? _GEN_9248 : valid_0_1; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10280 = 3'h5 == state ? _GEN_9249 : valid_0_2; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10281 = 3'h5 == state ? _GEN_9250 : valid_0_3; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10282 = 3'h5 == state ? _GEN_9251 : valid_0_4; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10283 = 3'h5 == state ? _GEN_9252 : valid_0_5; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10284 = 3'h5 == state ? _GEN_9253 : valid_0_6; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10285 = 3'h5 == state ? _GEN_9254 : valid_0_7; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10286 = 3'h5 == state ? _GEN_9255 : valid_0_8; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10287 = 3'h5 == state ? _GEN_9256 : valid_0_9; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10288 = 3'h5 == state ? _GEN_9257 : valid_0_10; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10289 = 3'h5 == state ? _GEN_9258 : valid_0_11; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10290 = 3'h5 == state ? _GEN_9259 : valid_0_12; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10291 = 3'h5 == state ? _GEN_9260 : valid_0_13; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10292 = 3'h5 == state ? _GEN_9261 : valid_0_14; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10293 = 3'h5 == state ? _GEN_9262 : valid_0_15; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10294 = 3'h5 == state ? _GEN_9263 : valid_0_16; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10295 = 3'h5 == state ? _GEN_9264 : valid_0_17; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10296 = 3'h5 == state ? _GEN_9265 : valid_0_18; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10297 = 3'h5 == state ? _GEN_9266 : valid_0_19; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10298 = 3'h5 == state ? _GEN_9267 : valid_0_20; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10299 = 3'h5 == state ? _GEN_9268 : valid_0_21; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10300 = 3'h5 == state ? _GEN_9269 : valid_0_22; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10301 = 3'h5 == state ? _GEN_9270 : valid_0_23; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10302 = 3'h5 == state ? _GEN_9271 : valid_0_24; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10303 = 3'h5 == state ? _GEN_9272 : valid_0_25; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10304 = 3'h5 == state ? _GEN_9273 : valid_0_26; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10305 = 3'h5 == state ? _GEN_9274 : valid_0_27; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10306 = 3'h5 == state ? _GEN_9275 : valid_0_28; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10307 = 3'h5 == state ? _GEN_9276 : valid_0_29; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10308 = 3'h5 == state ? _GEN_9277 : valid_0_30; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10309 = 3'h5 == state ? _GEN_9278 : valid_0_31; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10310 = 3'h5 == state ? _GEN_9279 : valid_0_32; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10311 = 3'h5 == state ? _GEN_9280 : valid_0_33; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10312 = 3'h5 == state ? _GEN_9281 : valid_0_34; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10313 = 3'h5 == state ? _GEN_9282 : valid_0_35; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10314 = 3'h5 == state ? _GEN_9283 : valid_0_36; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10315 = 3'h5 == state ? _GEN_9284 : valid_0_37; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10316 = 3'h5 == state ? _GEN_9285 : valid_0_38; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10317 = 3'h5 == state ? _GEN_9286 : valid_0_39; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10318 = 3'h5 == state ? _GEN_9287 : valid_0_40; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10319 = 3'h5 == state ? _GEN_9288 : valid_0_41; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10320 = 3'h5 == state ? _GEN_9289 : valid_0_42; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10321 = 3'h5 == state ? _GEN_9290 : valid_0_43; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10322 = 3'h5 == state ? _GEN_9291 : valid_0_44; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10323 = 3'h5 == state ? _GEN_9292 : valid_0_45; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10324 = 3'h5 == state ? _GEN_9293 : valid_0_46; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10325 = 3'h5 == state ? _GEN_9294 : valid_0_47; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10326 = 3'h5 == state ? _GEN_9295 : valid_0_48; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10327 = 3'h5 == state ? _GEN_9296 : valid_0_49; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10328 = 3'h5 == state ? _GEN_9297 : valid_0_50; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10329 = 3'h5 == state ? _GEN_9298 : valid_0_51; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10330 = 3'h5 == state ? _GEN_9299 : valid_0_52; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10331 = 3'h5 == state ? _GEN_9300 : valid_0_53; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10332 = 3'h5 == state ? _GEN_9301 : valid_0_54; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10333 = 3'h5 == state ? _GEN_9302 : valid_0_55; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10334 = 3'h5 == state ? _GEN_9303 : valid_0_56; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10335 = 3'h5 == state ? _GEN_9304 : valid_0_57; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10336 = 3'h5 == state ? _GEN_9305 : valid_0_58; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10337 = 3'h5 == state ? _GEN_9306 : valid_0_59; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10338 = 3'h5 == state ? _GEN_9307 : valid_0_60; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10339 = 3'h5 == state ? _GEN_9308 : valid_0_61; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10340 = 3'h5 == state ? _GEN_9309 : valid_0_62; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10341 = 3'h5 == state ? _GEN_9310 : valid_0_63; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10342 = 3'h5 == state ? _GEN_9311 : valid_0_64; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10343 = 3'h5 == state ? _GEN_9312 : valid_0_65; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10344 = 3'h5 == state ? _GEN_9313 : valid_0_66; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10345 = 3'h5 == state ? _GEN_9314 : valid_0_67; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10346 = 3'h5 == state ? _GEN_9315 : valid_0_68; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10347 = 3'h5 == state ? _GEN_9316 : valid_0_69; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10348 = 3'h5 == state ? _GEN_9317 : valid_0_70; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10349 = 3'h5 == state ? _GEN_9318 : valid_0_71; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10350 = 3'h5 == state ? _GEN_9319 : valid_0_72; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10351 = 3'h5 == state ? _GEN_9320 : valid_0_73; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10352 = 3'h5 == state ? _GEN_9321 : valid_0_74; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10353 = 3'h5 == state ? _GEN_9322 : valid_0_75; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10354 = 3'h5 == state ? _GEN_9323 : valid_0_76; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10355 = 3'h5 == state ? _GEN_9324 : valid_0_77; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10356 = 3'h5 == state ? _GEN_9325 : valid_0_78; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10357 = 3'h5 == state ? _GEN_9326 : valid_0_79; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10358 = 3'h5 == state ? _GEN_9327 : valid_0_80; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10359 = 3'h5 == state ? _GEN_9328 : valid_0_81; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10360 = 3'h5 == state ? _GEN_9329 : valid_0_82; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10361 = 3'h5 == state ? _GEN_9330 : valid_0_83; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10362 = 3'h5 == state ? _GEN_9331 : valid_0_84; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10363 = 3'h5 == state ? _GEN_9332 : valid_0_85; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10364 = 3'h5 == state ? _GEN_9333 : valid_0_86; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10365 = 3'h5 == state ? _GEN_9334 : valid_0_87; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10366 = 3'h5 == state ? _GEN_9335 : valid_0_88; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10367 = 3'h5 == state ? _GEN_9336 : valid_0_89; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10368 = 3'h5 == state ? _GEN_9337 : valid_0_90; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10369 = 3'h5 == state ? _GEN_9338 : valid_0_91; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10370 = 3'h5 == state ? _GEN_9339 : valid_0_92; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10371 = 3'h5 == state ? _GEN_9340 : valid_0_93; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10372 = 3'h5 == state ? _GEN_9341 : valid_0_94; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10373 = 3'h5 == state ? _GEN_9342 : valid_0_95; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10374 = 3'h5 == state ? _GEN_9343 : valid_0_96; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10375 = 3'h5 == state ? _GEN_9344 : valid_0_97; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10376 = 3'h5 == state ? _GEN_9345 : valid_0_98; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10377 = 3'h5 == state ? _GEN_9346 : valid_0_99; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10378 = 3'h5 == state ? _GEN_9347 : valid_0_100; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10379 = 3'h5 == state ? _GEN_9348 : valid_0_101; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10380 = 3'h5 == state ? _GEN_9349 : valid_0_102; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10381 = 3'h5 == state ? _GEN_9350 : valid_0_103; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10382 = 3'h5 == state ? _GEN_9351 : valid_0_104; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10383 = 3'h5 == state ? _GEN_9352 : valid_0_105; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10384 = 3'h5 == state ? _GEN_9353 : valid_0_106; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10385 = 3'h5 == state ? _GEN_9354 : valid_0_107; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10386 = 3'h5 == state ? _GEN_9355 : valid_0_108; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10387 = 3'h5 == state ? _GEN_9356 : valid_0_109; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10388 = 3'h5 == state ? _GEN_9357 : valid_0_110; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10389 = 3'h5 == state ? _GEN_9358 : valid_0_111; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10390 = 3'h5 == state ? _GEN_9359 : valid_0_112; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10391 = 3'h5 == state ? _GEN_9360 : valid_0_113; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10392 = 3'h5 == state ? _GEN_9361 : valid_0_114; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10393 = 3'h5 == state ? _GEN_9362 : valid_0_115; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10394 = 3'h5 == state ? _GEN_9363 : valid_0_116; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10395 = 3'h5 == state ? _GEN_9364 : valid_0_117; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10396 = 3'h5 == state ? _GEN_9365 : valid_0_118; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10397 = 3'h5 == state ? _GEN_9366 : valid_0_119; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10398 = 3'h5 == state ? _GEN_9367 : valid_0_120; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10399 = 3'h5 == state ? _GEN_9368 : valid_0_121; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10400 = 3'h5 == state ? _GEN_9369 : valid_0_122; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10401 = 3'h5 == state ? _GEN_9370 : valid_0_123; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10402 = 3'h5 == state ? _GEN_9371 : valid_0_124; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10403 = 3'h5 == state ? _GEN_9372 : valid_0_125; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10404 = 3'h5 == state ? _GEN_9373 : valid_0_126; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10405 = 3'h5 == state ? _GEN_9374 : valid_0_127; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_10406 = 3'h5 == state ? _GEN_9375 : quene; // @[d_cache.scala 78:18 35:24]
  wire [63:0] _GEN_10407 = 3'h5 == state ? _GEN_9376 : ram_1_0; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10408 = 3'h5 == state ? _GEN_9377 : ram_1_1; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10409 = 3'h5 == state ? _GEN_9378 : ram_1_2; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10410 = 3'h5 == state ? _GEN_9379 : ram_1_3; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10411 = 3'h5 == state ? _GEN_9380 : ram_1_4; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10412 = 3'h5 == state ? _GEN_9381 : ram_1_5; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10413 = 3'h5 == state ? _GEN_9382 : ram_1_6; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10414 = 3'h5 == state ? _GEN_9383 : ram_1_7; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10415 = 3'h5 == state ? _GEN_9384 : ram_1_8; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10416 = 3'h5 == state ? _GEN_9385 : ram_1_9; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10417 = 3'h5 == state ? _GEN_9386 : ram_1_10; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10418 = 3'h5 == state ? _GEN_9387 : ram_1_11; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10419 = 3'h5 == state ? _GEN_9388 : ram_1_12; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10420 = 3'h5 == state ? _GEN_9389 : ram_1_13; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10421 = 3'h5 == state ? _GEN_9390 : ram_1_14; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10422 = 3'h5 == state ? _GEN_9391 : ram_1_15; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10423 = 3'h5 == state ? _GEN_9392 : ram_1_16; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10424 = 3'h5 == state ? _GEN_9393 : ram_1_17; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10425 = 3'h5 == state ? _GEN_9394 : ram_1_18; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10426 = 3'h5 == state ? _GEN_9395 : ram_1_19; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10427 = 3'h5 == state ? _GEN_9396 : ram_1_20; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10428 = 3'h5 == state ? _GEN_9397 : ram_1_21; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10429 = 3'h5 == state ? _GEN_9398 : ram_1_22; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10430 = 3'h5 == state ? _GEN_9399 : ram_1_23; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10431 = 3'h5 == state ? _GEN_9400 : ram_1_24; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10432 = 3'h5 == state ? _GEN_9401 : ram_1_25; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10433 = 3'h5 == state ? _GEN_9402 : ram_1_26; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10434 = 3'h5 == state ? _GEN_9403 : ram_1_27; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10435 = 3'h5 == state ? _GEN_9404 : ram_1_28; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10436 = 3'h5 == state ? _GEN_9405 : ram_1_29; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10437 = 3'h5 == state ? _GEN_9406 : ram_1_30; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10438 = 3'h5 == state ? _GEN_9407 : ram_1_31; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10439 = 3'h5 == state ? _GEN_9408 : ram_1_32; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10440 = 3'h5 == state ? _GEN_9409 : ram_1_33; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10441 = 3'h5 == state ? _GEN_9410 : ram_1_34; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10442 = 3'h5 == state ? _GEN_9411 : ram_1_35; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10443 = 3'h5 == state ? _GEN_9412 : ram_1_36; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10444 = 3'h5 == state ? _GEN_9413 : ram_1_37; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10445 = 3'h5 == state ? _GEN_9414 : ram_1_38; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10446 = 3'h5 == state ? _GEN_9415 : ram_1_39; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10447 = 3'h5 == state ? _GEN_9416 : ram_1_40; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10448 = 3'h5 == state ? _GEN_9417 : ram_1_41; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10449 = 3'h5 == state ? _GEN_9418 : ram_1_42; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10450 = 3'h5 == state ? _GEN_9419 : ram_1_43; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10451 = 3'h5 == state ? _GEN_9420 : ram_1_44; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10452 = 3'h5 == state ? _GEN_9421 : ram_1_45; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10453 = 3'h5 == state ? _GEN_9422 : ram_1_46; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10454 = 3'h5 == state ? _GEN_9423 : ram_1_47; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10455 = 3'h5 == state ? _GEN_9424 : ram_1_48; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10456 = 3'h5 == state ? _GEN_9425 : ram_1_49; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10457 = 3'h5 == state ? _GEN_9426 : ram_1_50; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10458 = 3'h5 == state ? _GEN_9427 : ram_1_51; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10459 = 3'h5 == state ? _GEN_9428 : ram_1_52; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10460 = 3'h5 == state ? _GEN_9429 : ram_1_53; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10461 = 3'h5 == state ? _GEN_9430 : ram_1_54; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10462 = 3'h5 == state ? _GEN_9431 : ram_1_55; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10463 = 3'h5 == state ? _GEN_9432 : ram_1_56; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10464 = 3'h5 == state ? _GEN_9433 : ram_1_57; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10465 = 3'h5 == state ? _GEN_9434 : ram_1_58; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10466 = 3'h5 == state ? _GEN_9435 : ram_1_59; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10467 = 3'h5 == state ? _GEN_9436 : ram_1_60; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10468 = 3'h5 == state ? _GEN_9437 : ram_1_61; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10469 = 3'h5 == state ? _GEN_9438 : ram_1_62; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10470 = 3'h5 == state ? _GEN_9439 : ram_1_63; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10471 = 3'h5 == state ? _GEN_9440 : ram_1_64; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10472 = 3'h5 == state ? _GEN_9441 : ram_1_65; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10473 = 3'h5 == state ? _GEN_9442 : ram_1_66; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10474 = 3'h5 == state ? _GEN_9443 : ram_1_67; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10475 = 3'h5 == state ? _GEN_9444 : ram_1_68; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10476 = 3'h5 == state ? _GEN_9445 : ram_1_69; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10477 = 3'h5 == state ? _GEN_9446 : ram_1_70; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10478 = 3'h5 == state ? _GEN_9447 : ram_1_71; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10479 = 3'h5 == state ? _GEN_9448 : ram_1_72; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10480 = 3'h5 == state ? _GEN_9449 : ram_1_73; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10481 = 3'h5 == state ? _GEN_9450 : ram_1_74; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10482 = 3'h5 == state ? _GEN_9451 : ram_1_75; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10483 = 3'h5 == state ? _GEN_9452 : ram_1_76; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10484 = 3'h5 == state ? _GEN_9453 : ram_1_77; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10485 = 3'h5 == state ? _GEN_9454 : ram_1_78; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10486 = 3'h5 == state ? _GEN_9455 : ram_1_79; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10487 = 3'h5 == state ? _GEN_9456 : ram_1_80; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10488 = 3'h5 == state ? _GEN_9457 : ram_1_81; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10489 = 3'h5 == state ? _GEN_9458 : ram_1_82; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10490 = 3'h5 == state ? _GEN_9459 : ram_1_83; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10491 = 3'h5 == state ? _GEN_9460 : ram_1_84; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10492 = 3'h5 == state ? _GEN_9461 : ram_1_85; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10493 = 3'h5 == state ? _GEN_9462 : ram_1_86; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10494 = 3'h5 == state ? _GEN_9463 : ram_1_87; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10495 = 3'h5 == state ? _GEN_9464 : ram_1_88; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10496 = 3'h5 == state ? _GEN_9465 : ram_1_89; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10497 = 3'h5 == state ? _GEN_9466 : ram_1_90; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10498 = 3'h5 == state ? _GEN_9467 : ram_1_91; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10499 = 3'h5 == state ? _GEN_9468 : ram_1_92; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10500 = 3'h5 == state ? _GEN_9469 : ram_1_93; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10501 = 3'h5 == state ? _GEN_9470 : ram_1_94; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10502 = 3'h5 == state ? _GEN_9471 : ram_1_95; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10503 = 3'h5 == state ? _GEN_9472 : ram_1_96; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10504 = 3'h5 == state ? _GEN_9473 : ram_1_97; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10505 = 3'h5 == state ? _GEN_9474 : ram_1_98; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10506 = 3'h5 == state ? _GEN_9475 : ram_1_99; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10507 = 3'h5 == state ? _GEN_9476 : ram_1_100; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10508 = 3'h5 == state ? _GEN_9477 : ram_1_101; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10509 = 3'h5 == state ? _GEN_9478 : ram_1_102; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10510 = 3'h5 == state ? _GEN_9479 : ram_1_103; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10511 = 3'h5 == state ? _GEN_9480 : ram_1_104; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10512 = 3'h5 == state ? _GEN_9481 : ram_1_105; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10513 = 3'h5 == state ? _GEN_9482 : ram_1_106; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10514 = 3'h5 == state ? _GEN_9483 : ram_1_107; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10515 = 3'h5 == state ? _GEN_9484 : ram_1_108; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10516 = 3'h5 == state ? _GEN_9485 : ram_1_109; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10517 = 3'h5 == state ? _GEN_9486 : ram_1_110; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10518 = 3'h5 == state ? _GEN_9487 : ram_1_111; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10519 = 3'h5 == state ? _GEN_9488 : ram_1_112; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10520 = 3'h5 == state ? _GEN_9489 : ram_1_113; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10521 = 3'h5 == state ? _GEN_9490 : ram_1_114; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10522 = 3'h5 == state ? _GEN_9491 : ram_1_115; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10523 = 3'h5 == state ? _GEN_9492 : ram_1_116; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10524 = 3'h5 == state ? _GEN_9493 : ram_1_117; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10525 = 3'h5 == state ? _GEN_9494 : ram_1_118; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10526 = 3'h5 == state ? _GEN_9495 : ram_1_119; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10527 = 3'h5 == state ? _GEN_9496 : ram_1_120; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10528 = 3'h5 == state ? _GEN_9497 : ram_1_121; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10529 = 3'h5 == state ? _GEN_9498 : ram_1_122; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10530 = 3'h5 == state ? _GEN_9499 : ram_1_123; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10531 = 3'h5 == state ? _GEN_9500 : ram_1_124; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10532 = 3'h5 == state ? _GEN_9501 : ram_1_125; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10533 = 3'h5 == state ? _GEN_9502 : ram_1_126; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_10534 = 3'h5 == state ? _GEN_9503 : ram_1_127; // @[d_cache.scala 78:18 19:24]
  wire [31:0] _GEN_10535 = 3'h5 == state ? _GEN_9504 : tag_1_0; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10536 = 3'h5 == state ? _GEN_9505 : tag_1_1; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10537 = 3'h5 == state ? _GEN_9506 : tag_1_2; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10538 = 3'h5 == state ? _GEN_9507 : tag_1_3; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10539 = 3'h5 == state ? _GEN_9508 : tag_1_4; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10540 = 3'h5 == state ? _GEN_9509 : tag_1_5; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10541 = 3'h5 == state ? _GEN_9510 : tag_1_6; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10542 = 3'h5 == state ? _GEN_9511 : tag_1_7; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10543 = 3'h5 == state ? _GEN_9512 : tag_1_8; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10544 = 3'h5 == state ? _GEN_9513 : tag_1_9; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10545 = 3'h5 == state ? _GEN_9514 : tag_1_10; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10546 = 3'h5 == state ? _GEN_9515 : tag_1_11; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10547 = 3'h5 == state ? _GEN_9516 : tag_1_12; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10548 = 3'h5 == state ? _GEN_9517 : tag_1_13; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10549 = 3'h5 == state ? _GEN_9518 : tag_1_14; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10550 = 3'h5 == state ? _GEN_9519 : tag_1_15; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10551 = 3'h5 == state ? _GEN_9520 : tag_1_16; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10552 = 3'h5 == state ? _GEN_9521 : tag_1_17; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10553 = 3'h5 == state ? _GEN_9522 : tag_1_18; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10554 = 3'h5 == state ? _GEN_9523 : tag_1_19; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10555 = 3'h5 == state ? _GEN_9524 : tag_1_20; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10556 = 3'h5 == state ? _GEN_9525 : tag_1_21; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10557 = 3'h5 == state ? _GEN_9526 : tag_1_22; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10558 = 3'h5 == state ? _GEN_9527 : tag_1_23; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10559 = 3'h5 == state ? _GEN_9528 : tag_1_24; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10560 = 3'h5 == state ? _GEN_9529 : tag_1_25; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10561 = 3'h5 == state ? _GEN_9530 : tag_1_26; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10562 = 3'h5 == state ? _GEN_9531 : tag_1_27; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10563 = 3'h5 == state ? _GEN_9532 : tag_1_28; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10564 = 3'h5 == state ? _GEN_9533 : tag_1_29; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10565 = 3'h5 == state ? _GEN_9534 : tag_1_30; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10566 = 3'h5 == state ? _GEN_9535 : tag_1_31; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10567 = 3'h5 == state ? _GEN_9536 : tag_1_32; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10568 = 3'h5 == state ? _GEN_9537 : tag_1_33; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10569 = 3'h5 == state ? _GEN_9538 : tag_1_34; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10570 = 3'h5 == state ? _GEN_9539 : tag_1_35; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10571 = 3'h5 == state ? _GEN_9540 : tag_1_36; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10572 = 3'h5 == state ? _GEN_9541 : tag_1_37; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10573 = 3'h5 == state ? _GEN_9542 : tag_1_38; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10574 = 3'h5 == state ? _GEN_9543 : tag_1_39; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10575 = 3'h5 == state ? _GEN_9544 : tag_1_40; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10576 = 3'h5 == state ? _GEN_9545 : tag_1_41; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10577 = 3'h5 == state ? _GEN_9546 : tag_1_42; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10578 = 3'h5 == state ? _GEN_9547 : tag_1_43; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10579 = 3'h5 == state ? _GEN_9548 : tag_1_44; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10580 = 3'h5 == state ? _GEN_9549 : tag_1_45; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10581 = 3'h5 == state ? _GEN_9550 : tag_1_46; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10582 = 3'h5 == state ? _GEN_9551 : tag_1_47; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10583 = 3'h5 == state ? _GEN_9552 : tag_1_48; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10584 = 3'h5 == state ? _GEN_9553 : tag_1_49; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10585 = 3'h5 == state ? _GEN_9554 : tag_1_50; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10586 = 3'h5 == state ? _GEN_9555 : tag_1_51; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10587 = 3'h5 == state ? _GEN_9556 : tag_1_52; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10588 = 3'h5 == state ? _GEN_9557 : tag_1_53; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10589 = 3'h5 == state ? _GEN_9558 : tag_1_54; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10590 = 3'h5 == state ? _GEN_9559 : tag_1_55; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10591 = 3'h5 == state ? _GEN_9560 : tag_1_56; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10592 = 3'h5 == state ? _GEN_9561 : tag_1_57; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10593 = 3'h5 == state ? _GEN_9562 : tag_1_58; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10594 = 3'h5 == state ? _GEN_9563 : tag_1_59; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10595 = 3'h5 == state ? _GEN_9564 : tag_1_60; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10596 = 3'h5 == state ? _GEN_9565 : tag_1_61; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10597 = 3'h5 == state ? _GEN_9566 : tag_1_62; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10598 = 3'h5 == state ? _GEN_9567 : tag_1_63; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10599 = 3'h5 == state ? _GEN_9568 : tag_1_64; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10600 = 3'h5 == state ? _GEN_9569 : tag_1_65; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10601 = 3'h5 == state ? _GEN_9570 : tag_1_66; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10602 = 3'h5 == state ? _GEN_9571 : tag_1_67; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10603 = 3'h5 == state ? _GEN_9572 : tag_1_68; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10604 = 3'h5 == state ? _GEN_9573 : tag_1_69; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10605 = 3'h5 == state ? _GEN_9574 : tag_1_70; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10606 = 3'h5 == state ? _GEN_9575 : tag_1_71; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10607 = 3'h5 == state ? _GEN_9576 : tag_1_72; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10608 = 3'h5 == state ? _GEN_9577 : tag_1_73; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10609 = 3'h5 == state ? _GEN_9578 : tag_1_74; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10610 = 3'h5 == state ? _GEN_9579 : tag_1_75; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10611 = 3'h5 == state ? _GEN_9580 : tag_1_76; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10612 = 3'h5 == state ? _GEN_9581 : tag_1_77; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10613 = 3'h5 == state ? _GEN_9582 : tag_1_78; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10614 = 3'h5 == state ? _GEN_9583 : tag_1_79; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10615 = 3'h5 == state ? _GEN_9584 : tag_1_80; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10616 = 3'h5 == state ? _GEN_9585 : tag_1_81; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10617 = 3'h5 == state ? _GEN_9586 : tag_1_82; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10618 = 3'h5 == state ? _GEN_9587 : tag_1_83; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10619 = 3'h5 == state ? _GEN_9588 : tag_1_84; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10620 = 3'h5 == state ? _GEN_9589 : tag_1_85; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10621 = 3'h5 == state ? _GEN_9590 : tag_1_86; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10622 = 3'h5 == state ? _GEN_9591 : tag_1_87; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10623 = 3'h5 == state ? _GEN_9592 : tag_1_88; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10624 = 3'h5 == state ? _GEN_9593 : tag_1_89; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10625 = 3'h5 == state ? _GEN_9594 : tag_1_90; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10626 = 3'h5 == state ? _GEN_9595 : tag_1_91; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10627 = 3'h5 == state ? _GEN_9596 : tag_1_92; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10628 = 3'h5 == state ? _GEN_9597 : tag_1_93; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10629 = 3'h5 == state ? _GEN_9598 : tag_1_94; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10630 = 3'h5 == state ? _GEN_9599 : tag_1_95; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10631 = 3'h5 == state ? _GEN_9600 : tag_1_96; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10632 = 3'h5 == state ? _GEN_9601 : tag_1_97; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10633 = 3'h5 == state ? _GEN_9602 : tag_1_98; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10634 = 3'h5 == state ? _GEN_9603 : tag_1_99; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10635 = 3'h5 == state ? _GEN_9604 : tag_1_100; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10636 = 3'h5 == state ? _GEN_9605 : tag_1_101; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10637 = 3'h5 == state ? _GEN_9606 : tag_1_102; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10638 = 3'h5 == state ? _GEN_9607 : tag_1_103; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10639 = 3'h5 == state ? _GEN_9608 : tag_1_104; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10640 = 3'h5 == state ? _GEN_9609 : tag_1_105; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10641 = 3'h5 == state ? _GEN_9610 : tag_1_106; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10642 = 3'h5 == state ? _GEN_9611 : tag_1_107; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10643 = 3'h5 == state ? _GEN_9612 : tag_1_108; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10644 = 3'h5 == state ? _GEN_9613 : tag_1_109; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10645 = 3'h5 == state ? _GEN_9614 : tag_1_110; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10646 = 3'h5 == state ? _GEN_9615 : tag_1_111; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10647 = 3'h5 == state ? _GEN_9616 : tag_1_112; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10648 = 3'h5 == state ? _GEN_9617 : tag_1_113; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10649 = 3'h5 == state ? _GEN_9618 : tag_1_114; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10650 = 3'h5 == state ? _GEN_9619 : tag_1_115; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10651 = 3'h5 == state ? _GEN_9620 : tag_1_116; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10652 = 3'h5 == state ? _GEN_9621 : tag_1_117; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10653 = 3'h5 == state ? _GEN_9622 : tag_1_118; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10654 = 3'h5 == state ? _GEN_9623 : tag_1_119; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10655 = 3'h5 == state ? _GEN_9624 : tag_1_120; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10656 = 3'h5 == state ? _GEN_9625 : tag_1_121; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10657 = 3'h5 == state ? _GEN_9626 : tag_1_122; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10658 = 3'h5 == state ? _GEN_9627 : tag_1_123; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10659 = 3'h5 == state ? _GEN_9628 : tag_1_124; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10660 = 3'h5 == state ? _GEN_9629 : tag_1_125; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10661 = 3'h5 == state ? _GEN_9630 : tag_1_126; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_10662 = 3'h5 == state ? _GEN_9631 : tag_1_127; // @[d_cache.scala 78:18 21:24]
  wire  _GEN_10663 = 3'h5 == state ? _GEN_9632 : valid_1_0; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10664 = 3'h5 == state ? _GEN_9633 : valid_1_1; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10665 = 3'h5 == state ? _GEN_9634 : valid_1_2; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10666 = 3'h5 == state ? _GEN_9635 : valid_1_3; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10667 = 3'h5 == state ? _GEN_9636 : valid_1_4; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10668 = 3'h5 == state ? _GEN_9637 : valid_1_5; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10669 = 3'h5 == state ? _GEN_9638 : valid_1_6; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10670 = 3'h5 == state ? _GEN_9639 : valid_1_7; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10671 = 3'h5 == state ? _GEN_9640 : valid_1_8; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10672 = 3'h5 == state ? _GEN_9641 : valid_1_9; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10673 = 3'h5 == state ? _GEN_9642 : valid_1_10; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10674 = 3'h5 == state ? _GEN_9643 : valid_1_11; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10675 = 3'h5 == state ? _GEN_9644 : valid_1_12; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10676 = 3'h5 == state ? _GEN_9645 : valid_1_13; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10677 = 3'h5 == state ? _GEN_9646 : valid_1_14; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10678 = 3'h5 == state ? _GEN_9647 : valid_1_15; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10679 = 3'h5 == state ? _GEN_9648 : valid_1_16; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10680 = 3'h5 == state ? _GEN_9649 : valid_1_17; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10681 = 3'h5 == state ? _GEN_9650 : valid_1_18; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10682 = 3'h5 == state ? _GEN_9651 : valid_1_19; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10683 = 3'h5 == state ? _GEN_9652 : valid_1_20; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10684 = 3'h5 == state ? _GEN_9653 : valid_1_21; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10685 = 3'h5 == state ? _GEN_9654 : valid_1_22; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10686 = 3'h5 == state ? _GEN_9655 : valid_1_23; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10687 = 3'h5 == state ? _GEN_9656 : valid_1_24; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10688 = 3'h5 == state ? _GEN_9657 : valid_1_25; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10689 = 3'h5 == state ? _GEN_9658 : valid_1_26; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10690 = 3'h5 == state ? _GEN_9659 : valid_1_27; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10691 = 3'h5 == state ? _GEN_9660 : valid_1_28; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10692 = 3'h5 == state ? _GEN_9661 : valid_1_29; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10693 = 3'h5 == state ? _GEN_9662 : valid_1_30; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10694 = 3'h5 == state ? _GEN_9663 : valid_1_31; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10695 = 3'h5 == state ? _GEN_9664 : valid_1_32; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10696 = 3'h5 == state ? _GEN_9665 : valid_1_33; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10697 = 3'h5 == state ? _GEN_9666 : valid_1_34; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10698 = 3'h5 == state ? _GEN_9667 : valid_1_35; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10699 = 3'h5 == state ? _GEN_9668 : valid_1_36; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10700 = 3'h5 == state ? _GEN_9669 : valid_1_37; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10701 = 3'h5 == state ? _GEN_9670 : valid_1_38; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10702 = 3'h5 == state ? _GEN_9671 : valid_1_39; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10703 = 3'h5 == state ? _GEN_9672 : valid_1_40; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10704 = 3'h5 == state ? _GEN_9673 : valid_1_41; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10705 = 3'h5 == state ? _GEN_9674 : valid_1_42; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10706 = 3'h5 == state ? _GEN_9675 : valid_1_43; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10707 = 3'h5 == state ? _GEN_9676 : valid_1_44; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10708 = 3'h5 == state ? _GEN_9677 : valid_1_45; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10709 = 3'h5 == state ? _GEN_9678 : valid_1_46; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10710 = 3'h5 == state ? _GEN_9679 : valid_1_47; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10711 = 3'h5 == state ? _GEN_9680 : valid_1_48; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10712 = 3'h5 == state ? _GEN_9681 : valid_1_49; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10713 = 3'h5 == state ? _GEN_9682 : valid_1_50; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10714 = 3'h5 == state ? _GEN_9683 : valid_1_51; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10715 = 3'h5 == state ? _GEN_9684 : valid_1_52; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10716 = 3'h5 == state ? _GEN_9685 : valid_1_53; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10717 = 3'h5 == state ? _GEN_9686 : valid_1_54; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10718 = 3'h5 == state ? _GEN_9687 : valid_1_55; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10719 = 3'h5 == state ? _GEN_9688 : valid_1_56; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10720 = 3'h5 == state ? _GEN_9689 : valid_1_57; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10721 = 3'h5 == state ? _GEN_9690 : valid_1_58; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10722 = 3'h5 == state ? _GEN_9691 : valid_1_59; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10723 = 3'h5 == state ? _GEN_9692 : valid_1_60; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10724 = 3'h5 == state ? _GEN_9693 : valid_1_61; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10725 = 3'h5 == state ? _GEN_9694 : valid_1_62; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10726 = 3'h5 == state ? _GEN_9695 : valid_1_63; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10727 = 3'h5 == state ? _GEN_9696 : valid_1_64; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10728 = 3'h5 == state ? _GEN_9697 : valid_1_65; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10729 = 3'h5 == state ? _GEN_9698 : valid_1_66; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10730 = 3'h5 == state ? _GEN_9699 : valid_1_67; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10731 = 3'h5 == state ? _GEN_9700 : valid_1_68; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10732 = 3'h5 == state ? _GEN_9701 : valid_1_69; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10733 = 3'h5 == state ? _GEN_9702 : valid_1_70; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10734 = 3'h5 == state ? _GEN_9703 : valid_1_71; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10735 = 3'h5 == state ? _GEN_9704 : valid_1_72; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10736 = 3'h5 == state ? _GEN_9705 : valid_1_73; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10737 = 3'h5 == state ? _GEN_9706 : valid_1_74; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10738 = 3'h5 == state ? _GEN_9707 : valid_1_75; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10739 = 3'h5 == state ? _GEN_9708 : valid_1_76; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10740 = 3'h5 == state ? _GEN_9709 : valid_1_77; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10741 = 3'h5 == state ? _GEN_9710 : valid_1_78; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10742 = 3'h5 == state ? _GEN_9711 : valid_1_79; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10743 = 3'h5 == state ? _GEN_9712 : valid_1_80; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10744 = 3'h5 == state ? _GEN_9713 : valid_1_81; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10745 = 3'h5 == state ? _GEN_9714 : valid_1_82; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10746 = 3'h5 == state ? _GEN_9715 : valid_1_83; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10747 = 3'h5 == state ? _GEN_9716 : valid_1_84; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10748 = 3'h5 == state ? _GEN_9717 : valid_1_85; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10749 = 3'h5 == state ? _GEN_9718 : valid_1_86; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10750 = 3'h5 == state ? _GEN_9719 : valid_1_87; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10751 = 3'h5 == state ? _GEN_9720 : valid_1_88; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10752 = 3'h5 == state ? _GEN_9721 : valid_1_89; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10753 = 3'h5 == state ? _GEN_9722 : valid_1_90; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10754 = 3'h5 == state ? _GEN_9723 : valid_1_91; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10755 = 3'h5 == state ? _GEN_9724 : valid_1_92; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10756 = 3'h5 == state ? _GEN_9725 : valid_1_93; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10757 = 3'h5 == state ? _GEN_9726 : valid_1_94; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10758 = 3'h5 == state ? _GEN_9727 : valid_1_95; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10759 = 3'h5 == state ? _GEN_9728 : valid_1_96; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10760 = 3'h5 == state ? _GEN_9729 : valid_1_97; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10761 = 3'h5 == state ? _GEN_9730 : valid_1_98; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10762 = 3'h5 == state ? _GEN_9731 : valid_1_99; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10763 = 3'h5 == state ? _GEN_9732 : valid_1_100; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10764 = 3'h5 == state ? _GEN_9733 : valid_1_101; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10765 = 3'h5 == state ? _GEN_9734 : valid_1_102; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10766 = 3'h5 == state ? _GEN_9735 : valid_1_103; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10767 = 3'h5 == state ? _GEN_9736 : valid_1_104; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10768 = 3'h5 == state ? _GEN_9737 : valid_1_105; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10769 = 3'h5 == state ? _GEN_9738 : valid_1_106; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10770 = 3'h5 == state ? _GEN_9739 : valid_1_107; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10771 = 3'h5 == state ? _GEN_9740 : valid_1_108; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10772 = 3'h5 == state ? _GEN_9741 : valid_1_109; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10773 = 3'h5 == state ? _GEN_9742 : valid_1_110; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10774 = 3'h5 == state ? _GEN_9743 : valid_1_111; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10775 = 3'h5 == state ? _GEN_9744 : valid_1_112; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10776 = 3'h5 == state ? _GEN_9745 : valid_1_113; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10777 = 3'h5 == state ? _GEN_9746 : valid_1_114; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10778 = 3'h5 == state ? _GEN_9747 : valid_1_115; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10779 = 3'h5 == state ? _GEN_9748 : valid_1_116; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10780 = 3'h5 == state ? _GEN_9749 : valid_1_117; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10781 = 3'h5 == state ? _GEN_9750 : valid_1_118; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10782 = 3'h5 == state ? _GEN_9751 : valid_1_119; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10783 = 3'h5 == state ? _GEN_9752 : valid_1_120; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10784 = 3'h5 == state ? _GEN_9753 : valid_1_121; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10785 = 3'h5 == state ? _GEN_9754 : valid_1_122; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10786 = 3'h5 == state ? _GEN_9755 : valid_1_123; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10787 = 3'h5 == state ? _GEN_9756 : valid_1_124; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10788 = 3'h5 == state ? _GEN_9757 : valid_1_125; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10789 = 3'h5 == state ? _GEN_9758 : valid_1_126; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_10790 = 3'h5 == state ? _GEN_9759 : valid_1_127; // @[d_cache.scala 78:18 23:26]
  wire [63:0] _GEN_10791 = 3'h5 == state ? _GEN_9760 : write_back_data; // @[d_cache.scala 78:18 29:34]
  wire [41:0] _GEN_10792 = 3'h5 == state ? _GEN_9761 : {{10'd0}, write_back_addr}; // @[d_cache.scala 78:18 30:34]
  wire  _GEN_10793 = 3'h5 == state ? _GEN_9762 : dirty_0_0; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10794 = 3'h5 == state ? _GEN_9763 : dirty_0_1; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10795 = 3'h5 == state ? _GEN_9764 : dirty_0_2; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10796 = 3'h5 == state ? _GEN_9765 : dirty_0_3; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10797 = 3'h5 == state ? _GEN_9766 : dirty_0_4; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10798 = 3'h5 == state ? _GEN_9767 : dirty_0_5; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10799 = 3'h5 == state ? _GEN_9768 : dirty_0_6; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10800 = 3'h5 == state ? _GEN_9769 : dirty_0_7; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10801 = 3'h5 == state ? _GEN_9770 : dirty_0_8; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10802 = 3'h5 == state ? _GEN_9771 : dirty_0_9; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10803 = 3'h5 == state ? _GEN_9772 : dirty_0_10; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10804 = 3'h5 == state ? _GEN_9773 : dirty_0_11; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10805 = 3'h5 == state ? _GEN_9774 : dirty_0_12; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10806 = 3'h5 == state ? _GEN_9775 : dirty_0_13; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10807 = 3'h5 == state ? _GEN_9776 : dirty_0_14; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10808 = 3'h5 == state ? _GEN_9777 : dirty_0_15; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10809 = 3'h5 == state ? _GEN_9778 : dirty_0_16; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10810 = 3'h5 == state ? _GEN_9779 : dirty_0_17; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10811 = 3'h5 == state ? _GEN_9780 : dirty_0_18; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10812 = 3'h5 == state ? _GEN_9781 : dirty_0_19; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10813 = 3'h5 == state ? _GEN_9782 : dirty_0_20; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10814 = 3'h5 == state ? _GEN_9783 : dirty_0_21; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10815 = 3'h5 == state ? _GEN_9784 : dirty_0_22; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10816 = 3'h5 == state ? _GEN_9785 : dirty_0_23; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10817 = 3'h5 == state ? _GEN_9786 : dirty_0_24; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10818 = 3'h5 == state ? _GEN_9787 : dirty_0_25; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10819 = 3'h5 == state ? _GEN_9788 : dirty_0_26; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10820 = 3'h5 == state ? _GEN_9789 : dirty_0_27; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10821 = 3'h5 == state ? _GEN_9790 : dirty_0_28; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10822 = 3'h5 == state ? _GEN_9791 : dirty_0_29; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10823 = 3'h5 == state ? _GEN_9792 : dirty_0_30; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10824 = 3'h5 == state ? _GEN_9793 : dirty_0_31; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10825 = 3'h5 == state ? _GEN_9794 : dirty_0_32; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10826 = 3'h5 == state ? _GEN_9795 : dirty_0_33; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10827 = 3'h5 == state ? _GEN_9796 : dirty_0_34; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10828 = 3'h5 == state ? _GEN_9797 : dirty_0_35; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10829 = 3'h5 == state ? _GEN_9798 : dirty_0_36; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10830 = 3'h5 == state ? _GEN_9799 : dirty_0_37; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10831 = 3'h5 == state ? _GEN_9800 : dirty_0_38; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10832 = 3'h5 == state ? _GEN_9801 : dirty_0_39; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10833 = 3'h5 == state ? _GEN_9802 : dirty_0_40; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10834 = 3'h5 == state ? _GEN_9803 : dirty_0_41; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10835 = 3'h5 == state ? _GEN_9804 : dirty_0_42; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10836 = 3'h5 == state ? _GEN_9805 : dirty_0_43; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10837 = 3'h5 == state ? _GEN_9806 : dirty_0_44; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10838 = 3'h5 == state ? _GEN_9807 : dirty_0_45; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10839 = 3'h5 == state ? _GEN_9808 : dirty_0_46; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10840 = 3'h5 == state ? _GEN_9809 : dirty_0_47; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10841 = 3'h5 == state ? _GEN_9810 : dirty_0_48; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10842 = 3'h5 == state ? _GEN_9811 : dirty_0_49; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10843 = 3'h5 == state ? _GEN_9812 : dirty_0_50; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10844 = 3'h5 == state ? _GEN_9813 : dirty_0_51; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10845 = 3'h5 == state ? _GEN_9814 : dirty_0_52; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10846 = 3'h5 == state ? _GEN_9815 : dirty_0_53; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10847 = 3'h5 == state ? _GEN_9816 : dirty_0_54; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10848 = 3'h5 == state ? _GEN_9817 : dirty_0_55; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10849 = 3'h5 == state ? _GEN_9818 : dirty_0_56; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10850 = 3'h5 == state ? _GEN_9819 : dirty_0_57; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10851 = 3'h5 == state ? _GEN_9820 : dirty_0_58; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10852 = 3'h5 == state ? _GEN_9821 : dirty_0_59; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10853 = 3'h5 == state ? _GEN_9822 : dirty_0_60; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10854 = 3'h5 == state ? _GEN_9823 : dirty_0_61; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10855 = 3'h5 == state ? _GEN_9824 : dirty_0_62; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10856 = 3'h5 == state ? _GEN_9825 : dirty_0_63; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10857 = 3'h5 == state ? _GEN_9826 : dirty_0_64; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10858 = 3'h5 == state ? _GEN_9827 : dirty_0_65; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10859 = 3'h5 == state ? _GEN_9828 : dirty_0_66; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10860 = 3'h5 == state ? _GEN_9829 : dirty_0_67; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10861 = 3'h5 == state ? _GEN_9830 : dirty_0_68; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10862 = 3'h5 == state ? _GEN_9831 : dirty_0_69; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10863 = 3'h5 == state ? _GEN_9832 : dirty_0_70; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10864 = 3'h5 == state ? _GEN_9833 : dirty_0_71; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10865 = 3'h5 == state ? _GEN_9834 : dirty_0_72; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10866 = 3'h5 == state ? _GEN_9835 : dirty_0_73; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10867 = 3'h5 == state ? _GEN_9836 : dirty_0_74; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10868 = 3'h5 == state ? _GEN_9837 : dirty_0_75; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10869 = 3'h5 == state ? _GEN_9838 : dirty_0_76; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10870 = 3'h5 == state ? _GEN_9839 : dirty_0_77; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10871 = 3'h5 == state ? _GEN_9840 : dirty_0_78; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10872 = 3'h5 == state ? _GEN_9841 : dirty_0_79; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10873 = 3'h5 == state ? _GEN_9842 : dirty_0_80; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10874 = 3'h5 == state ? _GEN_9843 : dirty_0_81; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10875 = 3'h5 == state ? _GEN_9844 : dirty_0_82; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10876 = 3'h5 == state ? _GEN_9845 : dirty_0_83; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10877 = 3'h5 == state ? _GEN_9846 : dirty_0_84; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10878 = 3'h5 == state ? _GEN_9847 : dirty_0_85; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10879 = 3'h5 == state ? _GEN_9848 : dirty_0_86; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10880 = 3'h5 == state ? _GEN_9849 : dirty_0_87; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10881 = 3'h5 == state ? _GEN_9850 : dirty_0_88; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10882 = 3'h5 == state ? _GEN_9851 : dirty_0_89; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10883 = 3'h5 == state ? _GEN_9852 : dirty_0_90; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10884 = 3'h5 == state ? _GEN_9853 : dirty_0_91; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10885 = 3'h5 == state ? _GEN_9854 : dirty_0_92; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10886 = 3'h5 == state ? _GEN_9855 : dirty_0_93; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10887 = 3'h5 == state ? _GEN_9856 : dirty_0_94; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10888 = 3'h5 == state ? _GEN_9857 : dirty_0_95; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10889 = 3'h5 == state ? _GEN_9858 : dirty_0_96; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10890 = 3'h5 == state ? _GEN_9859 : dirty_0_97; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10891 = 3'h5 == state ? _GEN_9860 : dirty_0_98; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10892 = 3'h5 == state ? _GEN_9861 : dirty_0_99; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10893 = 3'h5 == state ? _GEN_9862 : dirty_0_100; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10894 = 3'h5 == state ? _GEN_9863 : dirty_0_101; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10895 = 3'h5 == state ? _GEN_9864 : dirty_0_102; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10896 = 3'h5 == state ? _GEN_9865 : dirty_0_103; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10897 = 3'h5 == state ? _GEN_9866 : dirty_0_104; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10898 = 3'h5 == state ? _GEN_9867 : dirty_0_105; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10899 = 3'h5 == state ? _GEN_9868 : dirty_0_106; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10900 = 3'h5 == state ? _GEN_9869 : dirty_0_107; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10901 = 3'h5 == state ? _GEN_9870 : dirty_0_108; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10902 = 3'h5 == state ? _GEN_9871 : dirty_0_109; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10903 = 3'h5 == state ? _GEN_9872 : dirty_0_110; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10904 = 3'h5 == state ? _GEN_9873 : dirty_0_111; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10905 = 3'h5 == state ? _GEN_9874 : dirty_0_112; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10906 = 3'h5 == state ? _GEN_9875 : dirty_0_113; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10907 = 3'h5 == state ? _GEN_9876 : dirty_0_114; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10908 = 3'h5 == state ? _GEN_9877 : dirty_0_115; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10909 = 3'h5 == state ? _GEN_9878 : dirty_0_116; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10910 = 3'h5 == state ? _GEN_9879 : dirty_0_117; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10911 = 3'h5 == state ? _GEN_9880 : dirty_0_118; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10912 = 3'h5 == state ? _GEN_9881 : dirty_0_119; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10913 = 3'h5 == state ? _GEN_9882 : dirty_0_120; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10914 = 3'h5 == state ? _GEN_9883 : dirty_0_121; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10915 = 3'h5 == state ? _GEN_9884 : dirty_0_122; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10916 = 3'h5 == state ? _GEN_9885 : dirty_0_123; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10917 = 3'h5 == state ? _GEN_9886 : dirty_0_124; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10918 = 3'h5 == state ? _GEN_9887 : dirty_0_125; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10919 = 3'h5 == state ? _GEN_9888 : dirty_0_126; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10920 = 3'h5 == state ? _GEN_9889 : dirty_0_127; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_10921 = 3'h5 == state ? _GEN_9890 : dirty_1_0; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10922 = 3'h5 == state ? _GEN_9891 : dirty_1_1; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10923 = 3'h5 == state ? _GEN_9892 : dirty_1_2; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10924 = 3'h5 == state ? _GEN_9893 : dirty_1_3; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10925 = 3'h5 == state ? _GEN_9894 : dirty_1_4; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10926 = 3'h5 == state ? _GEN_9895 : dirty_1_5; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10927 = 3'h5 == state ? _GEN_9896 : dirty_1_6; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10928 = 3'h5 == state ? _GEN_9897 : dirty_1_7; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10929 = 3'h5 == state ? _GEN_9898 : dirty_1_8; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10930 = 3'h5 == state ? _GEN_9899 : dirty_1_9; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10931 = 3'h5 == state ? _GEN_9900 : dirty_1_10; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10932 = 3'h5 == state ? _GEN_9901 : dirty_1_11; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10933 = 3'h5 == state ? _GEN_9902 : dirty_1_12; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10934 = 3'h5 == state ? _GEN_9903 : dirty_1_13; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10935 = 3'h5 == state ? _GEN_9904 : dirty_1_14; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10936 = 3'h5 == state ? _GEN_9905 : dirty_1_15; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10937 = 3'h5 == state ? _GEN_9906 : dirty_1_16; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10938 = 3'h5 == state ? _GEN_9907 : dirty_1_17; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10939 = 3'h5 == state ? _GEN_9908 : dirty_1_18; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10940 = 3'h5 == state ? _GEN_9909 : dirty_1_19; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10941 = 3'h5 == state ? _GEN_9910 : dirty_1_20; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10942 = 3'h5 == state ? _GEN_9911 : dirty_1_21; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10943 = 3'h5 == state ? _GEN_9912 : dirty_1_22; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10944 = 3'h5 == state ? _GEN_9913 : dirty_1_23; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10945 = 3'h5 == state ? _GEN_9914 : dirty_1_24; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10946 = 3'h5 == state ? _GEN_9915 : dirty_1_25; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10947 = 3'h5 == state ? _GEN_9916 : dirty_1_26; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10948 = 3'h5 == state ? _GEN_9917 : dirty_1_27; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10949 = 3'h5 == state ? _GEN_9918 : dirty_1_28; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10950 = 3'h5 == state ? _GEN_9919 : dirty_1_29; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10951 = 3'h5 == state ? _GEN_9920 : dirty_1_30; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10952 = 3'h5 == state ? _GEN_9921 : dirty_1_31; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10953 = 3'h5 == state ? _GEN_9922 : dirty_1_32; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10954 = 3'h5 == state ? _GEN_9923 : dirty_1_33; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10955 = 3'h5 == state ? _GEN_9924 : dirty_1_34; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10956 = 3'h5 == state ? _GEN_9925 : dirty_1_35; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10957 = 3'h5 == state ? _GEN_9926 : dirty_1_36; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10958 = 3'h5 == state ? _GEN_9927 : dirty_1_37; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10959 = 3'h5 == state ? _GEN_9928 : dirty_1_38; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10960 = 3'h5 == state ? _GEN_9929 : dirty_1_39; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10961 = 3'h5 == state ? _GEN_9930 : dirty_1_40; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10962 = 3'h5 == state ? _GEN_9931 : dirty_1_41; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10963 = 3'h5 == state ? _GEN_9932 : dirty_1_42; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10964 = 3'h5 == state ? _GEN_9933 : dirty_1_43; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10965 = 3'h5 == state ? _GEN_9934 : dirty_1_44; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10966 = 3'h5 == state ? _GEN_9935 : dirty_1_45; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10967 = 3'h5 == state ? _GEN_9936 : dirty_1_46; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10968 = 3'h5 == state ? _GEN_9937 : dirty_1_47; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10969 = 3'h5 == state ? _GEN_9938 : dirty_1_48; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10970 = 3'h5 == state ? _GEN_9939 : dirty_1_49; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10971 = 3'h5 == state ? _GEN_9940 : dirty_1_50; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10972 = 3'h5 == state ? _GEN_9941 : dirty_1_51; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10973 = 3'h5 == state ? _GEN_9942 : dirty_1_52; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10974 = 3'h5 == state ? _GEN_9943 : dirty_1_53; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10975 = 3'h5 == state ? _GEN_9944 : dirty_1_54; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10976 = 3'h5 == state ? _GEN_9945 : dirty_1_55; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10977 = 3'h5 == state ? _GEN_9946 : dirty_1_56; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10978 = 3'h5 == state ? _GEN_9947 : dirty_1_57; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10979 = 3'h5 == state ? _GEN_9948 : dirty_1_58; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10980 = 3'h5 == state ? _GEN_9949 : dirty_1_59; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10981 = 3'h5 == state ? _GEN_9950 : dirty_1_60; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10982 = 3'h5 == state ? _GEN_9951 : dirty_1_61; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10983 = 3'h5 == state ? _GEN_9952 : dirty_1_62; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10984 = 3'h5 == state ? _GEN_9953 : dirty_1_63; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10985 = 3'h5 == state ? _GEN_9954 : dirty_1_64; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10986 = 3'h5 == state ? _GEN_9955 : dirty_1_65; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10987 = 3'h5 == state ? _GEN_9956 : dirty_1_66; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10988 = 3'h5 == state ? _GEN_9957 : dirty_1_67; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10989 = 3'h5 == state ? _GEN_9958 : dirty_1_68; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10990 = 3'h5 == state ? _GEN_9959 : dirty_1_69; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10991 = 3'h5 == state ? _GEN_9960 : dirty_1_70; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10992 = 3'h5 == state ? _GEN_9961 : dirty_1_71; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10993 = 3'h5 == state ? _GEN_9962 : dirty_1_72; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10994 = 3'h5 == state ? _GEN_9963 : dirty_1_73; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10995 = 3'h5 == state ? _GEN_9964 : dirty_1_74; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10996 = 3'h5 == state ? _GEN_9965 : dirty_1_75; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10997 = 3'h5 == state ? _GEN_9966 : dirty_1_76; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10998 = 3'h5 == state ? _GEN_9967 : dirty_1_77; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_10999 = 3'h5 == state ? _GEN_9968 : dirty_1_78; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11000 = 3'h5 == state ? _GEN_9969 : dirty_1_79; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11001 = 3'h5 == state ? _GEN_9970 : dirty_1_80; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11002 = 3'h5 == state ? _GEN_9971 : dirty_1_81; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11003 = 3'h5 == state ? _GEN_9972 : dirty_1_82; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11004 = 3'h5 == state ? _GEN_9973 : dirty_1_83; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11005 = 3'h5 == state ? _GEN_9974 : dirty_1_84; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11006 = 3'h5 == state ? _GEN_9975 : dirty_1_85; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11007 = 3'h5 == state ? _GEN_9976 : dirty_1_86; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11008 = 3'h5 == state ? _GEN_9977 : dirty_1_87; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11009 = 3'h5 == state ? _GEN_9978 : dirty_1_88; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11010 = 3'h5 == state ? _GEN_9979 : dirty_1_89; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11011 = 3'h5 == state ? _GEN_9980 : dirty_1_90; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11012 = 3'h5 == state ? _GEN_9981 : dirty_1_91; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11013 = 3'h5 == state ? _GEN_9982 : dirty_1_92; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11014 = 3'h5 == state ? _GEN_9983 : dirty_1_93; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11015 = 3'h5 == state ? _GEN_9984 : dirty_1_94; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11016 = 3'h5 == state ? _GEN_9985 : dirty_1_95; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11017 = 3'h5 == state ? _GEN_9986 : dirty_1_96; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11018 = 3'h5 == state ? _GEN_9987 : dirty_1_97; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11019 = 3'h5 == state ? _GEN_9988 : dirty_1_98; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11020 = 3'h5 == state ? _GEN_9989 : dirty_1_99; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11021 = 3'h5 == state ? _GEN_9990 : dirty_1_100; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11022 = 3'h5 == state ? _GEN_9991 : dirty_1_101; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11023 = 3'h5 == state ? _GEN_9992 : dirty_1_102; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11024 = 3'h5 == state ? _GEN_9993 : dirty_1_103; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11025 = 3'h5 == state ? _GEN_9994 : dirty_1_104; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11026 = 3'h5 == state ? _GEN_9995 : dirty_1_105; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11027 = 3'h5 == state ? _GEN_9996 : dirty_1_106; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11028 = 3'h5 == state ? _GEN_9997 : dirty_1_107; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11029 = 3'h5 == state ? _GEN_9998 : dirty_1_108; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11030 = 3'h5 == state ? _GEN_9999 : dirty_1_109; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11031 = 3'h5 == state ? _GEN_10000 : dirty_1_110; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11032 = 3'h5 == state ? _GEN_10001 : dirty_1_111; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11033 = 3'h5 == state ? _GEN_10002 : dirty_1_112; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11034 = 3'h5 == state ? _GEN_10003 : dirty_1_113; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11035 = 3'h5 == state ? _GEN_10004 : dirty_1_114; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11036 = 3'h5 == state ? _GEN_10005 : dirty_1_115; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11037 = 3'h5 == state ? _GEN_10006 : dirty_1_116; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11038 = 3'h5 == state ? _GEN_10007 : dirty_1_117; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11039 = 3'h5 == state ? _GEN_10008 : dirty_1_118; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11040 = 3'h5 == state ? _GEN_10009 : dirty_1_119; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11041 = 3'h5 == state ? _GEN_10010 : dirty_1_120; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11042 = 3'h5 == state ? _GEN_10011 : dirty_1_121; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11043 = 3'h5 == state ? _GEN_10012 : dirty_1_122; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11044 = 3'h5 == state ? _GEN_10013 : dirty_1_123; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11045 = 3'h5 == state ? _GEN_10014 : dirty_1_124; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11046 = 3'h5 == state ? _GEN_10015 : dirty_1_125; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11047 = 3'h5 == state ? _GEN_10016 : dirty_1_126; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11048 = 3'h5 == state ? _GEN_10017 : dirty_1_127; // @[d_cache.scala 78:18 25:26]
  wire [2:0] _GEN_11049 = 3'h4 == state ? _GEN_2573 : _GEN_10021; // @[d_cache.scala 78:18]
  wire [63:0] _GEN_11050 = 3'h4 == state ? ram_0_0 : _GEN_10022; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11051 = 3'h4 == state ? ram_0_1 : _GEN_10023; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11052 = 3'h4 == state ? ram_0_2 : _GEN_10024; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11053 = 3'h4 == state ? ram_0_3 : _GEN_10025; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11054 = 3'h4 == state ? ram_0_4 : _GEN_10026; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11055 = 3'h4 == state ? ram_0_5 : _GEN_10027; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11056 = 3'h4 == state ? ram_0_6 : _GEN_10028; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11057 = 3'h4 == state ? ram_0_7 : _GEN_10029; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11058 = 3'h4 == state ? ram_0_8 : _GEN_10030; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11059 = 3'h4 == state ? ram_0_9 : _GEN_10031; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11060 = 3'h4 == state ? ram_0_10 : _GEN_10032; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11061 = 3'h4 == state ? ram_0_11 : _GEN_10033; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11062 = 3'h4 == state ? ram_0_12 : _GEN_10034; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11063 = 3'h4 == state ? ram_0_13 : _GEN_10035; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11064 = 3'h4 == state ? ram_0_14 : _GEN_10036; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11065 = 3'h4 == state ? ram_0_15 : _GEN_10037; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11066 = 3'h4 == state ? ram_0_16 : _GEN_10038; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11067 = 3'h4 == state ? ram_0_17 : _GEN_10039; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11068 = 3'h4 == state ? ram_0_18 : _GEN_10040; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11069 = 3'h4 == state ? ram_0_19 : _GEN_10041; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11070 = 3'h4 == state ? ram_0_20 : _GEN_10042; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11071 = 3'h4 == state ? ram_0_21 : _GEN_10043; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11072 = 3'h4 == state ? ram_0_22 : _GEN_10044; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11073 = 3'h4 == state ? ram_0_23 : _GEN_10045; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11074 = 3'h4 == state ? ram_0_24 : _GEN_10046; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11075 = 3'h4 == state ? ram_0_25 : _GEN_10047; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11076 = 3'h4 == state ? ram_0_26 : _GEN_10048; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11077 = 3'h4 == state ? ram_0_27 : _GEN_10049; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11078 = 3'h4 == state ? ram_0_28 : _GEN_10050; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11079 = 3'h4 == state ? ram_0_29 : _GEN_10051; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11080 = 3'h4 == state ? ram_0_30 : _GEN_10052; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11081 = 3'h4 == state ? ram_0_31 : _GEN_10053; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11082 = 3'h4 == state ? ram_0_32 : _GEN_10054; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11083 = 3'h4 == state ? ram_0_33 : _GEN_10055; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11084 = 3'h4 == state ? ram_0_34 : _GEN_10056; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11085 = 3'h4 == state ? ram_0_35 : _GEN_10057; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11086 = 3'h4 == state ? ram_0_36 : _GEN_10058; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11087 = 3'h4 == state ? ram_0_37 : _GEN_10059; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11088 = 3'h4 == state ? ram_0_38 : _GEN_10060; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11089 = 3'h4 == state ? ram_0_39 : _GEN_10061; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11090 = 3'h4 == state ? ram_0_40 : _GEN_10062; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11091 = 3'h4 == state ? ram_0_41 : _GEN_10063; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11092 = 3'h4 == state ? ram_0_42 : _GEN_10064; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11093 = 3'h4 == state ? ram_0_43 : _GEN_10065; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11094 = 3'h4 == state ? ram_0_44 : _GEN_10066; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11095 = 3'h4 == state ? ram_0_45 : _GEN_10067; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11096 = 3'h4 == state ? ram_0_46 : _GEN_10068; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11097 = 3'h4 == state ? ram_0_47 : _GEN_10069; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11098 = 3'h4 == state ? ram_0_48 : _GEN_10070; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11099 = 3'h4 == state ? ram_0_49 : _GEN_10071; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11100 = 3'h4 == state ? ram_0_50 : _GEN_10072; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11101 = 3'h4 == state ? ram_0_51 : _GEN_10073; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11102 = 3'h4 == state ? ram_0_52 : _GEN_10074; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11103 = 3'h4 == state ? ram_0_53 : _GEN_10075; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11104 = 3'h4 == state ? ram_0_54 : _GEN_10076; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11105 = 3'h4 == state ? ram_0_55 : _GEN_10077; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11106 = 3'h4 == state ? ram_0_56 : _GEN_10078; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11107 = 3'h4 == state ? ram_0_57 : _GEN_10079; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11108 = 3'h4 == state ? ram_0_58 : _GEN_10080; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11109 = 3'h4 == state ? ram_0_59 : _GEN_10081; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11110 = 3'h4 == state ? ram_0_60 : _GEN_10082; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11111 = 3'h4 == state ? ram_0_61 : _GEN_10083; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11112 = 3'h4 == state ? ram_0_62 : _GEN_10084; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11113 = 3'h4 == state ? ram_0_63 : _GEN_10085; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11114 = 3'h4 == state ? ram_0_64 : _GEN_10086; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11115 = 3'h4 == state ? ram_0_65 : _GEN_10087; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11116 = 3'h4 == state ? ram_0_66 : _GEN_10088; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11117 = 3'h4 == state ? ram_0_67 : _GEN_10089; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11118 = 3'h4 == state ? ram_0_68 : _GEN_10090; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11119 = 3'h4 == state ? ram_0_69 : _GEN_10091; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11120 = 3'h4 == state ? ram_0_70 : _GEN_10092; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11121 = 3'h4 == state ? ram_0_71 : _GEN_10093; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11122 = 3'h4 == state ? ram_0_72 : _GEN_10094; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11123 = 3'h4 == state ? ram_0_73 : _GEN_10095; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11124 = 3'h4 == state ? ram_0_74 : _GEN_10096; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11125 = 3'h4 == state ? ram_0_75 : _GEN_10097; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11126 = 3'h4 == state ? ram_0_76 : _GEN_10098; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11127 = 3'h4 == state ? ram_0_77 : _GEN_10099; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11128 = 3'h4 == state ? ram_0_78 : _GEN_10100; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11129 = 3'h4 == state ? ram_0_79 : _GEN_10101; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11130 = 3'h4 == state ? ram_0_80 : _GEN_10102; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11131 = 3'h4 == state ? ram_0_81 : _GEN_10103; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11132 = 3'h4 == state ? ram_0_82 : _GEN_10104; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11133 = 3'h4 == state ? ram_0_83 : _GEN_10105; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11134 = 3'h4 == state ? ram_0_84 : _GEN_10106; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11135 = 3'h4 == state ? ram_0_85 : _GEN_10107; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11136 = 3'h4 == state ? ram_0_86 : _GEN_10108; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11137 = 3'h4 == state ? ram_0_87 : _GEN_10109; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11138 = 3'h4 == state ? ram_0_88 : _GEN_10110; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11139 = 3'h4 == state ? ram_0_89 : _GEN_10111; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11140 = 3'h4 == state ? ram_0_90 : _GEN_10112; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11141 = 3'h4 == state ? ram_0_91 : _GEN_10113; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11142 = 3'h4 == state ? ram_0_92 : _GEN_10114; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11143 = 3'h4 == state ? ram_0_93 : _GEN_10115; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11144 = 3'h4 == state ? ram_0_94 : _GEN_10116; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11145 = 3'h4 == state ? ram_0_95 : _GEN_10117; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11146 = 3'h4 == state ? ram_0_96 : _GEN_10118; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11147 = 3'h4 == state ? ram_0_97 : _GEN_10119; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11148 = 3'h4 == state ? ram_0_98 : _GEN_10120; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11149 = 3'h4 == state ? ram_0_99 : _GEN_10121; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11150 = 3'h4 == state ? ram_0_100 : _GEN_10122; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11151 = 3'h4 == state ? ram_0_101 : _GEN_10123; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11152 = 3'h4 == state ? ram_0_102 : _GEN_10124; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11153 = 3'h4 == state ? ram_0_103 : _GEN_10125; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11154 = 3'h4 == state ? ram_0_104 : _GEN_10126; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11155 = 3'h4 == state ? ram_0_105 : _GEN_10127; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11156 = 3'h4 == state ? ram_0_106 : _GEN_10128; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11157 = 3'h4 == state ? ram_0_107 : _GEN_10129; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11158 = 3'h4 == state ? ram_0_108 : _GEN_10130; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11159 = 3'h4 == state ? ram_0_109 : _GEN_10131; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11160 = 3'h4 == state ? ram_0_110 : _GEN_10132; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11161 = 3'h4 == state ? ram_0_111 : _GEN_10133; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11162 = 3'h4 == state ? ram_0_112 : _GEN_10134; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11163 = 3'h4 == state ? ram_0_113 : _GEN_10135; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11164 = 3'h4 == state ? ram_0_114 : _GEN_10136; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11165 = 3'h4 == state ? ram_0_115 : _GEN_10137; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11166 = 3'h4 == state ? ram_0_116 : _GEN_10138; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11167 = 3'h4 == state ? ram_0_117 : _GEN_10139; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11168 = 3'h4 == state ? ram_0_118 : _GEN_10140; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11169 = 3'h4 == state ? ram_0_119 : _GEN_10141; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11170 = 3'h4 == state ? ram_0_120 : _GEN_10142; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11171 = 3'h4 == state ? ram_0_121 : _GEN_10143; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11172 = 3'h4 == state ? ram_0_122 : _GEN_10144; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11173 = 3'h4 == state ? ram_0_123 : _GEN_10145; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11174 = 3'h4 == state ? ram_0_124 : _GEN_10146; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11175 = 3'h4 == state ? ram_0_125 : _GEN_10147; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11176 = 3'h4 == state ? ram_0_126 : _GEN_10148; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_11177 = 3'h4 == state ? ram_0_127 : _GEN_10149; // @[d_cache.scala 78:18 18:24]
  wire [31:0] _GEN_11178 = 3'h4 == state ? tag_0_0 : _GEN_10150; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11179 = 3'h4 == state ? tag_0_1 : _GEN_10151; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11180 = 3'h4 == state ? tag_0_2 : _GEN_10152; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11181 = 3'h4 == state ? tag_0_3 : _GEN_10153; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11182 = 3'h4 == state ? tag_0_4 : _GEN_10154; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11183 = 3'h4 == state ? tag_0_5 : _GEN_10155; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11184 = 3'h4 == state ? tag_0_6 : _GEN_10156; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11185 = 3'h4 == state ? tag_0_7 : _GEN_10157; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11186 = 3'h4 == state ? tag_0_8 : _GEN_10158; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11187 = 3'h4 == state ? tag_0_9 : _GEN_10159; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11188 = 3'h4 == state ? tag_0_10 : _GEN_10160; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11189 = 3'h4 == state ? tag_0_11 : _GEN_10161; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11190 = 3'h4 == state ? tag_0_12 : _GEN_10162; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11191 = 3'h4 == state ? tag_0_13 : _GEN_10163; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11192 = 3'h4 == state ? tag_0_14 : _GEN_10164; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11193 = 3'h4 == state ? tag_0_15 : _GEN_10165; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11194 = 3'h4 == state ? tag_0_16 : _GEN_10166; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11195 = 3'h4 == state ? tag_0_17 : _GEN_10167; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11196 = 3'h4 == state ? tag_0_18 : _GEN_10168; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11197 = 3'h4 == state ? tag_0_19 : _GEN_10169; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11198 = 3'h4 == state ? tag_0_20 : _GEN_10170; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11199 = 3'h4 == state ? tag_0_21 : _GEN_10171; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11200 = 3'h4 == state ? tag_0_22 : _GEN_10172; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11201 = 3'h4 == state ? tag_0_23 : _GEN_10173; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11202 = 3'h4 == state ? tag_0_24 : _GEN_10174; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11203 = 3'h4 == state ? tag_0_25 : _GEN_10175; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11204 = 3'h4 == state ? tag_0_26 : _GEN_10176; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11205 = 3'h4 == state ? tag_0_27 : _GEN_10177; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11206 = 3'h4 == state ? tag_0_28 : _GEN_10178; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11207 = 3'h4 == state ? tag_0_29 : _GEN_10179; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11208 = 3'h4 == state ? tag_0_30 : _GEN_10180; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11209 = 3'h4 == state ? tag_0_31 : _GEN_10181; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11210 = 3'h4 == state ? tag_0_32 : _GEN_10182; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11211 = 3'h4 == state ? tag_0_33 : _GEN_10183; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11212 = 3'h4 == state ? tag_0_34 : _GEN_10184; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11213 = 3'h4 == state ? tag_0_35 : _GEN_10185; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11214 = 3'h4 == state ? tag_0_36 : _GEN_10186; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11215 = 3'h4 == state ? tag_0_37 : _GEN_10187; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11216 = 3'h4 == state ? tag_0_38 : _GEN_10188; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11217 = 3'h4 == state ? tag_0_39 : _GEN_10189; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11218 = 3'h4 == state ? tag_0_40 : _GEN_10190; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11219 = 3'h4 == state ? tag_0_41 : _GEN_10191; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11220 = 3'h4 == state ? tag_0_42 : _GEN_10192; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11221 = 3'h4 == state ? tag_0_43 : _GEN_10193; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11222 = 3'h4 == state ? tag_0_44 : _GEN_10194; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11223 = 3'h4 == state ? tag_0_45 : _GEN_10195; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11224 = 3'h4 == state ? tag_0_46 : _GEN_10196; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11225 = 3'h4 == state ? tag_0_47 : _GEN_10197; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11226 = 3'h4 == state ? tag_0_48 : _GEN_10198; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11227 = 3'h4 == state ? tag_0_49 : _GEN_10199; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11228 = 3'h4 == state ? tag_0_50 : _GEN_10200; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11229 = 3'h4 == state ? tag_0_51 : _GEN_10201; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11230 = 3'h4 == state ? tag_0_52 : _GEN_10202; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11231 = 3'h4 == state ? tag_0_53 : _GEN_10203; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11232 = 3'h4 == state ? tag_0_54 : _GEN_10204; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11233 = 3'h4 == state ? tag_0_55 : _GEN_10205; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11234 = 3'h4 == state ? tag_0_56 : _GEN_10206; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11235 = 3'h4 == state ? tag_0_57 : _GEN_10207; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11236 = 3'h4 == state ? tag_0_58 : _GEN_10208; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11237 = 3'h4 == state ? tag_0_59 : _GEN_10209; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11238 = 3'h4 == state ? tag_0_60 : _GEN_10210; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11239 = 3'h4 == state ? tag_0_61 : _GEN_10211; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11240 = 3'h4 == state ? tag_0_62 : _GEN_10212; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11241 = 3'h4 == state ? tag_0_63 : _GEN_10213; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11242 = 3'h4 == state ? tag_0_64 : _GEN_10214; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11243 = 3'h4 == state ? tag_0_65 : _GEN_10215; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11244 = 3'h4 == state ? tag_0_66 : _GEN_10216; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11245 = 3'h4 == state ? tag_0_67 : _GEN_10217; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11246 = 3'h4 == state ? tag_0_68 : _GEN_10218; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11247 = 3'h4 == state ? tag_0_69 : _GEN_10219; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11248 = 3'h4 == state ? tag_0_70 : _GEN_10220; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11249 = 3'h4 == state ? tag_0_71 : _GEN_10221; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11250 = 3'h4 == state ? tag_0_72 : _GEN_10222; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11251 = 3'h4 == state ? tag_0_73 : _GEN_10223; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11252 = 3'h4 == state ? tag_0_74 : _GEN_10224; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11253 = 3'h4 == state ? tag_0_75 : _GEN_10225; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11254 = 3'h4 == state ? tag_0_76 : _GEN_10226; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11255 = 3'h4 == state ? tag_0_77 : _GEN_10227; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11256 = 3'h4 == state ? tag_0_78 : _GEN_10228; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11257 = 3'h4 == state ? tag_0_79 : _GEN_10229; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11258 = 3'h4 == state ? tag_0_80 : _GEN_10230; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11259 = 3'h4 == state ? tag_0_81 : _GEN_10231; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11260 = 3'h4 == state ? tag_0_82 : _GEN_10232; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11261 = 3'h4 == state ? tag_0_83 : _GEN_10233; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11262 = 3'h4 == state ? tag_0_84 : _GEN_10234; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11263 = 3'h4 == state ? tag_0_85 : _GEN_10235; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11264 = 3'h4 == state ? tag_0_86 : _GEN_10236; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11265 = 3'h4 == state ? tag_0_87 : _GEN_10237; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11266 = 3'h4 == state ? tag_0_88 : _GEN_10238; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11267 = 3'h4 == state ? tag_0_89 : _GEN_10239; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11268 = 3'h4 == state ? tag_0_90 : _GEN_10240; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11269 = 3'h4 == state ? tag_0_91 : _GEN_10241; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11270 = 3'h4 == state ? tag_0_92 : _GEN_10242; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11271 = 3'h4 == state ? tag_0_93 : _GEN_10243; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11272 = 3'h4 == state ? tag_0_94 : _GEN_10244; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11273 = 3'h4 == state ? tag_0_95 : _GEN_10245; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11274 = 3'h4 == state ? tag_0_96 : _GEN_10246; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11275 = 3'h4 == state ? tag_0_97 : _GEN_10247; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11276 = 3'h4 == state ? tag_0_98 : _GEN_10248; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11277 = 3'h4 == state ? tag_0_99 : _GEN_10249; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11278 = 3'h4 == state ? tag_0_100 : _GEN_10250; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11279 = 3'h4 == state ? tag_0_101 : _GEN_10251; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11280 = 3'h4 == state ? tag_0_102 : _GEN_10252; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11281 = 3'h4 == state ? tag_0_103 : _GEN_10253; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11282 = 3'h4 == state ? tag_0_104 : _GEN_10254; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11283 = 3'h4 == state ? tag_0_105 : _GEN_10255; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11284 = 3'h4 == state ? tag_0_106 : _GEN_10256; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11285 = 3'h4 == state ? tag_0_107 : _GEN_10257; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11286 = 3'h4 == state ? tag_0_108 : _GEN_10258; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11287 = 3'h4 == state ? tag_0_109 : _GEN_10259; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11288 = 3'h4 == state ? tag_0_110 : _GEN_10260; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11289 = 3'h4 == state ? tag_0_111 : _GEN_10261; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11290 = 3'h4 == state ? tag_0_112 : _GEN_10262; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11291 = 3'h4 == state ? tag_0_113 : _GEN_10263; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11292 = 3'h4 == state ? tag_0_114 : _GEN_10264; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11293 = 3'h4 == state ? tag_0_115 : _GEN_10265; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11294 = 3'h4 == state ? tag_0_116 : _GEN_10266; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11295 = 3'h4 == state ? tag_0_117 : _GEN_10267; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11296 = 3'h4 == state ? tag_0_118 : _GEN_10268; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11297 = 3'h4 == state ? tag_0_119 : _GEN_10269; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11298 = 3'h4 == state ? tag_0_120 : _GEN_10270; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11299 = 3'h4 == state ? tag_0_121 : _GEN_10271; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11300 = 3'h4 == state ? tag_0_122 : _GEN_10272; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11301 = 3'h4 == state ? tag_0_123 : _GEN_10273; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11302 = 3'h4 == state ? tag_0_124 : _GEN_10274; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11303 = 3'h4 == state ? tag_0_125 : _GEN_10275; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11304 = 3'h4 == state ? tag_0_126 : _GEN_10276; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_11305 = 3'h4 == state ? tag_0_127 : _GEN_10277; // @[d_cache.scala 78:18 20:24]
  wire  _GEN_11306 = 3'h4 == state ? valid_0_0 : _GEN_10278; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11307 = 3'h4 == state ? valid_0_1 : _GEN_10279; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11308 = 3'h4 == state ? valid_0_2 : _GEN_10280; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11309 = 3'h4 == state ? valid_0_3 : _GEN_10281; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11310 = 3'h4 == state ? valid_0_4 : _GEN_10282; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11311 = 3'h4 == state ? valid_0_5 : _GEN_10283; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11312 = 3'h4 == state ? valid_0_6 : _GEN_10284; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11313 = 3'h4 == state ? valid_0_7 : _GEN_10285; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11314 = 3'h4 == state ? valid_0_8 : _GEN_10286; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11315 = 3'h4 == state ? valid_0_9 : _GEN_10287; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11316 = 3'h4 == state ? valid_0_10 : _GEN_10288; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11317 = 3'h4 == state ? valid_0_11 : _GEN_10289; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11318 = 3'h4 == state ? valid_0_12 : _GEN_10290; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11319 = 3'h4 == state ? valid_0_13 : _GEN_10291; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11320 = 3'h4 == state ? valid_0_14 : _GEN_10292; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11321 = 3'h4 == state ? valid_0_15 : _GEN_10293; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11322 = 3'h4 == state ? valid_0_16 : _GEN_10294; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11323 = 3'h4 == state ? valid_0_17 : _GEN_10295; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11324 = 3'h4 == state ? valid_0_18 : _GEN_10296; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11325 = 3'h4 == state ? valid_0_19 : _GEN_10297; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11326 = 3'h4 == state ? valid_0_20 : _GEN_10298; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11327 = 3'h4 == state ? valid_0_21 : _GEN_10299; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11328 = 3'h4 == state ? valid_0_22 : _GEN_10300; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11329 = 3'h4 == state ? valid_0_23 : _GEN_10301; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11330 = 3'h4 == state ? valid_0_24 : _GEN_10302; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11331 = 3'h4 == state ? valid_0_25 : _GEN_10303; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11332 = 3'h4 == state ? valid_0_26 : _GEN_10304; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11333 = 3'h4 == state ? valid_0_27 : _GEN_10305; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11334 = 3'h4 == state ? valid_0_28 : _GEN_10306; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11335 = 3'h4 == state ? valid_0_29 : _GEN_10307; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11336 = 3'h4 == state ? valid_0_30 : _GEN_10308; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11337 = 3'h4 == state ? valid_0_31 : _GEN_10309; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11338 = 3'h4 == state ? valid_0_32 : _GEN_10310; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11339 = 3'h4 == state ? valid_0_33 : _GEN_10311; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11340 = 3'h4 == state ? valid_0_34 : _GEN_10312; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11341 = 3'h4 == state ? valid_0_35 : _GEN_10313; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11342 = 3'h4 == state ? valid_0_36 : _GEN_10314; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11343 = 3'h4 == state ? valid_0_37 : _GEN_10315; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11344 = 3'h4 == state ? valid_0_38 : _GEN_10316; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11345 = 3'h4 == state ? valid_0_39 : _GEN_10317; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11346 = 3'h4 == state ? valid_0_40 : _GEN_10318; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11347 = 3'h4 == state ? valid_0_41 : _GEN_10319; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11348 = 3'h4 == state ? valid_0_42 : _GEN_10320; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11349 = 3'h4 == state ? valid_0_43 : _GEN_10321; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11350 = 3'h4 == state ? valid_0_44 : _GEN_10322; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11351 = 3'h4 == state ? valid_0_45 : _GEN_10323; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11352 = 3'h4 == state ? valid_0_46 : _GEN_10324; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11353 = 3'h4 == state ? valid_0_47 : _GEN_10325; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11354 = 3'h4 == state ? valid_0_48 : _GEN_10326; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11355 = 3'h4 == state ? valid_0_49 : _GEN_10327; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11356 = 3'h4 == state ? valid_0_50 : _GEN_10328; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11357 = 3'h4 == state ? valid_0_51 : _GEN_10329; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11358 = 3'h4 == state ? valid_0_52 : _GEN_10330; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11359 = 3'h4 == state ? valid_0_53 : _GEN_10331; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11360 = 3'h4 == state ? valid_0_54 : _GEN_10332; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11361 = 3'h4 == state ? valid_0_55 : _GEN_10333; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11362 = 3'h4 == state ? valid_0_56 : _GEN_10334; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11363 = 3'h4 == state ? valid_0_57 : _GEN_10335; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11364 = 3'h4 == state ? valid_0_58 : _GEN_10336; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11365 = 3'h4 == state ? valid_0_59 : _GEN_10337; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11366 = 3'h4 == state ? valid_0_60 : _GEN_10338; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11367 = 3'h4 == state ? valid_0_61 : _GEN_10339; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11368 = 3'h4 == state ? valid_0_62 : _GEN_10340; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11369 = 3'h4 == state ? valid_0_63 : _GEN_10341; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11370 = 3'h4 == state ? valid_0_64 : _GEN_10342; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11371 = 3'h4 == state ? valid_0_65 : _GEN_10343; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11372 = 3'h4 == state ? valid_0_66 : _GEN_10344; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11373 = 3'h4 == state ? valid_0_67 : _GEN_10345; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11374 = 3'h4 == state ? valid_0_68 : _GEN_10346; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11375 = 3'h4 == state ? valid_0_69 : _GEN_10347; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11376 = 3'h4 == state ? valid_0_70 : _GEN_10348; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11377 = 3'h4 == state ? valid_0_71 : _GEN_10349; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11378 = 3'h4 == state ? valid_0_72 : _GEN_10350; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11379 = 3'h4 == state ? valid_0_73 : _GEN_10351; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11380 = 3'h4 == state ? valid_0_74 : _GEN_10352; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11381 = 3'h4 == state ? valid_0_75 : _GEN_10353; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11382 = 3'h4 == state ? valid_0_76 : _GEN_10354; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11383 = 3'h4 == state ? valid_0_77 : _GEN_10355; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11384 = 3'h4 == state ? valid_0_78 : _GEN_10356; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11385 = 3'h4 == state ? valid_0_79 : _GEN_10357; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11386 = 3'h4 == state ? valid_0_80 : _GEN_10358; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11387 = 3'h4 == state ? valid_0_81 : _GEN_10359; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11388 = 3'h4 == state ? valid_0_82 : _GEN_10360; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11389 = 3'h4 == state ? valid_0_83 : _GEN_10361; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11390 = 3'h4 == state ? valid_0_84 : _GEN_10362; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11391 = 3'h4 == state ? valid_0_85 : _GEN_10363; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11392 = 3'h4 == state ? valid_0_86 : _GEN_10364; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11393 = 3'h4 == state ? valid_0_87 : _GEN_10365; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11394 = 3'h4 == state ? valid_0_88 : _GEN_10366; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11395 = 3'h4 == state ? valid_0_89 : _GEN_10367; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11396 = 3'h4 == state ? valid_0_90 : _GEN_10368; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11397 = 3'h4 == state ? valid_0_91 : _GEN_10369; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11398 = 3'h4 == state ? valid_0_92 : _GEN_10370; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11399 = 3'h4 == state ? valid_0_93 : _GEN_10371; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11400 = 3'h4 == state ? valid_0_94 : _GEN_10372; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11401 = 3'h4 == state ? valid_0_95 : _GEN_10373; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11402 = 3'h4 == state ? valid_0_96 : _GEN_10374; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11403 = 3'h4 == state ? valid_0_97 : _GEN_10375; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11404 = 3'h4 == state ? valid_0_98 : _GEN_10376; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11405 = 3'h4 == state ? valid_0_99 : _GEN_10377; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11406 = 3'h4 == state ? valid_0_100 : _GEN_10378; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11407 = 3'h4 == state ? valid_0_101 : _GEN_10379; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11408 = 3'h4 == state ? valid_0_102 : _GEN_10380; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11409 = 3'h4 == state ? valid_0_103 : _GEN_10381; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11410 = 3'h4 == state ? valid_0_104 : _GEN_10382; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11411 = 3'h4 == state ? valid_0_105 : _GEN_10383; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11412 = 3'h4 == state ? valid_0_106 : _GEN_10384; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11413 = 3'h4 == state ? valid_0_107 : _GEN_10385; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11414 = 3'h4 == state ? valid_0_108 : _GEN_10386; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11415 = 3'h4 == state ? valid_0_109 : _GEN_10387; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11416 = 3'h4 == state ? valid_0_110 : _GEN_10388; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11417 = 3'h4 == state ? valid_0_111 : _GEN_10389; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11418 = 3'h4 == state ? valid_0_112 : _GEN_10390; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11419 = 3'h4 == state ? valid_0_113 : _GEN_10391; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11420 = 3'h4 == state ? valid_0_114 : _GEN_10392; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11421 = 3'h4 == state ? valid_0_115 : _GEN_10393; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11422 = 3'h4 == state ? valid_0_116 : _GEN_10394; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11423 = 3'h4 == state ? valid_0_117 : _GEN_10395; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11424 = 3'h4 == state ? valid_0_118 : _GEN_10396; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11425 = 3'h4 == state ? valid_0_119 : _GEN_10397; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11426 = 3'h4 == state ? valid_0_120 : _GEN_10398; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11427 = 3'h4 == state ? valid_0_121 : _GEN_10399; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11428 = 3'h4 == state ? valid_0_122 : _GEN_10400; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11429 = 3'h4 == state ? valid_0_123 : _GEN_10401; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11430 = 3'h4 == state ? valid_0_124 : _GEN_10402; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11431 = 3'h4 == state ? valid_0_125 : _GEN_10403; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11432 = 3'h4 == state ? valid_0_126 : _GEN_10404; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11433 = 3'h4 == state ? valid_0_127 : _GEN_10405; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_11434 = 3'h4 == state ? quene : _GEN_10406; // @[d_cache.scala 78:18 35:24]
  wire [63:0] _GEN_11435 = 3'h4 == state ? ram_1_0 : _GEN_10407; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11436 = 3'h4 == state ? ram_1_1 : _GEN_10408; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11437 = 3'h4 == state ? ram_1_2 : _GEN_10409; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11438 = 3'h4 == state ? ram_1_3 : _GEN_10410; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11439 = 3'h4 == state ? ram_1_4 : _GEN_10411; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11440 = 3'h4 == state ? ram_1_5 : _GEN_10412; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11441 = 3'h4 == state ? ram_1_6 : _GEN_10413; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11442 = 3'h4 == state ? ram_1_7 : _GEN_10414; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11443 = 3'h4 == state ? ram_1_8 : _GEN_10415; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11444 = 3'h4 == state ? ram_1_9 : _GEN_10416; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11445 = 3'h4 == state ? ram_1_10 : _GEN_10417; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11446 = 3'h4 == state ? ram_1_11 : _GEN_10418; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11447 = 3'h4 == state ? ram_1_12 : _GEN_10419; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11448 = 3'h4 == state ? ram_1_13 : _GEN_10420; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11449 = 3'h4 == state ? ram_1_14 : _GEN_10421; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11450 = 3'h4 == state ? ram_1_15 : _GEN_10422; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11451 = 3'h4 == state ? ram_1_16 : _GEN_10423; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11452 = 3'h4 == state ? ram_1_17 : _GEN_10424; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11453 = 3'h4 == state ? ram_1_18 : _GEN_10425; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11454 = 3'h4 == state ? ram_1_19 : _GEN_10426; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11455 = 3'h4 == state ? ram_1_20 : _GEN_10427; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11456 = 3'h4 == state ? ram_1_21 : _GEN_10428; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11457 = 3'h4 == state ? ram_1_22 : _GEN_10429; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11458 = 3'h4 == state ? ram_1_23 : _GEN_10430; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11459 = 3'h4 == state ? ram_1_24 : _GEN_10431; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11460 = 3'h4 == state ? ram_1_25 : _GEN_10432; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11461 = 3'h4 == state ? ram_1_26 : _GEN_10433; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11462 = 3'h4 == state ? ram_1_27 : _GEN_10434; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11463 = 3'h4 == state ? ram_1_28 : _GEN_10435; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11464 = 3'h4 == state ? ram_1_29 : _GEN_10436; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11465 = 3'h4 == state ? ram_1_30 : _GEN_10437; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11466 = 3'h4 == state ? ram_1_31 : _GEN_10438; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11467 = 3'h4 == state ? ram_1_32 : _GEN_10439; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11468 = 3'h4 == state ? ram_1_33 : _GEN_10440; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11469 = 3'h4 == state ? ram_1_34 : _GEN_10441; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11470 = 3'h4 == state ? ram_1_35 : _GEN_10442; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11471 = 3'h4 == state ? ram_1_36 : _GEN_10443; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11472 = 3'h4 == state ? ram_1_37 : _GEN_10444; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11473 = 3'h4 == state ? ram_1_38 : _GEN_10445; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11474 = 3'h4 == state ? ram_1_39 : _GEN_10446; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11475 = 3'h4 == state ? ram_1_40 : _GEN_10447; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11476 = 3'h4 == state ? ram_1_41 : _GEN_10448; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11477 = 3'h4 == state ? ram_1_42 : _GEN_10449; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11478 = 3'h4 == state ? ram_1_43 : _GEN_10450; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11479 = 3'h4 == state ? ram_1_44 : _GEN_10451; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11480 = 3'h4 == state ? ram_1_45 : _GEN_10452; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11481 = 3'h4 == state ? ram_1_46 : _GEN_10453; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11482 = 3'h4 == state ? ram_1_47 : _GEN_10454; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11483 = 3'h4 == state ? ram_1_48 : _GEN_10455; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11484 = 3'h4 == state ? ram_1_49 : _GEN_10456; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11485 = 3'h4 == state ? ram_1_50 : _GEN_10457; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11486 = 3'h4 == state ? ram_1_51 : _GEN_10458; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11487 = 3'h4 == state ? ram_1_52 : _GEN_10459; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11488 = 3'h4 == state ? ram_1_53 : _GEN_10460; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11489 = 3'h4 == state ? ram_1_54 : _GEN_10461; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11490 = 3'h4 == state ? ram_1_55 : _GEN_10462; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11491 = 3'h4 == state ? ram_1_56 : _GEN_10463; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11492 = 3'h4 == state ? ram_1_57 : _GEN_10464; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11493 = 3'h4 == state ? ram_1_58 : _GEN_10465; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11494 = 3'h4 == state ? ram_1_59 : _GEN_10466; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11495 = 3'h4 == state ? ram_1_60 : _GEN_10467; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11496 = 3'h4 == state ? ram_1_61 : _GEN_10468; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11497 = 3'h4 == state ? ram_1_62 : _GEN_10469; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11498 = 3'h4 == state ? ram_1_63 : _GEN_10470; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11499 = 3'h4 == state ? ram_1_64 : _GEN_10471; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11500 = 3'h4 == state ? ram_1_65 : _GEN_10472; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11501 = 3'h4 == state ? ram_1_66 : _GEN_10473; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11502 = 3'h4 == state ? ram_1_67 : _GEN_10474; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11503 = 3'h4 == state ? ram_1_68 : _GEN_10475; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11504 = 3'h4 == state ? ram_1_69 : _GEN_10476; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11505 = 3'h4 == state ? ram_1_70 : _GEN_10477; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11506 = 3'h4 == state ? ram_1_71 : _GEN_10478; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11507 = 3'h4 == state ? ram_1_72 : _GEN_10479; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11508 = 3'h4 == state ? ram_1_73 : _GEN_10480; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11509 = 3'h4 == state ? ram_1_74 : _GEN_10481; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11510 = 3'h4 == state ? ram_1_75 : _GEN_10482; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11511 = 3'h4 == state ? ram_1_76 : _GEN_10483; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11512 = 3'h4 == state ? ram_1_77 : _GEN_10484; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11513 = 3'h4 == state ? ram_1_78 : _GEN_10485; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11514 = 3'h4 == state ? ram_1_79 : _GEN_10486; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11515 = 3'h4 == state ? ram_1_80 : _GEN_10487; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11516 = 3'h4 == state ? ram_1_81 : _GEN_10488; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11517 = 3'h4 == state ? ram_1_82 : _GEN_10489; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11518 = 3'h4 == state ? ram_1_83 : _GEN_10490; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11519 = 3'h4 == state ? ram_1_84 : _GEN_10491; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11520 = 3'h4 == state ? ram_1_85 : _GEN_10492; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11521 = 3'h4 == state ? ram_1_86 : _GEN_10493; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11522 = 3'h4 == state ? ram_1_87 : _GEN_10494; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11523 = 3'h4 == state ? ram_1_88 : _GEN_10495; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11524 = 3'h4 == state ? ram_1_89 : _GEN_10496; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11525 = 3'h4 == state ? ram_1_90 : _GEN_10497; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11526 = 3'h4 == state ? ram_1_91 : _GEN_10498; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11527 = 3'h4 == state ? ram_1_92 : _GEN_10499; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11528 = 3'h4 == state ? ram_1_93 : _GEN_10500; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11529 = 3'h4 == state ? ram_1_94 : _GEN_10501; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11530 = 3'h4 == state ? ram_1_95 : _GEN_10502; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11531 = 3'h4 == state ? ram_1_96 : _GEN_10503; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11532 = 3'h4 == state ? ram_1_97 : _GEN_10504; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11533 = 3'h4 == state ? ram_1_98 : _GEN_10505; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11534 = 3'h4 == state ? ram_1_99 : _GEN_10506; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11535 = 3'h4 == state ? ram_1_100 : _GEN_10507; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11536 = 3'h4 == state ? ram_1_101 : _GEN_10508; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11537 = 3'h4 == state ? ram_1_102 : _GEN_10509; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11538 = 3'h4 == state ? ram_1_103 : _GEN_10510; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11539 = 3'h4 == state ? ram_1_104 : _GEN_10511; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11540 = 3'h4 == state ? ram_1_105 : _GEN_10512; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11541 = 3'h4 == state ? ram_1_106 : _GEN_10513; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11542 = 3'h4 == state ? ram_1_107 : _GEN_10514; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11543 = 3'h4 == state ? ram_1_108 : _GEN_10515; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11544 = 3'h4 == state ? ram_1_109 : _GEN_10516; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11545 = 3'h4 == state ? ram_1_110 : _GEN_10517; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11546 = 3'h4 == state ? ram_1_111 : _GEN_10518; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11547 = 3'h4 == state ? ram_1_112 : _GEN_10519; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11548 = 3'h4 == state ? ram_1_113 : _GEN_10520; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11549 = 3'h4 == state ? ram_1_114 : _GEN_10521; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11550 = 3'h4 == state ? ram_1_115 : _GEN_10522; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11551 = 3'h4 == state ? ram_1_116 : _GEN_10523; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11552 = 3'h4 == state ? ram_1_117 : _GEN_10524; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11553 = 3'h4 == state ? ram_1_118 : _GEN_10525; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11554 = 3'h4 == state ? ram_1_119 : _GEN_10526; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11555 = 3'h4 == state ? ram_1_120 : _GEN_10527; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11556 = 3'h4 == state ? ram_1_121 : _GEN_10528; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11557 = 3'h4 == state ? ram_1_122 : _GEN_10529; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11558 = 3'h4 == state ? ram_1_123 : _GEN_10530; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11559 = 3'h4 == state ? ram_1_124 : _GEN_10531; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11560 = 3'h4 == state ? ram_1_125 : _GEN_10532; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11561 = 3'h4 == state ? ram_1_126 : _GEN_10533; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_11562 = 3'h4 == state ? ram_1_127 : _GEN_10534; // @[d_cache.scala 78:18 19:24]
  wire [31:0] _GEN_11563 = 3'h4 == state ? tag_1_0 : _GEN_10535; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11564 = 3'h4 == state ? tag_1_1 : _GEN_10536; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11565 = 3'h4 == state ? tag_1_2 : _GEN_10537; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11566 = 3'h4 == state ? tag_1_3 : _GEN_10538; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11567 = 3'h4 == state ? tag_1_4 : _GEN_10539; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11568 = 3'h4 == state ? tag_1_5 : _GEN_10540; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11569 = 3'h4 == state ? tag_1_6 : _GEN_10541; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11570 = 3'h4 == state ? tag_1_7 : _GEN_10542; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11571 = 3'h4 == state ? tag_1_8 : _GEN_10543; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11572 = 3'h4 == state ? tag_1_9 : _GEN_10544; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11573 = 3'h4 == state ? tag_1_10 : _GEN_10545; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11574 = 3'h4 == state ? tag_1_11 : _GEN_10546; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11575 = 3'h4 == state ? tag_1_12 : _GEN_10547; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11576 = 3'h4 == state ? tag_1_13 : _GEN_10548; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11577 = 3'h4 == state ? tag_1_14 : _GEN_10549; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11578 = 3'h4 == state ? tag_1_15 : _GEN_10550; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11579 = 3'h4 == state ? tag_1_16 : _GEN_10551; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11580 = 3'h4 == state ? tag_1_17 : _GEN_10552; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11581 = 3'h4 == state ? tag_1_18 : _GEN_10553; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11582 = 3'h4 == state ? tag_1_19 : _GEN_10554; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11583 = 3'h4 == state ? tag_1_20 : _GEN_10555; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11584 = 3'h4 == state ? tag_1_21 : _GEN_10556; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11585 = 3'h4 == state ? tag_1_22 : _GEN_10557; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11586 = 3'h4 == state ? tag_1_23 : _GEN_10558; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11587 = 3'h4 == state ? tag_1_24 : _GEN_10559; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11588 = 3'h4 == state ? tag_1_25 : _GEN_10560; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11589 = 3'h4 == state ? tag_1_26 : _GEN_10561; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11590 = 3'h4 == state ? tag_1_27 : _GEN_10562; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11591 = 3'h4 == state ? tag_1_28 : _GEN_10563; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11592 = 3'h4 == state ? tag_1_29 : _GEN_10564; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11593 = 3'h4 == state ? tag_1_30 : _GEN_10565; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11594 = 3'h4 == state ? tag_1_31 : _GEN_10566; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11595 = 3'h4 == state ? tag_1_32 : _GEN_10567; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11596 = 3'h4 == state ? tag_1_33 : _GEN_10568; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11597 = 3'h4 == state ? tag_1_34 : _GEN_10569; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11598 = 3'h4 == state ? tag_1_35 : _GEN_10570; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11599 = 3'h4 == state ? tag_1_36 : _GEN_10571; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11600 = 3'h4 == state ? tag_1_37 : _GEN_10572; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11601 = 3'h4 == state ? tag_1_38 : _GEN_10573; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11602 = 3'h4 == state ? tag_1_39 : _GEN_10574; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11603 = 3'h4 == state ? tag_1_40 : _GEN_10575; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11604 = 3'h4 == state ? tag_1_41 : _GEN_10576; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11605 = 3'h4 == state ? tag_1_42 : _GEN_10577; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11606 = 3'h4 == state ? tag_1_43 : _GEN_10578; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11607 = 3'h4 == state ? tag_1_44 : _GEN_10579; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11608 = 3'h4 == state ? tag_1_45 : _GEN_10580; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11609 = 3'h4 == state ? tag_1_46 : _GEN_10581; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11610 = 3'h4 == state ? tag_1_47 : _GEN_10582; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11611 = 3'h4 == state ? tag_1_48 : _GEN_10583; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11612 = 3'h4 == state ? tag_1_49 : _GEN_10584; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11613 = 3'h4 == state ? tag_1_50 : _GEN_10585; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11614 = 3'h4 == state ? tag_1_51 : _GEN_10586; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11615 = 3'h4 == state ? tag_1_52 : _GEN_10587; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11616 = 3'h4 == state ? tag_1_53 : _GEN_10588; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11617 = 3'h4 == state ? tag_1_54 : _GEN_10589; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11618 = 3'h4 == state ? tag_1_55 : _GEN_10590; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11619 = 3'h4 == state ? tag_1_56 : _GEN_10591; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11620 = 3'h4 == state ? tag_1_57 : _GEN_10592; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11621 = 3'h4 == state ? tag_1_58 : _GEN_10593; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11622 = 3'h4 == state ? tag_1_59 : _GEN_10594; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11623 = 3'h4 == state ? tag_1_60 : _GEN_10595; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11624 = 3'h4 == state ? tag_1_61 : _GEN_10596; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11625 = 3'h4 == state ? tag_1_62 : _GEN_10597; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11626 = 3'h4 == state ? tag_1_63 : _GEN_10598; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11627 = 3'h4 == state ? tag_1_64 : _GEN_10599; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11628 = 3'h4 == state ? tag_1_65 : _GEN_10600; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11629 = 3'h4 == state ? tag_1_66 : _GEN_10601; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11630 = 3'h4 == state ? tag_1_67 : _GEN_10602; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11631 = 3'h4 == state ? tag_1_68 : _GEN_10603; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11632 = 3'h4 == state ? tag_1_69 : _GEN_10604; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11633 = 3'h4 == state ? tag_1_70 : _GEN_10605; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11634 = 3'h4 == state ? tag_1_71 : _GEN_10606; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11635 = 3'h4 == state ? tag_1_72 : _GEN_10607; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11636 = 3'h4 == state ? tag_1_73 : _GEN_10608; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11637 = 3'h4 == state ? tag_1_74 : _GEN_10609; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11638 = 3'h4 == state ? tag_1_75 : _GEN_10610; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11639 = 3'h4 == state ? tag_1_76 : _GEN_10611; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11640 = 3'h4 == state ? tag_1_77 : _GEN_10612; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11641 = 3'h4 == state ? tag_1_78 : _GEN_10613; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11642 = 3'h4 == state ? tag_1_79 : _GEN_10614; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11643 = 3'h4 == state ? tag_1_80 : _GEN_10615; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11644 = 3'h4 == state ? tag_1_81 : _GEN_10616; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11645 = 3'h4 == state ? tag_1_82 : _GEN_10617; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11646 = 3'h4 == state ? tag_1_83 : _GEN_10618; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11647 = 3'h4 == state ? tag_1_84 : _GEN_10619; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11648 = 3'h4 == state ? tag_1_85 : _GEN_10620; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11649 = 3'h4 == state ? tag_1_86 : _GEN_10621; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11650 = 3'h4 == state ? tag_1_87 : _GEN_10622; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11651 = 3'h4 == state ? tag_1_88 : _GEN_10623; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11652 = 3'h4 == state ? tag_1_89 : _GEN_10624; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11653 = 3'h4 == state ? tag_1_90 : _GEN_10625; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11654 = 3'h4 == state ? tag_1_91 : _GEN_10626; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11655 = 3'h4 == state ? tag_1_92 : _GEN_10627; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11656 = 3'h4 == state ? tag_1_93 : _GEN_10628; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11657 = 3'h4 == state ? tag_1_94 : _GEN_10629; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11658 = 3'h4 == state ? tag_1_95 : _GEN_10630; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11659 = 3'h4 == state ? tag_1_96 : _GEN_10631; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11660 = 3'h4 == state ? tag_1_97 : _GEN_10632; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11661 = 3'h4 == state ? tag_1_98 : _GEN_10633; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11662 = 3'h4 == state ? tag_1_99 : _GEN_10634; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11663 = 3'h4 == state ? tag_1_100 : _GEN_10635; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11664 = 3'h4 == state ? tag_1_101 : _GEN_10636; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11665 = 3'h4 == state ? tag_1_102 : _GEN_10637; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11666 = 3'h4 == state ? tag_1_103 : _GEN_10638; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11667 = 3'h4 == state ? tag_1_104 : _GEN_10639; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11668 = 3'h4 == state ? tag_1_105 : _GEN_10640; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11669 = 3'h4 == state ? tag_1_106 : _GEN_10641; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11670 = 3'h4 == state ? tag_1_107 : _GEN_10642; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11671 = 3'h4 == state ? tag_1_108 : _GEN_10643; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11672 = 3'h4 == state ? tag_1_109 : _GEN_10644; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11673 = 3'h4 == state ? tag_1_110 : _GEN_10645; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11674 = 3'h4 == state ? tag_1_111 : _GEN_10646; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11675 = 3'h4 == state ? tag_1_112 : _GEN_10647; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11676 = 3'h4 == state ? tag_1_113 : _GEN_10648; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11677 = 3'h4 == state ? tag_1_114 : _GEN_10649; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11678 = 3'h4 == state ? tag_1_115 : _GEN_10650; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11679 = 3'h4 == state ? tag_1_116 : _GEN_10651; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11680 = 3'h4 == state ? tag_1_117 : _GEN_10652; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11681 = 3'h4 == state ? tag_1_118 : _GEN_10653; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11682 = 3'h4 == state ? tag_1_119 : _GEN_10654; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11683 = 3'h4 == state ? tag_1_120 : _GEN_10655; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11684 = 3'h4 == state ? tag_1_121 : _GEN_10656; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11685 = 3'h4 == state ? tag_1_122 : _GEN_10657; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11686 = 3'h4 == state ? tag_1_123 : _GEN_10658; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11687 = 3'h4 == state ? tag_1_124 : _GEN_10659; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11688 = 3'h4 == state ? tag_1_125 : _GEN_10660; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11689 = 3'h4 == state ? tag_1_126 : _GEN_10661; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_11690 = 3'h4 == state ? tag_1_127 : _GEN_10662; // @[d_cache.scala 78:18 21:24]
  wire  _GEN_11691 = 3'h4 == state ? valid_1_0 : _GEN_10663; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11692 = 3'h4 == state ? valid_1_1 : _GEN_10664; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11693 = 3'h4 == state ? valid_1_2 : _GEN_10665; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11694 = 3'h4 == state ? valid_1_3 : _GEN_10666; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11695 = 3'h4 == state ? valid_1_4 : _GEN_10667; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11696 = 3'h4 == state ? valid_1_5 : _GEN_10668; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11697 = 3'h4 == state ? valid_1_6 : _GEN_10669; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11698 = 3'h4 == state ? valid_1_7 : _GEN_10670; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11699 = 3'h4 == state ? valid_1_8 : _GEN_10671; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11700 = 3'h4 == state ? valid_1_9 : _GEN_10672; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11701 = 3'h4 == state ? valid_1_10 : _GEN_10673; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11702 = 3'h4 == state ? valid_1_11 : _GEN_10674; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11703 = 3'h4 == state ? valid_1_12 : _GEN_10675; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11704 = 3'h4 == state ? valid_1_13 : _GEN_10676; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11705 = 3'h4 == state ? valid_1_14 : _GEN_10677; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11706 = 3'h4 == state ? valid_1_15 : _GEN_10678; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11707 = 3'h4 == state ? valid_1_16 : _GEN_10679; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11708 = 3'h4 == state ? valid_1_17 : _GEN_10680; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11709 = 3'h4 == state ? valid_1_18 : _GEN_10681; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11710 = 3'h4 == state ? valid_1_19 : _GEN_10682; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11711 = 3'h4 == state ? valid_1_20 : _GEN_10683; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11712 = 3'h4 == state ? valid_1_21 : _GEN_10684; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11713 = 3'h4 == state ? valid_1_22 : _GEN_10685; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11714 = 3'h4 == state ? valid_1_23 : _GEN_10686; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11715 = 3'h4 == state ? valid_1_24 : _GEN_10687; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11716 = 3'h4 == state ? valid_1_25 : _GEN_10688; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11717 = 3'h4 == state ? valid_1_26 : _GEN_10689; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11718 = 3'h4 == state ? valid_1_27 : _GEN_10690; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11719 = 3'h4 == state ? valid_1_28 : _GEN_10691; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11720 = 3'h4 == state ? valid_1_29 : _GEN_10692; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11721 = 3'h4 == state ? valid_1_30 : _GEN_10693; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11722 = 3'h4 == state ? valid_1_31 : _GEN_10694; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11723 = 3'h4 == state ? valid_1_32 : _GEN_10695; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11724 = 3'h4 == state ? valid_1_33 : _GEN_10696; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11725 = 3'h4 == state ? valid_1_34 : _GEN_10697; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11726 = 3'h4 == state ? valid_1_35 : _GEN_10698; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11727 = 3'h4 == state ? valid_1_36 : _GEN_10699; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11728 = 3'h4 == state ? valid_1_37 : _GEN_10700; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11729 = 3'h4 == state ? valid_1_38 : _GEN_10701; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11730 = 3'h4 == state ? valid_1_39 : _GEN_10702; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11731 = 3'h4 == state ? valid_1_40 : _GEN_10703; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11732 = 3'h4 == state ? valid_1_41 : _GEN_10704; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11733 = 3'h4 == state ? valid_1_42 : _GEN_10705; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11734 = 3'h4 == state ? valid_1_43 : _GEN_10706; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11735 = 3'h4 == state ? valid_1_44 : _GEN_10707; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11736 = 3'h4 == state ? valid_1_45 : _GEN_10708; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11737 = 3'h4 == state ? valid_1_46 : _GEN_10709; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11738 = 3'h4 == state ? valid_1_47 : _GEN_10710; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11739 = 3'h4 == state ? valid_1_48 : _GEN_10711; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11740 = 3'h4 == state ? valid_1_49 : _GEN_10712; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11741 = 3'h4 == state ? valid_1_50 : _GEN_10713; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11742 = 3'h4 == state ? valid_1_51 : _GEN_10714; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11743 = 3'h4 == state ? valid_1_52 : _GEN_10715; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11744 = 3'h4 == state ? valid_1_53 : _GEN_10716; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11745 = 3'h4 == state ? valid_1_54 : _GEN_10717; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11746 = 3'h4 == state ? valid_1_55 : _GEN_10718; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11747 = 3'h4 == state ? valid_1_56 : _GEN_10719; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11748 = 3'h4 == state ? valid_1_57 : _GEN_10720; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11749 = 3'h4 == state ? valid_1_58 : _GEN_10721; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11750 = 3'h4 == state ? valid_1_59 : _GEN_10722; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11751 = 3'h4 == state ? valid_1_60 : _GEN_10723; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11752 = 3'h4 == state ? valid_1_61 : _GEN_10724; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11753 = 3'h4 == state ? valid_1_62 : _GEN_10725; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11754 = 3'h4 == state ? valid_1_63 : _GEN_10726; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11755 = 3'h4 == state ? valid_1_64 : _GEN_10727; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11756 = 3'h4 == state ? valid_1_65 : _GEN_10728; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11757 = 3'h4 == state ? valid_1_66 : _GEN_10729; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11758 = 3'h4 == state ? valid_1_67 : _GEN_10730; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11759 = 3'h4 == state ? valid_1_68 : _GEN_10731; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11760 = 3'h4 == state ? valid_1_69 : _GEN_10732; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11761 = 3'h4 == state ? valid_1_70 : _GEN_10733; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11762 = 3'h4 == state ? valid_1_71 : _GEN_10734; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11763 = 3'h4 == state ? valid_1_72 : _GEN_10735; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11764 = 3'h4 == state ? valid_1_73 : _GEN_10736; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11765 = 3'h4 == state ? valid_1_74 : _GEN_10737; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11766 = 3'h4 == state ? valid_1_75 : _GEN_10738; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11767 = 3'h4 == state ? valid_1_76 : _GEN_10739; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11768 = 3'h4 == state ? valid_1_77 : _GEN_10740; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11769 = 3'h4 == state ? valid_1_78 : _GEN_10741; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11770 = 3'h4 == state ? valid_1_79 : _GEN_10742; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11771 = 3'h4 == state ? valid_1_80 : _GEN_10743; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11772 = 3'h4 == state ? valid_1_81 : _GEN_10744; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11773 = 3'h4 == state ? valid_1_82 : _GEN_10745; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11774 = 3'h4 == state ? valid_1_83 : _GEN_10746; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11775 = 3'h4 == state ? valid_1_84 : _GEN_10747; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11776 = 3'h4 == state ? valid_1_85 : _GEN_10748; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11777 = 3'h4 == state ? valid_1_86 : _GEN_10749; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11778 = 3'h4 == state ? valid_1_87 : _GEN_10750; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11779 = 3'h4 == state ? valid_1_88 : _GEN_10751; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11780 = 3'h4 == state ? valid_1_89 : _GEN_10752; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11781 = 3'h4 == state ? valid_1_90 : _GEN_10753; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11782 = 3'h4 == state ? valid_1_91 : _GEN_10754; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11783 = 3'h4 == state ? valid_1_92 : _GEN_10755; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11784 = 3'h4 == state ? valid_1_93 : _GEN_10756; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11785 = 3'h4 == state ? valid_1_94 : _GEN_10757; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11786 = 3'h4 == state ? valid_1_95 : _GEN_10758; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11787 = 3'h4 == state ? valid_1_96 : _GEN_10759; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11788 = 3'h4 == state ? valid_1_97 : _GEN_10760; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11789 = 3'h4 == state ? valid_1_98 : _GEN_10761; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11790 = 3'h4 == state ? valid_1_99 : _GEN_10762; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11791 = 3'h4 == state ? valid_1_100 : _GEN_10763; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11792 = 3'h4 == state ? valid_1_101 : _GEN_10764; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11793 = 3'h4 == state ? valid_1_102 : _GEN_10765; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11794 = 3'h4 == state ? valid_1_103 : _GEN_10766; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11795 = 3'h4 == state ? valid_1_104 : _GEN_10767; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11796 = 3'h4 == state ? valid_1_105 : _GEN_10768; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11797 = 3'h4 == state ? valid_1_106 : _GEN_10769; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11798 = 3'h4 == state ? valid_1_107 : _GEN_10770; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11799 = 3'h4 == state ? valid_1_108 : _GEN_10771; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11800 = 3'h4 == state ? valid_1_109 : _GEN_10772; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11801 = 3'h4 == state ? valid_1_110 : _GEN_10773; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11802 = 3'h4 == state ? valid_1_111 : _GEN_10774; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11803 = 3'h4 == state ? valid_1_112 : _GEN_10775; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11804 = 3'h4 == state ? valid_1_113 : _GEN_10776; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11805 = 3'h4 == state ? valid_1_114 : _GEN_10777; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11806 = 3'h4 == state ? valid_1_115 : _GEN_10778; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11807 = 3'h4 == state ? valid_1_116 : _GEN_10779; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11808 = 3'h4 == state ? valid_1_117 : _GEN_10780; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11809 = 3'h4 == state ? valid_1_118 : _GEN_10781; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11810 = 3'h4 == state ? valid_1_119 : _GEN_10782; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11811 = 3'h4 == state ? valid_1_120 : _GEN_10783; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11812 = 3'h4 == state ? valid_1_121 : _GEN_10784; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11813 = 3'h4 == state ? valid_1_122 : _GEN_10785; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11814 = 3'h4 == state ? valid_1_123 : _GEN_10786; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11815 = 3'h4 == state ? valid_1_124 : _GEN_10787; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11816 = 3'h4 == state ? valid_1_125 : _GEN_10788; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11817 = 3'h4 == state ? valid_1_126 : _GEN_10789; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_11818 = 3'h4 == state ? valid_1_127 : _GEN_10790; // @[d_cache.scala 78:18 23:26]
  wire [63:0] _GEN_11819 = 3'h4 == state ? write_back_data : _GEN_10791; // @[d_cache.scala 78:18 29:34]
  wire [41:0] _GEN_11820 = 3'h4 == state ? {{10'd0}, write_back_addr} : _GEN_10792; // @[d_cache.scala 78:18 30:34]
  wire  _GEN_11821 = 3'h4 == state ? dirty_0_0 : _GEN_10793; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11822 = 3'h4 == state ? dirty_0_1 : _GEN_10794; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11823 = 3'h4 == state ? dirty_0_2 : _GEN_10795; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11824 = 3'h4 == state ? dirty_0_3 : _GEN_10796; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11825 = 3'h4 == state ? dirty_0_4 : _GEN_10797; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11826 = 3'h4 == state ? dirty_0_5 : _GEN_10798; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11827 = 3'h4 == state ? dirty_0_6 : _GEN_10799; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11828 = 3'h4 == state ? dirty_0_7 : _GEN_10800; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11829 = 3'h4 == state ? dirty_0_8 : _GEN_10801; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11830 = 3'h4 == state ? dirty_0_9 : _GEN_10802; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11831 = 3'h4 == state ? dirty_0_10 : _GEN_10803; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11832 = 3'h4 == state ? dirty_0_11 : _GEN_10804; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11833 = 3'h4 == state ? dirty_0_12 : _GEN_10805; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11834 = 3'h4 == state ? dirty_0_13 : _GEN_10806; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11835 = 3'h4 == state ? dirty_0_14 : _GEN_10807; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11836 = 3'h4 == state ? dirty_0_15 : _GEN_10808; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11837 = 3'h4 == state ? dirty_0_16 : _GEN_10809; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11838 = 3'h4 == state ? dirty_0_17 : _GEN_10810; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11839 = 3'h4 == state ? dirty_0_18 : _GEN_10811; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11840 = 3'h4 == state ? dirty_0_19 : _GEN_10812; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11841 = 3'h4 == state ? dirty_0_20 : _GEN_10813; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11842 = 3'h4 == state ? dirty_0_21 : _GEN_10814; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11843 = 3'h4 == state ? dirty_0_22 : _GEN_10815; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11844 = 3'h4 == state ? dirty_0_23 : _GEN_10816; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11845 = 3'h4 == state ? dirty_0_24 : _GEN_10817; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11846 = 3'h4 == state ? dirty_0_25 : _GEN_10818; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11847 = 3'h4 == state ? dirty_0_26 : _GEN_10819; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11848 = 3'h4 == state ? dirty_0_27 : _GEN_10820; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11849 = 3'h4 == state ? dirty_0_28 : _GEN_10821; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11850 = 3'h4 == state ? dirty_0_29 : _GEN_10822; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11851 = 3'h4 == state ? dirty_0_30 : _GEN_10823; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11852 = 3'h4 == state ? dirty_0_31 : _GEN_10824; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11853 = 3'h4 == state ? dirty_0_32 : _GEN_10825; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11854 = 3'h4 == state ? dirty_0_33 : _GEN_10826; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11855 = 3'h4 == state ? dirty_0_34 : _GEN_10827; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11856 = 3'h4 == state ? dirty_0_35 : _GEN_10828; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11857 = 3'h4 == state ? dirty_0_36 : _GEN_10829; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11858 = 3'h4 == state ? dirty_0_37 : _GEN_10830; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11859 = 3'h4 == state ? dirty_0_38 : _GEN_10831; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11860 = 3'h4 == state ? dirty_0_39 : _GEN_10832; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11861 = 3'h4 == state ? dirty_0_40 : _GEN_10833; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11862 = 3'h4 == state ? dirty_0_41 : _GEN_10834; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11863 = 3'h4 == state ? dirty_0_42 : _GEN_10835; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11864 = 3'h4 == state ? dirty_0_43 : _GEN_10836; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11865 = 3'h4 == state ? dirty_0_44 : _GEN_10837; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11866 = 3'h4 == state ? dirty_0_45 : _GEN_10838; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11867 = 3'h4 == state ? dirty_0_46 : _GEN_10839; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11868 = 3'h4 == state ? dirty_0_47 : _GEN_10840; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11869 = 3'h4 == state ? dirty_0_48 : _GEN_10841; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11870 = 3'h4 == state ? dirty_0_49 : _GEN_10842; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11871 = 3'h4 == state ? dirty_0_50 : _GEN_10843; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11872 = 3'h4 == state ? dirty_0_51 : _GEN_10844; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11873 = 3'h4 == state ? dirty_0_52 : _GEN_10845; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11874 = 3'h4 == state ? dirty_0_53 : _GEN_10846; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11875 = 3'h4 == state ? dirty_0_54 : _GEN_10847; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11876 = 3'h4 == state ? dirty_0_55 : _GEN_10848; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11877 = 3'h4 == state ? dirty_0_56 : _GEN_10849; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11878 = 3'h4 == state ? dirty_0_57 : _GEN_10850; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11879 = 3'h4 == state ? dirty_0_58 : _GEN_10851; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11880 = 3'h4 == state ? dirty_0_59 : _GEN_10852; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11881 = 3'h4 == state ? dirty_0_60 : _GEN_10853; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11882 = 3'h4 == state ? dirty_0_61 : _GEN_10854; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11883 = 3'h4 == state ? dirty_0_62 : _GEN_10855; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11884 = 3'h4 == state ? dirty_0_63 : _GEN_10856; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11885 = 3'h4 == state ? dirty_0_64 : _GEN_10857; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11886 = 3'h4 == state ? dirty_0_65 : _GEN_10858; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11887 = 3'h4 == state ? dirty_0_66 : _GEN_10859; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11888 = 3'h4 == state ? dirty_0_67 : _GEN_10860; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11889 = 3'h4 == state ? dirty_0_68 : _GEN_10861; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11890 = 3'h4 == state ? dirty_0_69 : _GEN_10862; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11891 = 3'h4 == state ? dirty_0_70 : _GEN_10863; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11892 = 3'h4 == state ? dirty_0_71 : _GEN_10864; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11893 = 3'h4 == state ? dirty_0_72 : _GEN_10865; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11894 = 3'h4 == state ? dirty_0_73 : _GEN_10866; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11895 = 3'h4 == state ? dirty_0_74 : _GEN_10867; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11896 = 3'h4 == state ? dirty_0_75 : _GEN_10868; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11897 = 3'h4 == state ? dirty_0_76 : _GEN_10869; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11898 = 3'h4 == state ? dirty_0_77 : _GEN_10870; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11899 = 3'h4 == state ? dirty_0_78 : _GEN_10871; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11900 = 3'h4 == state ? dirty_0_79 : _GEN_10872; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11901 = 3'h4 == state ? dirty_0_80 : _GEN_10873; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11902 = 3'h4 == state ? dirty_0_81 : _GEN_10874; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11903 = 3'h4 == state ? dirty_0_82 : _GEN_10875; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11904 = 3'h4 == state ? dirty_0_83 : _GEN_10876; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11905 = 3'h4 == state ? dirty_0_84 : _GEN_10877; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11906 = 3'h4 == state ? dirty_0_85 : _GEN_10878; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11907 = 3'h4 == state ? dirty_0_86 : _GEN_10879; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11908 = 3'h4 == state ? dirty_0_87 : _GEN_10880; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11909 = 3'h4 == state ? dirty_0_88 : _GEN_10881; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11910 = 3'h4 == state ? dirty_0_89 : _GEN_10882; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11911 = 3'h4 == state ? dirty_0_90 : _GEN_10883; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11912 = 3'h4 == state ? dirty_0_91 : _GEN_10884; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11913 = 3'h4 == state ? dirty_0_92 : _GEN_10885; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11914 = 3'h4 == state ? dirty_0_93 : _GEN_10886; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11915 = 3'h4 == state ? dirty_0_94 : _GEN_10887; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11916 = 3'h4 == state ? dirty_0_95 : _GEN_10888; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11917 = 3'h4 == state ? dirty_0_96 : _GEN_10889; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11918 = 3'h4 == state ? dirty_0_97 : _GEN_10890; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11919 = 3'h4 == state ? dirty_0_98 : _GEN_10891; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11920 = 3'h4 == state ? dirty_0_99 : _GEN_10892; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11921 = 3'h4 == state ? dirty_0_100 : _GEN_10893; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11922 = 3'h4 == state ? dirty_0_101 : _GEN_10894; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11923 = 3'h4 == state ? dirty_0_102 : _GEN_10895; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11924 = 3'h4 == state ? dirty_0_103 : _GEN_10896; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11925 = 3'h4 == state ? dirty_0_104 : _GEN_10897; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11926 = 3'h4 == state ? dirty_0_105 : _GEN_10898; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11927 = 3'h4 == state ? dirty_0_106 : _GEN_10899; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11928 = 3'h4 == state ? dirty_0_107 : _GEN_10900; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11929 = 3'h4 == state ? dirty_0_108 : _GEN_10901; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11930 = 3'h4 == state ? dirty_0_109 : _GEN_10902; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11931 = 3'h4 == state ? dirty_0_110 : _GEN_10903; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11932 = 3'h4 == state ? dirty_0_111 : _GEN_10904; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11933 = 3'h4 == state ? dirty_0_112 : _GEN_10905; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11934 = 3'h4 == state ? dirty_0_113 : _GEN_10906; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11935 = 3'h4 == state ? dirty_0_114 : _GEN_10907; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11936 = 3'h4 == state ? dirty_0_115 : _GEN_10908; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11937 = 3'h4 == state ? dirty_0_116 : _GEN_10909; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11938 = 3'h4 == state ? dirty_0_117 : _GEN_10910; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11939 = 3'h4 == state ? dirty_0_118 : _GEN_10911; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11940 = 3'h4 == state ? dirty_0_119 : _GEN_10912; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11941 = 3'h4 == state ? dirty_0_120 : _GEN_10913; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11942 = 3'h4 == state ? dirty_0_121 : _GEN_10914; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11943 = 3'h4 == state ? dirty_0_122 : _GEN_10915; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11944 = 3'h4 == state ? dirty_0_123 : _GEN_10916; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11945 = 3'h4 == state ? dirty_0_124 : _GEN_10917; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11946 = 3'h4 == state ? dirty_0_125 : _GEN_10918; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11947 = 3'h4 == state ? dirty_0_126 : _GEN_10919; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11948 = 3'h4 == state ? dirty_0_127 : _GEN_10920; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_11949 = 3'h4 == state ? dirty_1_0 : _GEN_10921; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11950 = 3'h4 == state ? dirty_1_1 : _GEN_10922; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11951 = 3'h4 == state ? dirty_1_2 : _GEN_10923; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11952 = 3'h4 == state ? dirty_1_3 : _GEN_10924; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11953 = 3'h4 == state ? dirty_1_4 : _GEN_10925; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11954 = 3'h4 == state ? dirty_1_5 : _GEN_10926; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11955 = 3'h4 == state ? dirty_1_6 : _GEN_10927; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11956 = 3'h4 == state ? dirty_1_7 : _GEN_10928; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11957 = 3'h4 == state ? dirty_1_8 : _GEN_10929; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11958 = 3'h4 == state ? dirty_1_9 : _GEN_10930; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11959 = 3'h4 == state ? dirty_1_10 : _GEN_10931; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11960 = 3'h4 == state ? dirty_1_11 : _GEN_10932; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11961 = 3'h4 == state ? dirty_1_12 : _GEN_10933; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11962 = 3'h4 == state ? dirty_1_13 : _GEN_10934; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11963 = 3'h4 == state ? dirty_1_14 : _GEN_10935; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11964 = 3'h4 == state ? dirty_1_15 : _GEN_10936; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11965 = 3'h4 == state ? dirty_1_16 : _GEN_10937; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11966 = 3'h4 == state ? dirty_1_17 : _GEN_10938; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11967 = 3'h4 == state ? dirty_1_18 : _GEN_10939; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11968 = 3'h4 == state ? dirty_1_19 : _GEN_10940; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11969 = 3'h4 == state ? dirty_1_20 : _GEN_10941; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11970 = 3'h4 == state ? dirty_1_21 : _GEN_10942; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11971 = 3'h4 == state ? dirty_1_22 : _GEN_10943; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11972 = 3'h4 == state ? dirty_1_23 : _GEN_10944; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11973 = 3'h4 == state ? dirty_1_24 : _GEN_10945; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11974 = 3'h4 == state ? dirty_1_25 : _GEN_10946; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11975 = 3'h4 == state ? dirty_1_26 : _GEN_10947; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11976 = 3'h4 == state ? dirty_1_27 : _GEN_10948; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11977 = 3'h4 == state ? dirty_1_28 : _GEN_10949; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11978 = 3'h4 == state ? dirty_1_29 : _GEN_10950; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11979 = 3'h4 == state ? dirty_1_30 : _GEN_10951; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11980 = 3'h4 == state ? dirty_1_31 : _GEN_10952; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11981 = 3'h4 == state ? dirty_1_32 : _GEN_10953; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11982 = 3'h4 == state ? dirty_1_33 : _GEN_10954; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11983 = 3'h4 == state ? dirty_1_34 : _GEN_10955; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11984 = 3'h4 == state ? dirty_1_35 : _GEN_10956; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11985 = 3'h4 == state ? dirty_1_36 : _GEN_10957; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11986 = 3'h4 == state ? dirty_1_37 : _GEN_10958; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11987 = 3'h4 == state ? dirty_1_38 : _GEN_10959; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11988 = 3'h4 == state ? dirty_1_39 : _GEN_10960; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11989 = 3'h4 == state ? dirty_1_40 : _GEN_10961; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11990 = 3'h4 == state ? dirty_1_41 : _GEN_10962; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11991 = 3'h4 == state ? dirty_1_42 : _GEN_10963; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11992 = 3'h4 == state ? dirty_1_43 : _GEN_10964; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11993 = 3'h4 == state ? dirty_1_44 : _GEN_10965; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11994 = 3'h4 == state ? dirty_1_45 : _GEN_10966; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11995 = 3'h4 == state ? dirty_1_46 : _GEN_10967; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11996 = 3'h4 == state ? dirty_1_47 : _GEN_10968; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11997 = 3'h4 == state ? dirty_1_48 : _GEN_10969; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11998 = 3'h4 == state ? dirty_1_49 : _GEN_10970; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_11999 = 3'h4 == state ? dirty_1_50 : _GEN_10971; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12000 = 3'h4 == state ? dirty_1_51 : _GEN_10972; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12001 = 3'h4 == state ? dirty_1_52 : _GEN_10973; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12002 = 3'h4 == state ? dirty_1_53 : _GEN_10974; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12003 = 3'h4 == state ? dirty_1_54 : _GEN_10975; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12004 = 3'h4 == state ? dirty_1_55 : _GEN_10976; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12005 = 3'h4 == state ? dirty_1_56 : _GEN_10977; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12006 = 3'h4 == state ? dirty_1_57 : _GEN_10978; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12007 = 3'h4 == state ? dirty_1_58 : _GEN_10979; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12008 = 3'h4 == state ? dirty_1_59 : _GEN_10980; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12009 = 3'h4 == state ? dirty_1_60 : _GEN_10981; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12010 = 3'h4 == state ? dirty_1_61 : _GEN_10982; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12011 = 3'h4 == state ? dirty_1_62 : _GEN_10983; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12012 = 3'h4 == state ? dirty_1_63 : _GEN_10984; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12013 = 3'h4 == state ? dirty_1_64 : _GEN_10985; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12014 = 3'h4 == state ? dirty_1_65 : _GEN_10986; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12015 = 3'h4 == state ? dirty_1_66 : _GEN_10987; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12016 = 3'h4 == state ? dirty_1_67 : _GEN_10988; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12017 = 3'h4 == state ? dirty_1_68 : _GEN_10989; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12018 = 3'h4 == state ? dirty_1_69 : _GEN_10990; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12019 = 3'h4 == state ? dirty_1_70 : _GEN_10991; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12020 = 3'h4 == state ? dirty_1_71 : _GEN_10992; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12021 = 3'h4 == state ? dirty_1_72 : _GEN_10993; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12022 = 3'h4 == state ? dirty_1_73 : _GEN_10994; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12023 = 3'h4 == state ? dirty_1_74 : _GEN_10995; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12024 = 3'h4 == state ? dirty_1_75 : _GEN_10996; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12025 = 3'h4 == state ? dirty_1_76 : _GEN_10997; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12026 = 3'h4 == state ? dirty_1_77 : _GEN_10998; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12027 = 3'h4 == state ? dirty_1_78 : _GEN_10999; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12028 = 3'h4 == state ? dirty_1_79 : _GEN_11000; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12029 = 3'h4 == state ? dirty_1_80 : _GEN_11001; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12030 = 3'h4 == state ? dirty_1_81 : _GEN_11002; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12031 = 3'h4 == state ? dirty_1_82 : _GEN_11003; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12032 = 3'h4 == state ? dirty_1_83 : _GEN_11004; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12033 = 3'h4 == state ? dirty_1_84 : _GEN_11005; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12034 = 3'h4 == state ? dirty_1_85 : _GEN_11006; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12035 = 3'h4 == state ? dirty_1_86 : _GEN_11007; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12036 = 3'h4 == state ? dirty_1_87 : _GEN_11008; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12037 = 3'h4 == state ? dirty_1_88 : _GEN_11009; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12038 = 3'h4 == state ? dirty_1_89 : _GEN_11010; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12039 = 3'h4 == state ? dirty_1_90 : _GEN_11011; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12040 = 3'h4 == state ? dirty_1_91 : _GEN_11012; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12041 = 3'h4 == state ? dirty_1_92 : _GEN_11013; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12042 = 3'h4 == state ? dirty_1_93 : _GEN_11014; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12043 = 3'h4 == state ? dirty_1_94 : _GEN_11015; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12044 = 3'h4 == state ? dirty_1_95 : _GEN_11016; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12045 = 3'h4 == state ? dirty_1_96 : _GEN_11017; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12046 = 3'h4 == state ? dirty_1_97 : _GEN_11018; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12047 = 3'h4 == state ? dirty_1_98 : _GEN_11019; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12048 = 3'h4 == state ? dirty_1_99 : _GEN_11020; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12049 = 3'h4 == state ? dirty_1_100 : _GEN_11021; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12050 = 3'h4 == state ? dirty_1_101 : _GEN_11022; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12051 = 3'h4 == state ? dirty_1_102 : _GEN_11023; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12052 = 3'h4 == state ? dirty_1_103 : _GEN_11024; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12053 = 3'h4 == state ? dirty_1_104 : _GEN_11025; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12054 = 3'h4 == state ? dirty_1_105 : _GEN_11026; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12055 = 3'h4 == state ? dirty_1_106 : _GEN_11027; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12056 = 3'h4 == state ? dirty_1_107 : _GEN_11028; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12057 = 3'h4 == state ? dirty_1_108 : _GEN_11029; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12058 = 3'h4 == state ? dirty_1_109 : _GEN_11030; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12059 = 3'h4 == state ? dirty_1_110 : _GEN_11031; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12060 = 3'h4 == state ? dirty_1_111 : _GEN_11032; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12061 = 3'h4 == state ? dirty_1_112 : _GEN_11033; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12062 = 3'h4 == state ? dirty_1_113 : _GEN_11034; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12063 = 3'h4 == state ? dirty_1_114 : _GEN_11035; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12064 = 3'h4 == state ? dirty_1_115 : _GEN_11036; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12065 = 3'h4 == state ? dirty_1_116 : _GEN_11037; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12066 = 3'h4 == state ? dirty_1_117 : _GEN_11038; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12067 = 3'h4 == state ? dirty_1_118 : _GEN_11039; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12068 = 3'h4 == state ? dirty_1_119 : _GEN_11040; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12069 = 3'h4 == state ? dirty_1_120 : _GEN_11041; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12070 = 3'h4 == state ? dirty_1_121 : _GEN_11042; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12071 = 3'h4 == state ? dirty_1_122 : _GEN_11043; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12072 = 3'h4 == state ? dirty_1_123 : _GEN_11044; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12073 = 3'h4 == state ? dirty_1_124 : _GEN_11045; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12074 = 3'h4 == state ? dirty_1_125 : _GEN_11046; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12075 = 3'h4 == state ? dirty_1_126 : _GEN_11047; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12076 = 3'h4 == state ? dirty_1_127 : _GEN_11048; // @[d_cache.scala 78:18 25:26]
  wire [2:0] _GEN_12077 = 3'h3 == state ? _GEN_2571 : _GEN_11049; // @[d_cache.scala 78:18]
  wire [63:0] _GEN_12078 = 3'h3 == state ? _GEN_2572 : receive_data; // @[d_cache.scala 78:18 34:31]
  wire [63:0] _GEN_12079 = 3'h3 == state ? ram_0_0 : _GEN_11050; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12080 = 3'h3 == state ? ram_0_1 : _GEN_11051; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12081 = 3'h3 == state ? ram_0_2 : _GEN_11052; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12082 = 3'h3 == state ? ram_0_3 : _GEN_11053; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12083 = 3'h3 == state ? ram_0_4 : _GEN_11054; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12084 = 3'h3 == state ? ram_0_5 : _GEN_11055; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12085 = 3'h3 == state ? ram_0_6 : _GEN_11056; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12086 = 3'h3 == state ? ram_0_7 : _GEN_11057; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12087 = 3'h3 == state ? ram_0_8 : _GEN_11058; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12088 = 3'h3 == state ? ram_0_9 : _GEN_11059; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12089 = 3'h3 == state ? ram_0_10 : _GEN_11060; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12090 = 3'h3 == state ? ram_0_11 : _GEN_11061; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12091 = 3'h3 == state ? ram_0_12 : _GEN_11062; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12092 = 3'h3 == state ? ram_0_13 : _GEN_11063; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12093 = 3'h3 == state ? ram_0_14 : _GEN_11064; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12094 = 3'h3 == state ? ram_0_15 : _GEN_11065; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12095 = 3'h3 == state ? ram_0_16 : _GEN_11066; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12096 = 3'h3 == state ? ram_0_17 : _GEN_11067; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12097 = 3'h3 == state ? ram_0_18 : _GEN_11068; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12098 = 3'h3 == state ? ram_0_19 : _GEN_11069; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12099 = 3'h3 == state ? ram_0_20 : _GEN_11070; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12100 = 3'h3 == state ? ram_0_21 : _GEN_11071; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12101 = 3'h3 == state ? ram_0_22 : _GEN_11072; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12102 = 3'h3 == state ? ram_0_23 : _GEN_11073; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12103 = 3'h3 == state ? ram_0_24 : _GEN_11074; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12104 = 3'h3 == state ? ram_0_25 : _GEN_11075; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12105 = 3'h3 == state ? ram_0_26 : _GEN_11076; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12106 = 3'h3 == state ? ram_0_27 : _GEN_11077; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12107 = 3'h3 == state ? ram_0_28 : _GEN_11078; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12108 = 3'h3 == state ? ram_0_29 : _GEN_11079; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12109 = 3'h3 == state ? ram_0_30 : _GEN_11080; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12110 = 3'h3 == state ? ram_0_31 : _GEN_11081; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12111 = 3'h3 == state ? ram_0_32 : _GEN_11082; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12112 = 3'h3 == state ? ram_0_33 : _GEN_11083; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12113 = 3'h3 == state ? ram_0_34 : _GEN_11084; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12114 = 3'h3 == state ? ram_0_35 : _GEN_11085; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12115 = 3'h3 == state ? ram_0_36 : _GEN_11086; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12116 = 3'h3 == state ? ram_0_37 : _GEN_11087; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12117 = 3'h3 == state ? ram_0_38 : _GEN_11088; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12118 = 3'h3 == state ? ram_0_39 : _GEN_11089; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12119 = 3'h3 == state ? ram_0_40 : _GEN_11090; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12120 = 3'h3 == state ? ram_0_41 : _GEN_11091; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12121 = 3'h3 == state ? ram_0_42 : _GEN_11092; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12122 = 3'h3 == state ? ram_0_43 : _GEN_11093; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12123 = 3'h3 == state ? ram_0_44 : _GEN_11094; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12124 = 3'h3 == state ? ram_0_45 : _GEN_11095; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12125 = 3'h3 == state ? ram_0_46 : _GEN_11096; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12126 = 3'h3 == state ? ram_0_47 : _GEN_11097; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12127 = 3'h3 == state ? ram_0_48 : _GEN_11098; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12128 = 3'h3 == state ? ram_0_49 : _GEN_11099; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12129 = 3'h3 == state ? ram_0_50 : _GEN_11100; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12130 = 3'h3 == state ? ram_0_51 : _GEN_11101; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12131 = 3'h3 == state ? ram_0_52 : _GEN_11102; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12132 = 3'h3 == state ? ram_0_53 : _GEN_11103; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12133 = 3'h3 == state ? ram_0_54 : _GEN_11104; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12134 = 3'h3 == state ? ram_0_55 : _GEN_11105; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12135 = 3'h3 == state ? ram_0_56 : _GEN_11106; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12136 = 3'h3 == state ? ram_0_57 : _GEN_11107; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12137 = 3'h3 == state ? ram_0_58 : _GEN_11108; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12138 = 3'h3 == state ? ram_0_59 : _GEN_11109; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12139 = 3'h3 == state ? ram_0_60 : _GEN_11110; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12140 = 3'h3 == state ? ram_0_61 : _GEN_11111; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12141 = 3'h3 == state ? ram_0_62 : _GEN_11112; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12142 = 3'h3 == state ? ram_0_63 : _GEN_11113; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12143 = 3'h3 == state ? ram_0_64 : _GEN_11114; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12144 = 3'h3 == state ? ram_0_65 : _GEN_11115; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12145 = 3'h3 == state ? ram_0_66 : _GEN_11116; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12146 = 3'h3 == state ? ram_0_67 : _GEN_11117; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12147 = 3'h3 == state ? ram_0_68 : _GEN_11118; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12148 = 3'h3 == state ? ram_0_69 : _GEN_11119; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12149 = 3'h3 == state ? ram_0_70 : _GEN_11120; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12150 = 3'h3 == state ? ram_0_71 : _GEN_11121; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12151 = 3'h3 == state ? ram_0_72 : _GEN_11122; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12152 = 3'h3 == state ? ram_0_73 : _GEN_11123; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12153 = 3'h3 == state ? ram_0_74 : _GEN_11124; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12154 = 3'h3 == state ? ram_0_75 : _GEN_11125; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12155 = 3'h3 == state ? ram_0_76 : _GEN_11126; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12156 = 3'h3 == state ? ram_0_77 : _GEN_11127; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12157 = 3'h3 == state ? ram_0_78 : _GEN_11128; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12158 = 3'h3 == state ? ram_0_79 : _GEN_11129; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12159 = 3'h3 == state ? ram_0_80 : _GEN_11130; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12160 = 3'h3 == state ? ram_0_81 : _GEN_11131; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12161 = 3'h3 == state ? ram_0_82 : _GEN_11132; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12162 = 3'h3 == state ? ram_0_83 : _GEN_11133; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12163 = 3'h3 == state ? ram_0_84 : _GEN_11134; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12164 = 3'h3 == state ? ram_0_85 : _GEN_11135; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12165 = 3'h3 == state ? ram_0_86 : _GEN_11136; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12166 = 3'h3 == state ? ram_0_87 : _GEN_11137; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12167 = 3'h3 == state ? ram_0_88 : _GEN_11138; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12168 = 3'h3 == state ? ram_0_89 : _GEN_11139; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12169 = 3'h3 == state ? ram_0_90 : _GEN_11140; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12170 = 3'h3 == state ? ram_0_91 : _GEN_11141; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12171 = 3'h3 == state ? ram_0_92 : _GEN_11142; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12172 = 3'h3 == state ? ram_0_93 : _GEN_11143; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12173 = 3'h3 == state ? ram_0_94 : _GEN_11144; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12174 = 3'h3 == state ? ram_0_95 : _GEN_11145; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12175 = 3'h3 == state ? ram_0_96 : _GEN_11146; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12176 = 3'h3 == state ? ram_0_97 : _GEN_11147; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12177 = 3'h3 == state ? ram_0_98 : _GEN_11148; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12178 = 3'h3 == state ? ram_0_99 : _GEN_11149; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12179 = 3'h3 == state ? ram_0_100 : _GEN_11150; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12180 = 3'h3 == state ? ram_0_101 : _GEN_11151; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12181 = 3'h3 == state ? ram_0_102 : _GEN_11152; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12182 = 3'h3 == state ? ram_0_103 : _GEN_11153; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12183 = 3'h3 == state ? ram_0_104 : _GEN_11154; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12184 = 3'h3 == state ? ram_0_105 : _GEN_11155; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12185 = 3'h3 == state ? ram_0_106 : _GEN_11156; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12186 = 3'h3 == state ? ram_0_107 : _GEN_11157; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12187 = 3'h3 == state ? ram_0_108 : _GEN_11158; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12188 = 3'h3 == state ? ram_0_109 : _GEN_11159; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12189 = 3'h3 == state ? ram_0_110 : _GEN_11160; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12190 = 3'h3 == state ? ram_0_111 : _GEN_11161; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12191 = 3'h3 == state ? ram_0_112 : _GEN_11162; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12192 = 3'h3 == state ? ram_0_113 : _GEN_11163; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12193 = 3'h3 == state ? ram_0_114 : _GEN_11164; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12194 = 3'h3 == state ? ram_0_115 : _GEN_11165; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12195 = 3'h3 == state ? ram_0_116 : _GEN_11166; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12196 = 3'h3 == state ? ram_0_117 : _GEN_11167; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12197 = 3'h3 == state ? ram_0_118 : _GEN_11168; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12198 = 3'h3 == state ? ram_0_119 : _GEN_11169; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12199 = 3'h3 == state ? ram_0_120 : _GEN_11170; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12200 = 3'h3 == state ? ram_0_121 : _GEN_11171; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12201 = 3'h3 == state ? ram_0_122 : _GEN_11172; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12202 = 3'h3 == state ? ram_0_123 : _GEN_11173; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12203 = 3'h3 == state ? ram_0_124 : _GEN_11174; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12204 = 3'h3 == state ? ram_0_125 : _GEN_11175; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12205 = 3'h3 == state ? ram_0_126 : _GEN_11176; // @[d_cache.scala 78:18 18:24]
  wire [63:0] _GEN_12206 = 3'h3 == state ? ram_0_127 : _GEN_11177; // @[d_cache.scala 78:18 18:24]
  wire [31:0] _GEN_12207 = 3'h3 == state ? tag_0_0 : _GEN_11178; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12208 = 3'h3 == state ? tag_0_1 : _GEN_11179; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12209 = 3'h3 == state ? tag_0_2 : _GEN_11180; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12210 = 3'h3 == state ? tag_0_3 : _GEN_11181; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12211 = 3'h3 == state ? tag_0_4 : _GEN_11182; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12212 = 3'h3 == state ? tag_0_5 : _GEN_11183; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12213 = 3'h3 == state ? tag_0_6 : _GEN_11184; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12214 = 3'h3 == state ? tag_0_7 : _GEN_11185; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12215 = 3'h3 == state ? tag_0_8 : _GEN_11186; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12216 = 3'h3 == state ? tag_0_9 : _GEN_11187; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12217 = 3'h3 == state ? tag_0_10 : _GEN_11188; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12218 = 3'h3 == state ? tag_0_11 : _GEN_11189; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12219 = 3'h3 == state ? tag_0_12 : _GEN_11190; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12220 = 3'h3 == state ? tag_0_13 : _GEN_11191; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12221 = 3'h3 == state ? tag_0_14 : _GEN_11192; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12222 = 3'h3 == state ? tag_0_15 : _GEN_11193; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12223 = 3'h3 == state ? tag_0_16 : _GEN_11194; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12224 = 3'h3 == state ? tag_0_17 : _GEN_11195; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12225 = 3'h3 == state ? tag_0_18 : _GEN_11196; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12226 = 3'h3 == state ? tag_0_19 : _GEN_11197; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12227 = 3'h3 == state ? tag_0_20 : _GEN_11198; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12228 = 3'h3 == state ? tag_0_21 : _GEN_11199; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12229 = 3'h3 == state ? tag_0_22 : _GEN_11200; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12230 = 3'h3 == state ? tag_0_23 : _GEN_11201; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12231 = 3'h3 == state ? tag_0_24 : _GEN_11202; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12232 = 3'h3 == state ? tag_0_25 : _GEN_11203; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12233 = 3'h3 == state ? tag_0_26 : _GEN_11204; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12234 = 3'h3 == state ? tag_0_27 : _GEN_11205; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12235 = 3'h3 == state ? tag_0_28 : _GEN_11206; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12236 = 3'h3 == state ? tag_0_29 : _GEN_11207; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12237 = 3'h3 == state ? tag_0_30 : _GEN_11208; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12238 = 3'h3 == state ? tag_0_31 : _GEN_11209; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12239 = 3'h3 == state ? tag_0_32 : _GEN_11210; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12240 = 3'h3 == state ? tag_0_33 : _GEN_11211; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12241 = 3'h3 == state ? tag_0_34 : _GEN_11212; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12242 = 3'h3 == state ? tag_0_35 : _GEN_11213; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12243 = 3'h3 == state ? tag_0_36 : _GEN_11214; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12244 = 3'h3 == state ? tag_0_37 : _GEN_11215; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12245 = 3'h3 == state ? tag_0_38 : _GEN_11216; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12246 = 3'h3 == state ? tag_0_39 : _GEN_11217; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12247 = 3'h3 == state ? tag_0_40 : _GEN_11218; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12248 = 3'h3 == state ? tag_0_41 : _GEN_11219; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12249 = 3'h3 == state ? tag_0_42 : _GEN_11220; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12250 = 3'h3 == state ? tag_0_43 : _GEN_11221; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12251 = 3'h3 == state ? tag_0_44 : _GEN_11222; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12252 = 3'h3 == state ? tag_0_45 : _GEN_11223; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12253 = 3'h3 == state ? tag_0_46 : _GEN_11224; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12254 = 3'h3 == state ? tag_0_47 : _GEN_11225; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12255 = 3'h3 == state ? tag_0_48 : _GEN_11226; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12256 = 3'h3 == state ? tag_0_49 : _GEN_11227; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12257 = 3'h3 == state ? tag_0_50 : _GEN_11228; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12258 = 3'h3 == state ? tag_0_51 : _GEN_11229; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12259 = 3'h3 == state ? tag_0_52 : _GEN_11230; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12260 = 3'h3 == state ? tag_0_53 : _GEN_11231; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12261 = 3'h3 == state ? tag_0_54 : _GEN_11232; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12262 = 3'h3 == state ? tag_0_55 : _GEN_11233; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12263 = 3'h3 == state ? tag_0_56 : _GEN_11234; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12264 = 3'h3 == state ? tag_0_57 : _GEN_11235; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12265 = 3'h3 == state ? tag_0_58 : _GEN_11236; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12266 = 3'h3 == state ? tag_0_59 : _GEN_11237; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12267 = 3'h3 == state ? tag_0_60 : _GEN_11238; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12268 = 3'h3 == state ? tag_0_61 : _GEN_11239; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12269 = 3'h3 == state ? tag_0_62 : _GEN_11240; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12270 = 3'h3 == state ? tag_0_63 : _GEN_11241; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12271 = 3'h3 == state ? tag_0_64 : _GEN_11242; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12272 = 3'h3 == state ? tag_0_65 : _GEN_11243; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12273 = 3'h3 == state ? tag_0_66 : _GEN_11244; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12274 = 3'h3 == state ? tag_0_67 : _GEN_11245; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12275 = 3'h3 == state ? tag_0_68 : _GEN_11246; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12276 = 3'h3 == state ? tag_0_69 : _GEN_11247; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12277 = 3'h3 == state ? tag_0_70 : _GEN_11248; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12278 = 3'h3 == state ? tag_0_71 : _GEN_11249; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12279 = 3'h3 == state ? tag_0_72 : _GEN_11250; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12280 = 3'h3 == state ? tag_0_73 : _GEN_11251; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12281 = 3'h3 == state ? tag_0_74 : _GEN_11252; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12282 = 3'h3 == state ? tag_0_75 : _GEN_11253; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12283 = 3'h3 == state ? tag_0_76 : _GEN_11254; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12284 = 3'h3 == state ? tag_0_77 : _GEN_11255; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12285 = 3'h3 == state ? tag_0_78 : _GEN_11256; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12286 = 3'h3 == state ? tag_0_79 : _GEN_11257; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12287 = 3'h3 == state ? tag_0_80 : _GEN_11258; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12288 = 3'h3 == state ? tag_0_81 : _GEN_11259; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12289 = 3'h3 == state ? tag_0_82 : _GEN_11260; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12290 = 3'h3 == state ? tag_0_83 : _GEN_11261; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12291 = 3'h3 == state ? tag_0_84 : _GEN_11262; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12292 = 3'h3 == state ? tag_0_85 : _GEN_11263; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12293 = 3'h3 == state ? tag_0_86 : _GEN_11264; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12294 = 3'h3 == state ? tag_0_87 : _GEN_11265; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12295 = 3'h3 == state ? tag_0_88 : _GEN_11266; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12296 = 3'h3 == state ? tag_0_89 : _GEN_11267; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12297 = 3'h3 == state ? tag_0_90 : _GEN_11268; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12298 = 3'h3 == state ? tag_0_91 : _GEN_11269; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12299 = 3'h3 == state ? tag_0_92 : _GEN_11270; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12300 = 3'h3 == state ? tag_0_93 : _GEN_11271; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12301 = 3'h3 == state ? tag_0_94 : _GEN_11272; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12302 = 3'h3 == state ? tag_0_95 : _GEN_11273; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12303 = 3'h3 == state ? tag_0_96 : _GEN_11274; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12304 = 3'h3 == state ? tag_0_97 : _GEN_11275; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12305 = 3'h3 == state ? tag_0_98 : _GEN_11276; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12306 = 3'h3 == state ? tag_0_99 : _GEN_11277; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12307 = 3'h3 == state ? tag_0_100 : _GEN_11278; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12308 = 3'h3 == state ? tag_0_101 : _GEN_11279; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12309 = 3'h3 == state ? tag_0_102 : _GEN_11280; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12310 = 3'h3 == state ? tag_0_103 : _GEN_11281; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12311 = 3'h3 == state ? tag_0_104 : _GEN_11282; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12312 = 3'h3 == state ? tag_0_105 : _GEN_11283; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12313 = 3'h3 == state ? tag_0_106 : _GEN_11284; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12314 = 3'h3 == state ? tag_0_107 : _GEN_11285; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12315 = 3'h3 == state ? tag_0_108 : _GEN_11286; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12316 = 3'h3 == state ? tag_0_109 : _GEN_11287; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12317 = 3'h3 == state ? tag_0_110 : _GEN_11288; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12318 = 3'h3 == state ? tag_0_111 : _GEN_11289; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12319 = 3'h3 == state ? tag_0_112 : _GEN_11290; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12320 = 3'h3 == state ? tag_0_113 : _GEN_11291; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12321 = 3'h3 == state ? tag_0_114 : _GEN_11292; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12322 = 3'h3 == state ? tag_0_115 : _GEN_11293; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12323 = 3'h3 == state ? tag_0_116 : _GEN_11294; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12324 = 3'h3 == state ? tag_0_117 : _GEN_11295; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12325 = 3'h3 == state ? tag_0_118 : _GEN_11296; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12326 = 3'h3 == state ? tag_0_119 : _GEN_11297; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12327 = 3'h3 == state ? tag_0_120 : _GEN_11298; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12328 = 3'h3 == state ? tag_0_121 : _GEN_11299; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12329 = 3'h3 == state ? tag_0_122 : _GEN_11300; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12330 = 3'h3 == state ? tag_0_123 : _GEN_11301; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12331 = 3'h3 == state ? tag_0_124 : _GEN_11302; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12332 = 3'h3 == state ? tag_0_125 : _GEN_11303; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12333 = 3'h3 == state ? tag_0_126 : _GEN_11304; // @[d_cache.scala 78:18 20:24]
  wire [31:0] _GEN_12334 = 3'h3 == state ? tag_0_127 : _GEN_11305; // @[d_cache.scala 78:18 20:24]
  wire  _GEN_12335 = 3'h3 == state ? valid_0_0 : _GEN_11306; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12336 = 3'h3 == state ? valid_0_1 : _GEN_11307; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12337 = 3'h3 == state ? valid_0_2 : _GEN_11308; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12338 = 3'h3 == state ? valid_0_3 : _GEN_11309; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12339 = 3'h3 == state ? valid_0_4 : _GEN_11310; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12340 = 3'h3 == state ? valid_0_5 : _GEN_11311; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12341 = 3'h3 == state ? valid_0_6 : _GEN_11312; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12342 = 3'h3 == state ? valid_0_7 : _GEN_11313; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12343 = 3'h3 == state ? valid_0_8 : _GEN_11314; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12344 = 3'h3 == state ? valid_0_9 : _GEN_11315; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12345 = 3'h3 == state ? valid_0_10 : _GEN_11316; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12346 = 3'h3 == state ? valid_0_11 : _GEN_11317; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12347 = 3'h3 == state ? valid_0_12 : _GEN_11318; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12348 = 3'h3 == state ? valid_0_13 : _GEN_11319; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12349 = 3'h3 == state ? valid_0_14 : _GEN_11320; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12350 = 3'h3 == state ? valid_0_15 : _GEN_11321; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12351 = 3'h3 == state ? valid_0_16 : _GEN_11322; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12352 = 3'h3 == state ? valid_0_17 : _GEN_11323; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12353 = 3'h3 == state ? valid_0_18 : _GEN_11324; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12354 = 3'h3 == state ? valid_0_19 : _GEN_11325; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12355 = 3'h3 == state ? valid_0_20 : _GEN_11326; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12356 = 3'h3 == state ? valid_0_21 : _GEN_11327; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12357 = 3'h3 == state ? valid_0_22 : _GEN_11328; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12358 = 3'h3 == state ? valid_0_23 : _GEN_11329; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12359 = 3'h3 == state ? valid_0_24 : _GEN_11330; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12360 = 3'h3 == state ? valid_0_25 : _GEN_11331; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12361 = 3'h3 == state ? valid_0_26 : _GEN_11332; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12362 = 3'h3 == state ? valid_0_27 : _GEN_11333; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12363 = 3'h3 == state ? valid_0_28 : _GEN_11334; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12364 = 3'h3 == state ? valid_0_29 : _GEN_11335; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12365 = 3'h3 == state ? valid_0_30 : _GEN_11336; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12366 = 3'h3 == state ? valid_0_31 : _GEN_11337; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12367 = 3'h3 == state ? valid_0_32 : _GEN_11338; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12368 = 3'h3 == state ? valid_0_33 : _GEN_11339; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12369 = 3'h3 == state ? valid_0_34 : _GEN_11340; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12370 = 3'h3 == state ? valid_0_35 : _GEN_11341; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12371 = 3'h3 == state ? valid_0_36 : _GEN_11342; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12372 = 3'h3 == state ? valid_0_37 : _GEN_11343; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12373 = 3'h3 == state ? valid_0_38 : _GEN_11344; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12374 = 3'h3 == state ? valid_0_39 : _GEN_11345; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12375 = 3'h3 == state ? valid_0_40 : _GEN_11346; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12376 = 3'h3 == state ? valid_0_41 : _GEN_11347; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12377 = 3'h3 == state ? valid_0_42 : _GEN_11348; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12378 = 3'h3 == state ? valid_0_43 : _GEN_11349; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12379 = 3'h3 == state ? valid_0_44 : _GEN_11350; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12380 = 3'h3 == state ? valid_0_45 : _GEN_11351; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12381 = 3'h3 == state ? valid_0_46 : _GEN_11352; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12382 = 3'h3 == state ? valid_0_47 : _GEN_11353; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12383 = 3'h3 == state ? valid_0_48 : _GEN_11354; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12384 = 3'h3 == state ? valid_0_49 : _GEN_11355; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12385 = 3'h3 == state ? valid_0_50 : _GEN_11356; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12386 = 3'h3 == state ? valid_0_51 : _GEN_11357; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12387 = 3'h3 == state ? valid_0_52 : _GEN_11358; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12388 = 3'h3 == state ? valid_0_53 : _GEN_11359; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12389 = 3'h3 == state ? valid_0_54 : _GEN_11360; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12390 = 3'h3 == state ? valid_0_55 : _GEN_11361; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12391 = 3'h3 == state ? valid_0_56 : _GEN_11362; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12392 = 3'h3 == state ? valid_0_57 : _GEN_11363; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12393 = 3'h3 == state ? valid_0_58 : _GEN_11364; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12394 = 3'h3 == state ? valid_0_59 : _GEN_11365; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12395 = 3'h3 == state ? valid_0_60 : _GEN_11366; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12396 = 3'h3 == state ? valid_0_61 : _GEN_11367; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12397 = 3'h3 == state ? valid_0_62 : _GEN_11368; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12398 = 3'h3 == state ? valid_0_63 : _GEN_11369; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12399 = 3'h3 == state ? valid_0_64 : _GEN_11370; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12400 = 3'h3 == state ? valid_0_65 : _GEN_11371; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12401 = 3'h3 == state ? valid_0_66 : _GEN_11372; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12402 = 3'h3 == state ? valid_0_67 : _GEN_11373; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12403 = 3'h3 == state ? valid_0_68 : _GEN_11374; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12404 = 3'h3 == state ? valid_0_69 : _GEN_11375; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12405 = 3'h3 == state ? valid_0_70 : _GEN_11376; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12406 = 3'h3 == state ? valid_0_71 : _GEN_11377; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12407 = 3'h3 == state ? valid_0_72 : _GEN_11378; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12408 = 3'h3 == state ? valid_0_73 : _GEN_11379; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12409 = 3'h3 == state ? valid_0_74 : _GEN_11380; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12410 = 3'h3 == state ? valid_0_75 : _GEN_11381; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12411 = 3'h3 == state ? valid_0_76 : _GEN_11382; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12412 = 3'h3 == state ? valid_0_77 : _GEN_11383; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12413 = 3'h3 == state ? valid_0_78 : _GEN_11384; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12414 = 3'h3 == state ? valid_0_79 : _GEN_11385; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12415 = 3'h3 == state ? valid_0_80 : _GEN_11386; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12416 = 3'h3 == state ? valid_0_81 : _GEN_11387; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12417 = 3'h3 == state ? valid_0_82 : _GEN_11388; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12418 = 3'h3 == state ? valid_0_83 : _GEN_11389; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12419 = 3'h3 == state ? valid_0_84 : _GEN_11390; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12420 = 3'h3 == state ? valid_0_85 : _GEN_11391; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12421 = 3'h3 == state ? valid_0_86 : _GEN_11392; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12422 = 3'h3 == state ? valid_0_87 : _GEN_11393; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12423 = 3'h3 == state ? valid_0_88 : _GEN_11394; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12424 = 3'h3 == state ? valid_0_89 : _GEN_11395; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12425 = 3'h3 == state ? valid_0_90 : _GEN_11396; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12426 = 3'h3 == state ? valid_0_91 : _GEN_11397; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12427 = 3'h3 == state ? valid_0_92 : _GEN_11398; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12428 = 3'h3 == state ? valid_0_93 : _GEN_11399; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12429 = 3'h3 == state ? valid_0_94 : _GEN_11400; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12430 = 3'h3 == state ? valid_0_95 : _GEN_11401; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12431 = 3'h3 == state ? valid_0_96 : _GEN_11402; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12432 = 3'h3 == state ? valid_0_97 : _GEN_11403; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12433 = 3'h3 == state ? valid_0_98 : _GEN_11404; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12434 = 3'h3 == state ? valid_0_99 : _GEN_11405; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12435 = 3'h3 == state ? valid_0_100 : _GEN_11406; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12436 = 3'h3 == state ? valid_0_101 : _GEN_11407; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12437 = 3'h3 == state ? valid_0_102 : _GEN_11408; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12438 = 3'h3 == state ? valid_0_103 : _GEN_11409; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12439 = 3'h3 == state ? valid_0_104 : _GEN_11410; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12440 = 3'h3 == state ? valid_0_105 : _GEN_11411; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12441 = 3'h3 == state ? valid_0_106 : _GEN_11412; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12442 = 3'h3 == state ? valid_0_107 : _GEN_11413; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12443 = 3'h3 == state ? valid_0_108 : _GEN_11414; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12444 = 3'h3 == state ? valid_0_109 : _GEN_11415; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12445 = 3'h3 == state ? valid_0_110 : _GEN_11416; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12446 = 3'h3 == state ? valid_0_111 : _GEN_11417; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12447 = 3'h3 == state ? valid_0_112 : _GEN_11418; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12448 = 3'h3 == state ? valid_0_113 : _GEN_11419; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12449 = 3'h3 == state ? valid_0_114 : _GEN_11420; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12450 = 3'h3 == state ? valid_0_115 : _GEN_11421; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12451 = 3'h3 == state ? valid_0_116 : _GEN_11422; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12452 = 3'h3 == state ? valid_0_117 : _GEN_11423; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12453 = 3'h3 == state ? valid_0_118 : _GEN_11424; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12454 = 3'h3 == state ? valid_0_119 : _GEN_11425; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12455 = 3'h3 == state ? valid_0_120 : _GEN_11426; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12456 = 3'h3 == state ? valid_0_121 : _GEN_11427; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12457 = 3'h3 == state ? valid_0_122 : _GEN_11428; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12458 = 3'h3 == state ? valid_0_123 : _GEN_11429; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12459 = 3'h3 == state ? valid_0_124 : _GEN_11430; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12460 = 3'h3 == state ? valid_0_125 : _GEN_11431; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12461 = 3'h3 == state ? valid_0_126 : _GEN_11432; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12462 = 3'h3 == state ? valid_0_127 : _GEN_11433; // @[d_cache.scala 78:18 22:26]
  wire  _GEN_12463 = 3'h3 == state ? quene : _GEN_11434; // @[d_cache.scala 78:18 35:24]
  wire [63:0] _GEN_12464 = 3'h3 == state ? ram_1_0 : _GEN_11435; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12465 = 3'h3 == state ? ram_1_1 : _GEN_11436; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12466 = 3'h3 == state ? ram_1_2 : _GEN_11437; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12467 = 3'h3 == state ? ram_1_3 : _GEN_11438; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12468 = 3'h3 == state ? ram_1_4 : _GEN_11439; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12469 = 3'h3 == state ? ram_1_5 : _GEN_11440; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12470 = 3'h3 == state ? ram_1_6 : _GEN_11441; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12471 = 3'h3 == state ? ram_1_7 : _GEN_11442; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12472 = 3'h3 == state ? ram_1_8 : _GEN_11443; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12473 = 3'h3 == state ? ram_1_9 : _GEN_11444; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12474 = 3'h3 == state ? ram_1_10 : _GEN_11445; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12475 = 3'h3 == state ? ram_1_11 : _GEN_11446; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12476 = 3'h3 == state ? ram_1_12 : _GEN_11447; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12477 = 3'h3 == state ? ram_1_13 : _GEN_11448; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12478 = 3'h3 == state ? ram_1_14 : _GEN_11449; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12479 = 3'h3 == state ? ram_1_15 : _GEN_11450; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12480 = 3'h3 == state ? ram_1_16 : _GEN_11451; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12481 = 3'h3 == state ? ram_1_17 : _GEN_11452; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12482 = 3'h3 == state ? ram_1_18 : _GEN_11453; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12483 = 3'h3 == state ? ram_1_19 : _GEN_11454; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12484 = 3'h3 == state ? ram_1_20 : _GEN_11455; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12485 = 3'h3 == state ? ram_1_21 : _GEN_11456; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12486 = 3'h3 == state ? ram_1_22 : _GEN_11457; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12487 = 3'h3 == state ? ram_1_23 : _GEN_11458; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12488 = 3'h3 == state ? ram_1_24 : _GEN_11459; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12489 = 3'h3 == state ? ram_1_25 : _GEN_11460; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12490 = 3'h3 == state ? ram_1_26 : _GEN_11461; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12491 = 3'h3 == state ? ram_1_27 : _GEN_11462; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12492 = 3'h3 == state ? ram_1_28 : _GEN_11463; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12493 = 3'h3 == state ? ram_1_29 : _GEN_11464; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12494 = 3'h3 == state ? ram_1_30 : _GEN_11465; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12495 = 3'h3 == state ? ram_1_31 : _GEN_11466; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12496 = 3'h3 == state ? ram_1_32 : _GEN_11467; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12497 = 3'h3 == state ? ram_1_33 : _GEN_11468; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12498 = 3'h3 == state ? ram_1_34 : _GEN_11469; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12499 = 3'h3 == state ? ram_1_35 : _GEN_11470; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12500 = 3'h3 == state ? ram_1_36 : _GEN_11471; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12501 = 3'h3 == state ? ram_1_37 : _GEN_11472; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12502 = 3'h3 == state ? ram_1_38 : _GEN_11473; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12503 = 3'h3 == state ? ram_1_39 : _GEN_11474; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12504 = 3'h3 == state ? ram_1_40 : _GEN_11475; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12505 = 3'h3 == state ? ram_1_41 : _GEN_11476; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12506 = 3'h3 == state ? ram_1_42 : _GEN_11477; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12507 = 3'h3 == state ? ram_1_43 : _GEN_11478; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12508 = 3'h3 == state ? ram_1_44 : _GEN_11479; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12509 = 3'h3 == state ? ram_1_45 : _GEN_11480; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12510 = 3'h3 == state ? ram_1_46 : _GEN_11481; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12511 = 3'h3 == state ? ram_1_47 : _GEN_11482; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12512 = 3'h3 == state ? ram_1_48 : _GEN_11483; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12513 = 3'h3 == state ? ram_1_49 : _GEN_11484; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12514 = 3'h3 == state ? ram_1_50 : _GEN_11485; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12515 = 3'h3 == state ? ram_1_51 : _GEN_11486; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12516 = 3'h3 == state ? ram_1_52 : _GEN_11487; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12517 = 3'h3 == state ? ram_1_53 : _GEN_11488; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12518 = 3'h3 == state ? ram_1_54 : _GEN_11489; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12519 = 3'h3 == state ? ram_1_55 : _GEN_11490; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12520 = 3'h3 == state ? ram_1_56 : _GEN_11491; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12521 = 3'h3 == state ? ram_1_57 : _GEN_11492; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12522 = 3'h3 == state ? ram_1_58 : _GEN_11493; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12523 = 3'h3 == state ? ram_1_59 : _GEN_11494; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12524 = 3'h3 == state ? ram_1_60 : _GEN_11495; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12525 = 3'h3 == state ? ram_1_61 : _GEN_11496; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12526 = 3'h3 == state ? ram_1_62 : _GEN_11497; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12527 = 3'h3 == state ? ram_1_63 : _GEN_11498; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12528 = 3'h3 == state ? ram_1_64 : _GEN_11499; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12529 = 3'h3 == state ? ram_1_65 : _GEN_11500; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12530 = 3'h3 == state ? ram_1_66 : _GEN_11501; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12531 = 3'h3 == state ? ram_1_67 : _GEN_11502; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12532 = 3'h3 == state ? ram_1_68 : _GEN_11503; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12533 = 3'h3 == state ? ram_1_69 : _GEN_11504; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12534 = 3'h3 == state ? ram_1_70 : _GEN_11505; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12535 = 3'h3 == state ? ram_1_71 : _GEN_11506; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12536 = 3'h3 == state ? ram_1_72 : _GEN_11507; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12537 = 3'h3 == state ? ram_1_73 : _GEN_11508; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12538 = 3'h3 == state ? ram_1_74 : _GEN_11509; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12539 = 3'h3 == state ? ram_1_75 : _GEN_11510; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12540 = 3'h3 == state ? ram_1_76 : _GEN_11511; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12541 = 3'h3 == state ? ram_1_77 : _GEN_11512; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12542 = 3'h3 == state ? ram_1_78 : _GEN_11513; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12543 = 3'h3 == state ? ram_1_79 : _GEN_11514; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12544 = 3'h3 == state ? ram_1_80 : _GEN_11515; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12545 = 3'h3 == state ? ram_1_81 : _GEN_11516; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12546 = 3'h3 == state ? ram_1_82 : _GEN_11517; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12547 = 3'h3 == state ? ram_1_83 : _GEN_11518; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12548 = 3'h3 == state ? ram_1_84 : _GEN_11519; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12549 = 3'h3 == state ? ram_1_85 : _GEN_11520; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12550 = 3'h3 == state ? ram_1_86 : _GEN_11521; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12551 = 3'h3 == state ? ram_1_87 : _GEN_11522; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12552 = 3'h3 == state ? ram_1_88 : _GEN_11523; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12553 = 3'h3 == state ? ram_1_89 : _GEN_11524; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12554 = 3'h3 == state ? ram_1_90 : _GEN_11525; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12555 = 3'h3 == state ? ram_1_91 : _GEN_11526; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12556 = 3'h3 == state ? ram_1_92 : _GEN_11527; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12557 = 3'h3 == state ? ram_1_93 : _GEN_11528; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12558 = 3'h3 == state ? ram_1_94 : _GEN_11529; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12559 = 3'h3 == state ? ram_1_95 : _GEN_11530; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12560 = 3'h3 == state ? ram_1_96 : _GEN_11531; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12561 = 3'h3 == state ? ram_1_97 : _GEN_11532; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12562 = 3'h3 == state ? ram_1_98 : _GEN_11533; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12563 = 3'h3 == state ? ram_1_99 : _GEN_11534; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12564 = 3'h3 == state ? ram_1_100 : _GEN_11535; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12565 = 3'h3 == state ? ram_1_101 : _GEN_11536; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12566 = 3'h3 == state ? ram_1_102 : _GEN_11537; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12567 = 3'h3 == state ? ram_1_103 : _GEN_11538; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12568 = 3'h3 == state ? ram_1_104 : _GEN_11539; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12569 = 3'h3 == state ? ram_1_105 : _GEN_11540; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12570 = 3'h3 == state ? ram_1_106 : _GEN_11541; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12571 = 3'h3 == state ? ram_1_107 : _GEN_11542; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12572 = 3'h3 == state ? ram_1_108 : _GEN_11543; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12573 = 3'h3 == state ? ram_1_109 : _GEN_11544; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12574 = 3'h3 == state ? ram_1_110 : _GEN_11545; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12575 = 3'h3 == state ? ram_1_111 : _GEN_11546; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12576 = 3'h3 == state ? ram_1_112 : _GEN_11547; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12577 = 3'h3 == state ? ram_1_113 : _GEN_11548; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12578 = 3'h3 == state ? ram_1_114 : _GEN_11549; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12579 = 3'h3 == state ? ram_1_115 : _GEN_11550; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12580 = 3'h3 == state ? ram_1_116 : _GEN_11551; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12581 = 3'h3 == state ? ram_1_117 : _GEN_11552; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12582 = 3'h3 == state ? ram_1_118 : _GEN_11553; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12583 = 3'h3 == state ? ram_1_119 : _GEN_11554; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12584 = 3'h3 == state ? ram_1_120 : _GEN_11555; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12585 = 3'h3 == state ? ram_1_121 : _GEN_11556; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12586 = 3'h3 == state ? ram_1_122 : _GEN_11557; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12587 = 3'h3 == state ? ram_1_123 : _GEN_11558; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12588 = 3'h3 == state ? ram_1_124 : _GEN_11559; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12589 = 3'h3 == state ? ram_1_125 : _GEN_11560; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12590 = 3'h3 == state ? ram_1_126 : _GEN_11561; // @[d_cache.scala 78:18 19:24]
  wire [63:0] _GEN_12591 = 3'h3 == state ? ram_1_127 : _GEN_11562; // @[d_cache.scala 78:18 19:24]
  wire [31:0] _GEN_12592 = 3'h3 == state ? tag_1_0 : _GEN_11563; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12593 = 3'h3 == state ? tag_1_1 : _GEN_11564; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12594 = 3'h3 == state ? tag_1_2 : _GEN_11565; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12595 = 3'h3 == state ? tag_1_3 : _GEN_11566; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12596 = 3'h3 == state ? tag_1_4 : _GEN_11567; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12597 = 3'h3 == state ? tag_1_5 : _GEN_11568; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12598 = 3'h3 == state ? tag_1_6 : _GEN_11569; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12599 = 3'h3 == state ? tag_1_7 : _GEN_11570; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12600 = 3'h3 == state ? tag_1_8 : _GEN_11571; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12601 = 3'h3 == state ? tag_1_9 : _GEN_11572; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12602 = 3'h3 == state ? tag_1_10 : _GEN_11573; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12603 = 3'h3 == state ? tag_1_11 : _GEN_11574; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12604 = 3'h3 == state ? tag_1_12 : _GEN_11575; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12605 = 3'h3 == state ? tag_1_13 : _GEN_11576; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12606 = 3'h3 == state ? tag_1_14 : _GEN_11577; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12607 = 3'h3 == state ? tag_1_15 : _GEN_11578; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12608 = 3'h3 == state ? tag_1_16 : _GEN_11579; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12609 = 3'h3 == state ? tag_1_17 : _GEN_11580; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12610 = 3'h3 == state ? tag_1_18 : _GEN_11581; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12611 = 3'h3 == state ? tag_1_19 : _GEN_11582; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12612 = 3'h3 == state ? tag_1_20 : _GEN_11583; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12613 = 3'h3 == state ? tag_1_21 : _GEN_11584; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12614 = 3'h3 == state ? tag_1_22 : _GEN_11585; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12615 = 3'h3 == state ? tag_1_23 : _GEN_11586; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12616 = 3'h3 == state ? tag_1_24 : _GEN_11587; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12617 = 3'h3 == state ? tag_1_25 : _GEN_11588; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12618 = 3'h3 == state ? tag_1_26 : _GEN_11589; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12619 = 3'h3 == state ? tag_1_27 : _GEN_11590; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12620 = 3'h3 == state ? tag_1_28 : _GEN_11591; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12621 = 3'h3 == state ? tag_1_29 : _GEN_11592; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12622 = 3'h3 == state ? tag_1_30 : _GEN_11593; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12623 = 3'h3 == state ? tag_1_31 : _GEN_11594; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12624 = 3'h3 == state ? tag_1_32 : _GEN_11595; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12625 = 3'h3 == state ? tag_1_33 : _GEN_11596; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12626 = 3'h3 == state ? tag_1_34 : _GEN_11597; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12627 = 3'h3 == state ? tag_1_35 : _GEN_11598; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12628 = 3'h3 == state ? tag_1_36 : _GEN_11599; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12629 = 3'h3 == state ? tag_1_37 : _GEN_11600; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12630 = 3'h3 == state ? tag_1_38 : _GEN_11601; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12631 = 3'h3 == state ? tag_1_39 : _GEN_11602; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12632 = 3'h3 == state ? tag_1_40 : _GEN_11603; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12633 = 3'h3 == state ? tag_1_41 : _GEN_11604; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12634 = 3'h3 == state ? tag_1_42 : _GEN_11605; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12635 = 3'h3 == state ? tag_1_43 : _GEN_11606; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12636 = 3'h3 == state ? tag_1_44 : _GEN_11607; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12637 = 3'h3 == state ? tag_1_45 : _GEN_11608; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12638 = 3'h3 == state ? tag_1_46 : _GEN_11609; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12639 = 3'h3 == state ? tag_1_47 : _GEN_11610; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12640 = 3'h3 == state ? tag_1_48 : _GEN_11611; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12641 = 3'h3 == state ? tag_1_49 : _GEN_11612; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12642 = 3'h3 == state ? tag_1_50 : _GEN_11613; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12643 = 3'h3 == state ? tag_1_51 : _GEN_11614; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12644 = 3'h3 == state ? tag_1_52 : _GEN_11615; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12645 = 3'h3 == state ? tag_1_53 : _GEN_11616; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12646 = 3'h3 == state ? tag_1_54 : _GEN_11617; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12647 = 3'h3 == state ? tag_1_55 : _GEN_11618; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12648 = 3'h3 == state ? tag_1_56 : _GEN_11619; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12649 = 3'h3 == state ? tag_1_57 : _GEN_11620; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12650 = 3'h3 == state ? tag_1_58 : _GEN_11621; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12651 = 3'h3 == state ? tag_1_59 : _GEN_11622; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12652 = 3'h3 == state ? tag_1_60 : _GEN_11623; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12653 = 3'h3 == state ? tag_1_61 : _GEN_11624; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12654 = 3'h3 == state ? tag_1_62 : _GEN_11625; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12655 = 3'h3 == state ? tag_1_63 : _GEN_11626; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12656 = 3'h3 == state ? tag_1_64 : _GEN_11627; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12657 = 3'h3 == state ? tag_1_65 : _GEN_11628; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12658 = 3'h3 == state ? tag_1_66 : _GEN_11629; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12659 = 3'h3 == state ? tag_1_67 : _GEN_11630; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12660 = 3'h3 == state ? tag_1_68 : _GEN_11631; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12661 = 3'h3 == state ? tag_1_69 : _GEN_11632; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12662 = 3'h3 == state ? tag_1_70 : _GEN_11633; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12663 = 3'h3 == state ? tag_1_71 : _GEN_11634; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12664 = 3'h3 == state ? tag_1_72 : _GEN_11635; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12665 = 3'h3 == state ? tag_1_73 : _GEN_11636; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12666 = 3'h3 == state ? tag_1_74 : _GEN_11637; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12667 = 3'h3 == state ? tag_1_75 : _GEN_11638; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12668 = 3'h3 == state ? tag_1_76 : _GEN_11639; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12669 = 3'h3 == state ? tag_1_77 : _GEN_11640; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12670 = 3'h3 == state ? tag_1_78 : _GEN_11641; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12671 = 3'h3 == state ? tag_1_79 : _GEN_11642; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12672 = 3'h3 == state ? tag_1_80 : _GEN_11643; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12673 = 3'h3 == state ? tag_1_81 : _GEN_11644; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12674 = 3'h3 == state ? tag_1_82 : _GEN_11645; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12675 = 3'h3 == state ? tag_1_83 : _GEN_11646; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12676 = 3'h3 == state ? tag_1_84 : _GEN_11647; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12677 = 3'h3 == state ? tag_1_85 : _GEN_11648; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12678 = 3'h3 == state ? tag_1_86 : _GEN_11649; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12679 = 3'h3 == state ? tag_1_87 : _GEN_11650; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12680 = 3'h3 == state ? tag_1_88 : _GEN_11651; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12681 = 3'h3 == state ? tag_1_89 : _GEN_11652; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12682 = 3'h3 == state ? tag_1_90 : _GEN_11653; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12683 = 3'h3 == state ? tag_1_91 : _GEN_11654; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12684 = 3'h3 == state ? tag_1_92 : _GEN_11655; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12685 = 3'h3 == state ? tag_1_93 : _GEN_11656; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12686 = 3'h3 == state ? tag_1_94 : _GEN_11657; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12687 = 3'h3 == state ? tag_1_95 : _GEN_11658; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12688 = 3'h3 == state ? tag_1_96 : _GEN_11659; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12689 = 3'h3 == state ? tag_1_97 : _GEN_11660; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12690 = 3'h3 == state ? tag_1_98 : _GEN_11661; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12691 = 3'h3 == state ? tag_1_99 : _GEN_11662; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12692 = 3'h3 == state ? tag_1_100 : _GEN_11663; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12693 = 3'h3 == state ? tag_1_101 : _GEN_11664; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12694 = 3'h3 == state ? tag_1_102 : _GEN_11665; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12695 = 3'h3 == state ? tag_1_103 : _GEN_11666; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12696 = 3'h3 == state ? tag_1_104 : _GEN_11667; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12697 = 3'h3 == state ? tag_1_105 : _GEN_11668; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12698 = 3'h3 == state ? tag_1_106 : _GEN_11669; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12699 = 3'h3 == state ? tag_1_107 : _GEN_11670; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12700 = 3'h3 == state ? tag_1_108 : _GEN_11671; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12701 = 3'h3 == state ? tag_1_109 : _GEN_11672; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12702 = 3'h3 == state ? tag_1_110 : _GEN_11673; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12703 = 3'h3 == state ? tag_1_111 : _GEN_11674; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12704 = 3'h3 == state ? tag_1_112 : _GEN_11675; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12705 = 3'h3 == state ? tag_1_113 : _GEN_11676; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12706 = 3'h3 == state ? tag_1_114 : _GEN_11677; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12707 = 3'h3 == state ? tag_1_115 : _GEN_11678; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12708 = 3'h3 == state ? tag_1_116 : _GEN_11679; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12709 = 3'h3 == state ? tag_1_117 : _GEN_11680; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12710 = 3'h3 == state ? tag_1_118 : _GEN_11681; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12711 = 3'h3 == state ? tag_1_119 : _GEN_11682; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12712 = 3'h3 == state ? tag_1_120 : _GEN_11683; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12713 = 3'h3 == state ? tag_1_121 : _GEN_11684; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12714 = 3'h3 == state ? tag_1_122 : _GEN_11685; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12715 = 3'h3 == state ? tag_1_123 : _GEN_11686; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12716 = 3'h3 == state ? tag_1_124 : _GEN_11687; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12717 = 3'h3 == state ? tag_1_125 : _GEN_11688; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12718 = 3'h3 == state ? tag_1_126 : _GEN_11689; // @[d_cache.scala 78:18 21:24]
  wire [31:0] _GEN_12719 = 3'h3 == state ? tag_1_127 : _GEN_11690; // @[d_cache.scala 78:18 21:24]
  wire  _GEN_12720 = 3'h3 == state ? valid_1_0 : _GEN_11691; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12721 = 3'h3 == state ? valid_1_1 : _GEN_11692; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12722 = 3'h3 == state ? valid_1_2 : _GEN_11693; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12723 = 3'h3 == state ? valid_1_3 : _GEN_11694; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12724 = 3'h3 == state ? valid_1_4 : _GEN_11695; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12725 = 3'h3 == state ? valid_1_5 : _GEN_11696; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12726 = 3'h3 == state ? valid_1_6 : _GEN_11697; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12727 = 3'h3 == state ? valid_1_7 : _GEN_11698; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12728 = 3'h3 == state ? valid_1_8 : _GEN_11699; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12729 = 3'h3 == state ? valid_1_9 : _GEN_11700; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12730 = 3'h3 == state ? valid_1_10 : _GEN_11701; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12731 = 3'h3 == state ? valid_1_11 : _GEN_11702; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12732 = 3'h3 == state ? valid_1_12 : _GEN_11703; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12733 = 3'h3 == state ? valid_1_13 : _GEN_11704; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12734 = 3'h3 == state ? valid_1_14 : _GEN_11705; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12735 = 3'h3 == state ? valid_1_15 : _GEN_11706; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12736 = 3'h3 == state ? valid_1_16 : _GEN_11707; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12737 = 3'h3 == state ? valid_1_17 : _GEN_11708; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12738 = 3'h3 == state ? valid_1_18 : _GEN_11709; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12739 = 3'h3 == state ? valid_1_19 : _GEN_11710; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12740 = 3'h3 == state ? valid_1_20 : _GEN_11711; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12741 = 3'h3 == state ? valid_1_21 : _GEN_11712; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12742 = 3'h3 == state ? valid_1_22 : _GEN_11713; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12743 = 3'h3 == state ? valid_1_23 : _GEN_11714; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12744 = 3'h3 == state ? valid_1_24 : _GEN_11715; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12745 = 3'h3 == state ? valid_1_25 : _GEN_11716; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12746 = 3'h3 == state ? valid_1_26 : _GEN_11717; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12747 = 3'h3 == state ? valid_1_27 : _GEN_11718; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12748 = 3'h3 == state ? valid_1_28 : _GEN_11719; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12749 = 3'h3 == state ? valid_1_29 : _GEN_11720; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12750 = 3'h3 == state ? valid_1_30 : _GEN_11721; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12751 = 3'h3 == state ? valid_1_31 : _GEN_11722; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12752 = 3'h3 == state ? valid_1_32 : _GEN_11723; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12753 = 3'h3 == state ? valid_1_33 : _GEN_11724; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12754 = 3'h3 == state ? valid_1_34 : _GEN_11725; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12755 = 3'h3 == state ? valid_1_35 : _GEN_11726; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12756 = 3'h3 == state ? valid_1_36 : _GEN_11727; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12757 = 3'h3 == state ? valid_1_37 : _GEN_11728; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12758 = 3'h3 == state ? valid_1_38 : _GEN_11729; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12759 = 3'h3 == state ? valid_1_39 : _GEN_11730; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12760 = 3'h3 == state ? valid_1_40 : _GEN_11731; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12761 = 3'h3 == state ? valid_1_41 : _GEN_11732; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12762 = 3'h3 == state ? valid_1_42 : _GEN_11733; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12763 = 3'h3 == state ? valid_1_43 : _GEN_11734; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12764 = 3'h3 == state ? valid_1_44 : _GEN_11735; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12765 = 3'h3 == state ? valid_1_45 : _GEN_11736; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12766 = 3'h3 == state ? valid_1_46 : _GEN_11737; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12767 = 3'h3 == state ? valid_1_47 : _GEN_11738; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12768 = 3'h3 == state ? valid_1_48 : _GEN_11739; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12769 = 3'h3 == state ? valid_1_49 : _GEN_11740; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12770 = 3'h3 == state ? valid_1_50 : _GEN_11741; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12771 = 3'h3 == state ? valid_1_51 : _GEN_11742; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12772 = 3'h3 == state ? valid_1_52 : _GEN_11743; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12773 = 3'h3 == state ? valid_1_53 : _GEN_11744; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12774 = 3'h3 == state ? valid_1_54 : _GEN_11745; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12775 = 3'h3 == state ? valid_1_55 : _GEN_11746; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12776 = 3'h3 == state ? valid_1_56 : _GEN_11747; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12777 = 3'h3 == state ? valid_1_57 : _GEN_11748; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12778 = 3'h3 == state ? valid_1_58 : _GEN_11749; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12779 = 3'h3 == state ? valid_1_59 : _GEN_11750; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12780 = 3'h3 == state ? valid_1_60 : _GEN_11751; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12781 = 3'h3 == state ? valid_1_61 : _GEN_11752; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12782 = 3'h3 == state ? valid_1_62 : _GEN_11753; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12783 = 3'h3 == state ? valid_1_63 : _GEN_11754; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12784 = 3'h3 == state ? valid_1_64 : _GEN_11755; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12785 = 3'h3 == state ? valid_1_65 : _GEN_11756; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12786 = 3'h3 == state ? valid_1_66 : _GEN_11757; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12787 = 3'h3 == state ? valid_1_67 : _GEN_11758; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12788 = 3'h3 == state ? valid_1_68 : _GEN_11759; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12789 = 3'h3 == state ? valid_1_69 : _GEN_11760; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12790 = 3'h3 == state ? valid_1_70 : _GEN_11761; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12791 = 3'h3 == state ? valid_1_71 : _GEN_11762; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12792 = 3'h3 == state ? valid_1_72 : _GEN_11763; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12793 = 3'h3 == state ? valid_1_73 : _GEN_11764; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12794 = 3'h3 == state ? valid_1_74 : _GEN_11765; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12795 = 3'h3 == state ? valid_1_75 : _GEN_11766; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12796 = 3'h3 == state ? valid_1_76 : _GEN_11767; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12797 = 3'h3 == state ? valid_1_77 : _GEN_11768; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12798 = 3'h3 == state ? valid_1_78 : _GEN_11769; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12799 = 3'h3 == state ? valid_1_79 : _GEN_11770; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12800 = 3'h3 == state ? valid_1_80 : _GEN_11771; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12801 = 3'h3 == state ? valid_1_81 : _GEN_11772; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12802 = 3'h3 == state ? valid_1_82 : _GEN_11773; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12803 = 3'h3 == state ? valid_1_83 : _GEN_11774; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12804 = 3'h3 == state ? valid_1_84 : _GEN_11775; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12805 = 3'h3 == state ? valid_1_85 : _GEN_11776; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12806 = 3'h3 == state ? valid_1_86 : _GEN_11777; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12807 = 3'h3 == state ? valid_1_87 : _GEN_11778; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12808 = 3'h3 == state ? valid_1_88 : _GEN_11779; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12809 = 3'h3 == state ? valid_1_89 : _GEN_11780; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12810 = 3'h3 == state ? valid_1_90 : _GEN_11781; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12811 = 3'h3 == state ? valid_1_91 : _GEN_11782; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12812 = 3'h3 == state ? valid_1_92 : _GEN_11783; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12813 = 3'h3 == state ? valid_1_93 : _GEN_11784; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12814 = 3'h3 == state ? valid_1_94 : _GEN_11785; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12815 = 3'h3 == state ? valid_1_95 : _GEN_11786; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12816 = 3'h3 == state ? valid_1_96 : _GEN_11787; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12817 = 3'h3 == state ? valid_1_97 : _GEN_11788; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12818 = 3'h3 == state ? valid_1_98 : _GEN_11789; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12819 = 3'h3 == state ? valid_1_99 : _GEN_11790; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12820 = 3'h3 == state ? valid_1_100 : _GEN_11791; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12821 = 3'h3 == state ? valid_1_101 : _GEN_11792; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12822 = 3'h3 == state ? valid_1_102 : _GEN_11793; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12823 = 3'h3 == state ? valid_1_103 : _GEN_11794; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12824 = 3'h3 == state ? valid_1_104 : _GEN_11795; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12825 = 3'h3 == state ? valid_1_105 : _GEN_11796; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12826 = 3'h3 == state ? valid_1_106 : _GEN_11797; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12827 = 3'h3 == state ? valid_1_107 : _GEN_11798; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12828 = 3'h3 == state ? valid_1_108 : _GEN_11799; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12829 = 3'h3 == state ? valid_1_109 : _GEN_11800; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12830 = 3'h3 == state ? valid_1_110 : _GEN_11801; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12831 = 3'h3 == state ? valid_1_111 : _GEN_11802; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12832 = 3'h3 == state ? valid_1_112 : _GEN_11803; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12833 = 3'h3 == state ? valid_1_113 : _GEN_11804; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12834 = 3'h3 == state ? valid_1_114 : _GEN_11805; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12835 = 3'h3 == state ? valid_1_115 : _GEN_11806; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12836 = 3'h3 == state ? valid_1_116 : _GEN_11807; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12837 = 3'h3 == state ? valid_1_117 : _GEN_11808; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12838 = 3'h3 == state ? valid_1_118 : _GEN_11809; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12839 = 3'h3 == state ? valid_1_119 : _GEN_11810; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12840 = 3'h3 == state ? valid_1_120 : _GEN_11811; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12841 = 3'h3 == state ? valid_1_121 : _GEN_11812; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12842 = 3'h3 == state ? valid_1_122 : _GEN_11813; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12843 = 3'h3 == state ? valid_1_123 : _GEN_11814; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12844 = 3'h3 == state ? valid_1_124 : _GEN_11815; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12845 = 3'h3 == state ? valid_1_125 : _GEN_11816; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12846 = 3'h3 == state ? valid_1_126 : _GEN_11817; // @[d_cache.scala 78:18 23:26]
  wire  _GEN_12847 = 3'h3 == state ? valid_1_127 : _GEN_11818; // @[d_cache.scala 78:18 23:26]
  wire [63:0] _GEN_12848 = 3'h3 == state ? write_back_data : _GEN_11819; // @[d_cache.scala 78:18 29:34]
  wire [41:0] _GEN_12849 = 3'h3 == state ? {{10'd0}, write_back_addr} : _GEN_11820; // @[d_cache.scala 78:18 30:34]
  wire  _GEN_12850 = 3'h3 == state ? dirty_0_0 : _GEN_11821; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12851 = 3'h3 == state ? dirty_0_1 : _GEN_11822; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12852 = 3'h3 == state ? dirty_0_2 : _GEN_11823; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12853 = 3'h3 == state ? dirty_0_3 : _GEN_11824; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12854 = 3'h3 == state ? dirty_0_4 : _GEN_11825; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12855 = 3'h3 == state ? dirty_0_5 : _GEN_11826; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12856 = 3'h3 == state ? dirty_0_6 : _GEN_11827; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12857 = 3'h3 == state ? dirty_0_7 : _GEN_11828; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12858 = 3'h3 == state ? dirty_0_8 : _GEN_11829; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12859 = 3'h3 == state ? dirty_0_9 : _GEN_11830; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12860 = 3'h3 == state ? dirty_0_10 : _GEN_11831; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12861 = 3'h3 == state ? dirty_0_11 : _GEN_11832; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12862 = 3'h3 == state ? dirty_0_12 : _GEN_11833; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12863 = 3'h3 == state ? dirty_0_13 : _GEN_11834; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12864 = 3'h3 == state ? dirty_0_14 : _GEN_11835; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12865 = 3'h3 == state ? dirty_0_15 : _GEN_11836; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12866 = 3'h3 == state ? dirty_0_16 : _GEN_11837; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12867 = 3'h3 == state ? dirty_0_17 : _GEN_11838; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12868 = 3'h3 == state ? dirty_0_18 : _GEN_11839; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12869 = 3'h3 == state ? dirty_0_19 : _GEN_11840; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12870 = 3'h3 == state ? dirty_0_20 : _GEN_11841; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12871 = 3'h3 == state ? dirty_0_21 : _GEN_11842; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12872 = 3'h3 == state ? dirty_0_22 : _GEN_11843; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12873 = 3'h3 == state ? dirty_0_23 : _GEN_11844; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12874 = 3'h3 == state ? dirty_0_24 : _GEN_11845; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12875 = 3'h3 == state ? dirty_0_25 : _GEN_11846; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12876 = 3'h3 == state ? dirty_0_26 : _GEN_11847; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12877 = 3'h3 == state ? dirty_0_27 : _GEN_11848; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12878 = 3'h3 == state ? dirty_0_28 : _GEN_11849; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12879 = 3'h3 == state ? dirty_0_29 : _GEN_11850; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12880 = 3'h3 == state ? dirty_0_30 : _GEN_11851; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12881 = 3'h3 == state ? dirty_0_31 : _GEN_11852; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12882 = 3'h3 == state ? dirty_0_32 : _GEN_11853; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12883 = 3'h3 == state ? dirty_0_33 : _GEN_11854; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12884 = 3'h3 == state ? dirty_0_34 : _GEN_11855; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12885 = 3'h3 == state ? dirty_0_35 : _GEN_11856; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12886 = 3'h3 == state ? dirty_0_36 : _GEN_11857; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12887 = 3'h3 == state ? dirty_0_37 : _GEN_11858; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12888 = 3'h3 == state ? dirty_0_38 : _GEN_11859; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12889 = 3'h3 == state ? dirty_0_39 : _GEN_11860; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12890 = 3'h3 == state ? dirty_0_40 : _GEN_11861; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12891 = 3'h3 == state ? dirty_0_41 : _GEN_11862; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12892 = 3'h3 == state ? dirty_0_42 : _GEN_11863; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12893 = 3'h3 == state ? dirty_0_43 : _GEN_11864; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12894 = 3'h3 == state ? dirty_0_44 : _GEN_11865; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12895 = 3'h3 == state ? dirty_0_45 : _GEN_11866; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12896 = 3'h3 == state ? dirty_0_46 : _GEN_11867; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12897 = 3'h3 == state ? dirty_0_47 : _GEN_11868; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12898 = 3'h3 == state ? dirty_0_48 : _GEN_11869; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12899 = 3'h3 == state ? dirty_0_49 : _GEN_11870; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12900 = 3'h3 == state ? dirty_0_50 : _GEN_11871; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12901 = 3'h3 == state ? dirty_0_51 : _GEN_11872; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12902 = 3'h3 == state ? dirty_0_52 : _GEN_11873; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12903 = 3'h3 == state ? dirty_0_53 : _GEN_11874; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12904 = 3'h3 == state ? dirty_0_54 : _GEN_11875; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12905 = 3'h3 == state ? dirty_0_55 : _GEN_11876; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12906 = 3'h3 == state ? dirty_0_56 : _GEN_11877; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12907 = 3'h3 == state ? dirty_0_57 : _GEN_11878; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12908 = 3'h3 == state ? dirty_0_58 : _GEN_11879; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12909 = 3'h3 == state ? dirty_0_59 : _GEN_11880; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12910 = 3'h3 == state ? dirty_0_60 : _GEN_11881; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12911 = 3'h3 == state ? dirty_0_61 : _GEN_11882; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12912 = 3'h3 == state ? dirty_0_62 : _GEN_11883; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12913 = 3'h3 == state ? dirty_0_63 : _GEN_11884; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12914 = 3'h3 == state ? dirty_0_64 : _GEN_11885; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12915 = 3'h3 == state ? dirty_0_65 : _GEN_11886; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12916 = 3'h3 == state ? dirty_0_66 : _GEN_11887; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12917 = 3'h3 == state ? dirty_0_67 : _GEN_11888; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12918 = 3'h3 == state ? dirty_0_68 : _GEN_11889; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12919 = 3'h3 == state ? dirty_0_69 : _GEN_11890; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12920 = 3'h3 == state ? dirty_0_70 : _GEN_11891; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12921 = 3'h3 == state ? dirty_0_71 : _GEN_11892; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12922 = 3'h3 == state ? dirty_0_72 : _GEN_11893; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12923 = 3'h3 == state ? dirty_0_73 : _GEN_11894; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12924 = 3'h3 == state ? dirty_0_74 : _GEN_11895; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12925 = 3'h3 == state ? dirty_0_75 : _GEN_11896; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12926 = 3'h3 == state ? dirty_0_76 : _GEN_11897; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12927 = 3'h3 == state ? dirty_0_77 : _GEN_11898; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12928 = 3'h3 == state ? dirty_0_78 : _GEN_11899; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12929 = 3'h3 == state ? dirty_0_79 : _GEN_11900; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12930 = 3'h3 == state ? dirty_0_80 : _GEN_11901; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12931 = 3'h3 == state ? dirty_0_81 : _GEN_11902; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12932 = 3'h3 == state ? dirty_0_82 : _GEN_11903; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12933 = 3'h3 == state ? dirty_0_83 : _GEN_11904; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12934 = 3'h3 == state ? dirty_0_84 : _GEN_11905; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12935 = 3'h3 == state ? dirty_0_85 : _GEN_11906; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12936 = 3'h3 == state ? dirty_0_86 : _GEN_11907; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12937 = 3'h3 == state ? dirty_0_87 : _GEN_11908; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12938 = 3'h3 == state ? dirty_0_88 : _GEN_11909; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12939 = 3'h3 == state ? dirty_0_89 : _GEN_11910; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12940 = 3'h3 == state ? dirty_0_90 : _GEN_11911; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12941 = 3'h3 == state ? dirty_0_91 : _GEN_11912; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12942 = 3'h3 == state ? dirty_0_92 : _GEN_11913; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12943 = 3'h3 == state ? dirty_0_93 : _GEN_11914; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12944 = 3'h3 == state ? dirty_0_94 : _GEN_11915; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12945 = 3'h3 == state ? dirty_0_95 : _GEN_11916; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12946 = 3'h3 == state ? dirty_0_96 : _GEN_11917; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12947 = 3'h3 == state ? dirty_0_97 : _GEN_11918; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12948 = 3'h3 == state ? dirty_0_98 : _GEN_11919; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12949 = 3'h3 == state ? dirty_0_99 : _GEN_11920; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12950 = 3'h3 == state ? dirty_0_100 : _GEN_11921; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12951 = 3'h3 == state ? dirty_0_101 : _GEN_11922; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12952 = 3'h3 == state ? dirty_0_102 : _GEN_11923; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12953 = 3'h3 == state ? dirty_0_103 : _GEN_11924; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12954 = 3'h3 == state ? dirty_0_104 : _GEN_11925; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12955 = 3'h3 == state ? dirty_0_105 : _GEN_11926; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12956 = 3'h3 == state ? dirty_0_106 : _GEN_11927; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12957 = 3'h3 == state ? dirty_0_107 : _GEN_11928; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12958 = 3'h3 == state ? dirty_0_108 : _GEN_11929; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12959 = 3'h3 == state ? dirty_0_109 : _GEN_11930; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12960 = 3'h3 == state ? dirty_0_110 : _GEN_11931; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12961 = 3'h3 == state ? dirty_0_111 : _GEN_11932; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12962 = 3'h3 == state ? dirty_0_112 : _GEN_11933; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12963 = 3'h3 == state ? dirty_0_113 : _GEN_11934; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12964 = 3'h3 == state ? dirty_0_114 : _GEN_11935; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12965 = 3'h3 == state ? dirty_0_115 : _GEN_11936; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12966 = 3'h3 == state ? dirty_0_116 : _GEN_11937; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12967 = 3'h3 == state ? dirty_0_117 : _GEN_11938; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12968 = 3'h3 == state ? dirty_0_118 : _GEN_11939; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12969 = 3'h3 == state ? dirty_0_119 : _GEN_11940; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12970 = 3'h3 == state ? dirty_0_120 : _GEN_11941; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12971 = 3'h3 == state ? dirty_0_121 : _GEN_11942; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12972 = 3'h3 == state ? dirty_0_122 : _GEN_11943; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12973 = 3'h3 == state ? dirty_0_123 : _GEN_11944; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12974 = 3'h3 == state ? dirty_0_124 : _GEN_11945; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12975 = 3'h3 == state ? dirty_0_125 : _GEN_11946; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12976 = 3'h3 == state ? dirty_0_126 : _GEN_11947; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12977 = 3'h3 == state ? dirty_0_127 : _GEN_11948; // @[d_cache.scala 78:18 24:26]
  wire  _GEN_12978 = 3'h3 == state ? dirty_1_0 : _GEN_11949; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12979 = 3'h3 == state ? dirty_1_1 : _GEN_11950; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12980 = 3'h3 == state ? dirty_1_2 : _GEN_11951; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12981 = 3'h3 == state ? dirty_1_3 : _GEN_11952; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12982 = 3'h3 == state ? dirty_1_4 : _GEN_11953; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12983 = 3'h3 == state ? dirty_1_5 : _GEN_11954; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12984 = 3'h3 == state ? dirty_1_6 : _GEN_11955; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12985 = 3'h3 == state ? dirty_1_7 : _GEN_11956; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12986 = 3'h3 == state ? dirty_1_8 : _GEN_11957; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12987 = 3'h3 == state ? dirty_1_9 : _GEN_11958; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12988 = 3'h3 == state ? dirty_1_10 : _GEN_11959; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12989 = 3'h3 == state ? dirty_1_11 : _GEN_11960; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12990 = 3'h3 == state ? dirty_1_12 : _GEN_11961; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12991 = 3'h3 == state ? dirty_1_13 : _GEN_11962; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12992 = 3'h3 == state ? dirty_1_14 : _GEN_11963; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12993 = 3'h3 == state ? dirty_1_15 : _GEN_11964; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12994 = 3'h3 == state ? dirty_1_16 : _GEN_11965; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12995 = 3'h3 == state ? dirty_1_17 : _GEN_11966; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12996 = 3'h3 == state ? dirty_1_18 : _GEN_11967; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12997 = 3'h3 == state ? dirty_1_19 : _GEN_11968; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12998 = 3'h3 == state ? dirty_1_20 : _GEN_11969; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_12999 = 3'h3 == state ? dirty_1_21 : _GEN_11970; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13000 = 3'h3 == state ? dirty_1_22 : _GEN_11971; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13001 = 3'h3 == state ? dirty_1_23 : _GEN_11972; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13002 = 3'h3 == state ? dirty_1_24 : _GEN_11973; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13003 = 3'h3 == state ? dirty_1_25 : _GEN_11974; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13004 = 3'h3 == state ? dirty_1_26 : _GEN_11975; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13005 = 3'h3 == state ? dirty_1_27 : _GEN_11976; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13006 = 3'h3 == state ? dirty_1_28 : _GEN_11977; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13007 = 3'h3 == state ? dirty_1_29 : _GEN_11978; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13008 = 3'h3 == state ? dirty_1_30 : _GEN_11979; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13009 = 3'h3 == state ? dirty_1_31 : _GEN_11980; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13010 = 3'h3 == state ? dirty_1_32 : _GEN_11981; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13011 = 3'h3 == state ? dirty_1_33 : _GEN_11982; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13012 = 3'h3 == state ? dirty_1_34 : _GEN_11983; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13013 = 3'h3 == state ? dirty_1_35 : _GEN_11984; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13014 = 3'h3 == state ? dirty_1_36 : _GEN_11985; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13015 = 3'h3 == state ? dirty_1_37 : _GEN_11986; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13016 = 3'h3 == state ? dirty_1_38 : _GEN_11987; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13017 = 3'h3 == state ? dirty_1_39 : _GEN_11988; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13018 = 3'h3 == state ? dirty_1_40 : _GEN_11989; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13019 = 3'h3 == state ? dirty_1_41 : _GEN_11990; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13020 = 3'h3 == state ? dirty_1_42 : _GEN_11991; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13021 = 3'h3 == state ? dirty_1_43 : _GEN_11992; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13022 = 3'h3 == state ? dirty_1_44 : _GEN_11993; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13023 = 3'h3 == state ? dirty_1_45 : _GEN_11994; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13024 = 3'h3 == state ? dirty_1_46 : _GEN_11995; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13025 = 3'h3 == state ? dirty_1_47 : _GEN_11996; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13026 = 3'h3 == state ? dirty_1_48 : _GEN_11997; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13027 = 3'h3 == state ? dirty_1_49 : _GEN_11998; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13028 = 3'h3 == state ? dirty_1_50 : _GEN_11999; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13029 = 3'h3 == state ? dirty_1_51 : _GEN_12000; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13030 = 3'h3 == state ? dirty_1_52 : _GEN_12001; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13031 = 3'h3 == state ? dirty_1_53 : _GEN_12002; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13032 = 3'h3 == state ? dirty_1_54 : _GEN_12003; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13033 = 3'h3 == state ? dirty_1_55 : _GEN_12004; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13034 = 3'h3 == state ? dirty_1_56 : _GEN_12005; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13035 = 3'h3 == state ? dirty_1_57 : _GEN_12006; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13036 = 3'h3 == state ? dirty_1_58 : _GEN_12007; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13037 = 3'h3 == state ? dirty_1_59 : _GEN_12008; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13038 = 3'h3 == state ? dirty_1_60 : _GEN_12009; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13039 = 3'h3 == state ? dirty_1_61 : _GEN_12010; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13040 = 3'h3 == state ? dirty_1_62 : _GEN_12011; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13041 = 3'h3 == state ? dirty_1_63 : _GEN_12012; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13042 = 3'h3 == state ? dirty_1_64 : _GEN_12013; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13043 = 3'h3 == state ? dirty_1_65 : _GEN_12014; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13044 = 3'h3 == state ? dirty_1_66 : _GEN_12015; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13045 = 3'h3 == state ? dirty_1_67 : _GEN_12016; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13046 = 3'h3 == state ? dirty_1_68 : _GEN_12017; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13047 = 3'h3 == state ? dirty_1_69 : _GEN_12018; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13048 = 3'h3 == state ? dirty_1_70 : _GEN_12019; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13049 = 3'h3 == state ? dirty_1_71 : _GEN_12020; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13050 = 3'h3 == state ? dirty_1_72 : _GEN_12021; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13051 = 3'h3 == state ? dirty_1_73 : _GEN_12022; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13052 = 3'h3 == state ? dirty_1_74 : _GEN_12023; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13053 = 3'h3 == state ? dirty_1_75 : _GEN_12024; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13054 = 3'h3 == state ? dirty_1_76 : _GEN_12025; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13055 = 3'h3 == state ? dirty_1_77 : _GEN_12026; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13056 = 3'h3 == state ? dirty_1_78 : _GEN_12027; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13057 = 3'h3 == state ? dirty_1_79 : _GEN_12028; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13058 = 3'h3 == state ? dirty_1_80 : _GEN_12029; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13059 = 3'h3 == state ? dirty_1_81 : _GEN_12030; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13060 = 3'h3 == state ? dirty_1_82 : _GEN_12031; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13061 = 3'h3 == state ? dirty_1_83 : _GEN_12032; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13062 = 3'h3 == state ? dirty_1_84 : _GEN_12033; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13063 = 3'h3 == state ? dirty_1_85 : _GEN_12034; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13064 = 3'h3 == state ? dirty_1_86 : _GEN_12035; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13065 = 3'h3 == state ? dirty_1_87 : _GEN_12036; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13066 = 3'h3 == state ? dirty_1_88 : _GEN_12037; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13067 = 3'h3 == state ? dirty_1_89 : _GEN_12038; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13068 = 3'h3 == state ? dirty_1_90 : _GEN_12039; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13069 = 3'h3 == state ? dirty_1_91 : _GEN_12040; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13070 = 3'h3 == state ? dirty_1_92 : _GEN_12041; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13071 = 3'h3 == state ? dirty_1_93 : _GEN_12042; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13072 = 3'h3 == state ? dirty_1_94 : _GEN_12043; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13073 = 3'h3 == state ? dirty_1_95 : _GEN_12044; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13074 = 3'h3 == state ? dirty_1_96 : _GEN_12045; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13075 = 3'h3 == state ? dirty_1_97 : _GEN_12046; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13076 = 3'h3 == state ? dirty_1_98 : _GEN_12047; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13077 = 3'h3 == state ? dirty_1_99 : _GEN_12048; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13078 = 3'h3 == state ? dirty_1_100 : _GEN_12049; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13079 = 3'h3 == state ? dirty_1_101 : _GEN_12050; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13080 = 3'h3 == state ? dirty_1_102 : _GEN_12051; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13081 = 3'h3 == state ? dirty_1_103 : _GEN_12052; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13082 = 3'h3 == state ? dirty_1_104 : _GEN_12053; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13083 = 3'h3 == state ? dirty_1_105 : _GEN_12054; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13084 = 3'h3 == state ? dirty_1_106 : _GEN_12055; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13085 = 3'h3 == state ? dirty_1_107 : _GEN_12056; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13086 = 3'h3 == state ? dirty_1_108 : _GEN_12057; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13087 = 3'h3 == state ? dirty_1_109 : _GEN_12058; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13088 = 3'h3 == state ? dirty_1_110 : _GEN_12059; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13089 = 3'h3 == state ? dirty_1_111 : _GEN_12060; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13090 = 3'h3 == state ? dirty_1_112 : _GEN_12061; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13091 = 3'h3 == state ? dirty_1_113 : _GEN_12062; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13092 = 3'h3 == state ? dirty_1_114 : _GEN_12063; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13093 = 3'h3 == state ? dirty_1_115 : _GEN_12064; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13094 = 3'h3 == state ? dirty_1_116 : _GEN_12065; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13095 = 3'h3 == state ? dirty_1_117 : _GEN_12066; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13096 = 3'h3 == state ? dirty_1_118 : _GEN_12067; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13097 = 3'h3 == state ? dirty_1_119 : _GEN_12068; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13098 = 3'h3 == state ? dirty_1_120 : _GEN_12069; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13099 = 3'h3 == state ? dirty_1_121 : _GEN_12070; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13100 = 3'h3 == state ? dirty_1_122 : _GEN_12071; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13101 = 3'h3 == state ? dirty_1_123 : _GEN_12072; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13102 = 3'h3 == state ? dirty_1_124 : _GEN_12073; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13103 = 3'h3 == state ? dirty_1_125 : _GEN_12074; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13104 = 3'h3 == state ? dirty_1_126 : _GEN_12075; // @[d_cache.scala 78:18 25:26]
  wire  _GEN_13105 = 3'h3 == state ? dirty_1_127 : _GEN_12076; // @[d_cache.scala 78:18 25:26]
  wire [41:0] _GEN_14134 = 3'h2 == state ? {{10'd0}, write_back_addr} : _GEN_12849; // @[d_cache.scala 78:18 30:34]
  wire [41:0] _GEN_15163 = 3'h1 == state ? {{10'd0}, write_back_addr} : _GEN_14134; // @[d_cache.scala 78:18 30:34]
  wire [41:0] _GEN_16192 = 3'h0 == state ? {{10'd0}, write_back_addr} : _GEN_15163; // @[d_cache.scala 78:18 30:34]
  wire [63:0] _io_to_lsu_rdata_T_1 = _GEN_1160 >> offset; // @[d_cache.scala 221:49]
  wire [63:0] _io_to_lsu_rdata_T_3 = _GEN_5393 >> offset; // @[d_cache.scala 228:49]
  wire [63:0] _GEN_16449 = way1_hit ? _io_to_lsu_rdata_T_3 : 64'h0; // @[d_cache.scala 227:33 228:33 235:33]
  wire [63:0] _GEN_16453 = way0_hit ? _io_to_lsu_rdata_T_1 : _GEN_16449; // @[d_cache.scala 220:23 221:33]
  wire  _GEN_16455 = way0_hit | way1_hit; // @[d_cache.scala 220:23 223:34]
  wire  _GEN_16457 = way1_hit ? 1'h0 : 1'h1; // @[d_cache.scala 259:33 261:35 268:35]
  wire  _GEN_16458 = way0_hit ? 1'h0 : _GEN_16457; // @[d_cache.scala 252:23 254:35]
  wire  _T_72 = state == 3'h3; // @[d_cache.scala 274:21]
  wire  _T_75 = state == 3'h6; // @[d_cache.scala 323:21]
  wire [31:0] _GEN_16461 = state == 3'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 323:35 331:26 347:26]
  wire  _GEN_16462 = state == 3'h6 ? 1'h0 : io_from_lsu_rready; // @[d_cache.scala 323:35 332:26 348:26]
  wire [31:0] _GEN_16463 = state == 3'h6 ? write_back_addr : 32'h0; // @[d_cache.scala 323:35 333:26 349:26]
  wire [63:0] _GEN_16464 = state == 3'h6 ? write_back_data : 64'h0; // @[d_cache.scala 323:35 335:25 351:25]
  wire [31:0] _GEN_16465 = state == 3'h6 ? 32'hffffffff : 32'h0; // @[d_cache.scala 323:35 336:25 352:25]
  wire  _GEN_16467 = state == 3'h5 | _T_75; // @[d_cache.scala 307:31 309:27]
  wire [31:0] _GEN_16468 = state == 3'h5 ? io_from_lsu_araddr : _GEN_16461; // @[d_cache.scala 307:31 315:26]
  wire  _GEN_16469 = state == 3'h5 ? io_from_lsu_rready : _GEN_16462; // @[d_cache.scala 307:31 316:26]
  wire [31:0] _GEN_16470 = state == 3'h5 ? 32'h0 : _GEN_16463; // @[d_cache.scala 307:31 317:26]
  wire  _GEN_16471 = state == 3'h5 ? 1'h0 : _T_75; // @[d_cache.scala 307:31 318:27]
  wire [63:0] _GEN_16472 = state == 3'h5 ? 64'h0 : _GEN_16464; // @[d_cache.scala 307:31 319:25]
  wire [31:0] _GEN_16473 = state == 3'h5 ? 32'h0 : _GEN_16465; // @[d_cache.scala 307:31 320:25]
  wire  _GEN_16475 = state == 3'h4 | _GEN_16467; // @[d_cache.scala 290:31 292:27]
  wire  _GEN_16476 = state == 3'h4 & io_from_axi_wready; // @[d_cache.scala 290:31 294:26]
  wire  _GEN_16477 = state == 3'h4 & io_from_axi_bvalid; // @[d_cache.scala 290:31 295:26]
  wire  _GEN_16478 = state == 3'h4 & io_from_axi_awready; // @[d_cache.scala 290:31 296:27]
  wire [31:0] _GEN_16479 = state == 3'h4 ? 32'h0 : _GEN_16468; // @[d_cache.scala 290:31 298:26]
  wire  _GEN_16480 = state == 3'h4 ? io_from_lsu_rready : _GEN_16469; // @[d_cache.scala 290:31 299:26]
  wire [31:0] _GEN_16481 = state == 3'h4 ? io_from_lsu_awaddr : _GEN_16470; // @[d_cache.scala 290:31 300:26]
  wire  _GEN_16482 = state == 3'h4 ? io_from_lsu_awvalid : _GEN_16471; // @[d_cache.scala 290:31 301:27]
  wire [63:0] _GEN_16483 = state == 3'h4 ? {{32'd0}, io_from_lsu_wdata} : _GEN_16472; // @[d_cache.scala 290:31 302:25]
  wire [31:0] _GEN_16484 = state == 3'h4 ? {{24'd0}, io_from_lsu_wstrb} : _GEN_16473; // @[d_cache.scala 290:31 303:25]
  wire  _GEN_16485 = state == 3'h4 ? io_from_lsu_wvalid : _GEN_16471; // @[d_cache.scala 290:31 304:26]
  wire  _GEN_16486 = state == 3'h4 ? io_from_lsu_bready : _GEN_16471; // @[d_cache.scala 290:31 305:26]
  wire  _GEN_16488 = state == 3'h3 | _GEN_16475; // @[d_cache.scala 274:31 276:27]
  wire  _GEN_16489 = state == 3'h3 ? 1'h0 : _GEN_16476; // @[d_cache.scala 274:31 278:26]
  wire  _GEN_16490 = state == 3'h3 ? 1'h0 : _GEN_16477; // @[d_cache.scala 274:31 279:26]
  wire  _GEN_16491 = state == 3'h3 ? 1'h0 : _GEN_16478; // @[d_cache.scala 274:31 280:27]
  wire [31:0] _GEN_16493 = state == 3'h3 ? io_from_lsu_araddr : _GEN_16479; // @[d_cache.scala 274:31 282:26]
  wire  _GEN_16494 = state == 3'h3 ? io_from_lsu_rready : _GEN_16480; // @[d_cache.scala 274:31 283:26]
  wire [31:0] _GEN_16495 = state == 3'h3 ? 32'h0 : _GEN_16481; // @[d_cache.scala 274:31 284:26]
  wire  _GEN_16496 = state == 3'h3 ? 1'h0 : _GEN_16482; // @[d_cache.scala 274:31 285:27]
  wire [63:0] _GEN_16497 = state == 3'h3 ? 64'h0 : _GEN_16483; // @[d_cache.scala 274:31 286:25]
  wire [31:0] _GEN_16498 = state == 3'h3 ? 32'h0 : _GEN_16484; // @[d_cache.scala 274:31 287:25]
  wire  _GEN_16499 = state == 3'h3 ? 1'h0 : _GEN_16485; // @[d_cache.scala 274:31 288:26]
  wire  _GEN_16500 = state == 3'h3 ? 1'h0 : _GEN_16486; // @[d_cache.scala 274:31 289:26]
  wire  _GEN_16501 = state == 3'h2 ? 1'h0 : _T_72; // @[d_cache.scala 242:33 243:27]
  wire [31:0] _GEN_16502 = state == 3'h2 ? io_from_lsu_araddr : _GEN_16493; // @[d_cache.scala 242:33 244:26]
  wire  _GEN_16503 = state == 3'h2 ? 1'h0 : _GEN_16494; // @[d_cache.scala 242:33 245:26]
  wire [31:0] _GEN_16504 = state == 3'h2 ? 32'h0 : _GEN_16495; // @[d_cache.scala 242:33 246:26]
  wire  _GEN_16505 = state == 3'h2 ? 1'h0 : _GEN_16496; // @[d_cache.scala 242:33 247:27]
  wire [63:0] _GEN_16506 = state == 3'h2 ? 64'h0 : _GEN_16497; // @[d_cache.scala 242:33 248:25]
  wire [31:0] _GEN_16507 = state == 3'h2 ? 32'h0 : _GEN_16498; // @[d_cache.scala 242:33 249:25]
  wire  _GEN_16508 = state == 3'h2 ? 1'h0 : _GEN_16499; // @[d_cache.scala 242:33 250:26]
  wire  _GEN_16509 = state == 3'h2 ? 1'h0 : _GEN_16500; // @[d_cache.scala 242:33 251:26]
  wire  _GEN_16511 = state == 3'h2 ? _GEN_16458 : _GEN_16488; // @[d_cache.scala 242:33]
  wire  _GEN_16512 = state == 3'h2 ? _GEN_16455 : _GEN_16489; // @[d_cache.scala 242:33]
  wire  _GEN_16513 = state == 3'h2 ? _GEN_16455 : _GEN_16491; // @[d_cache.scala 242:33]
  wire  _GEN_16514 = state == 3'h2 ? _GEN_16455 : _GEN_16490; // @[d_cache.scala 242:33]
  wire  _GEN_16515 = state == 3'h1 ? 1'h0 : _GEN_16501; // @[d_cache.scala 210:33 211:27]
  wire [31:0] _GEN_16516 = state == 3'h1 ? io_from_lsu_araddr : _GEN_16502; // @[d_cache.scala 210:33 212:26]
  wire  _GEN_16517 = state == 3'h1 ? io_from_lsu_rready : _GEN_16503; // @[d_cache.scala 210:33 213:26]
  wire [31:0] _GEN_16518 = state == 3'h1 ? 32'h0 : _GEN_16504; // @[d_cache.scala 210:33 214:26]
  wire  _GEN_16519 = state == 3'h1 ? 1'h0 : _GEN_16505; // @[d_cache.scala 210:33 215:27]
  wire [63:0] _GEN_16520 = state == 3'h1 ? 64'h0 : _GEN_16506; // @[d_cache.scala 210:33 216:25]
  wire [31:0] _GEN_16521 = state == 3'h1 ? 32'h0 : _GEN_16507; // @[d_cache.scala 210:33 217:25]
  wire  _GEN_16522 = state == 3'h1 ? 1'h0 : _GEN_16508; // @[d_cache.scala 210:33 218:26]
  wire  _GEN_16523 = state == 3'h1 ? io_from_lsu_bready : _GEN_16509; // @[d_cache.scala 210:33 219:26]
  wire [63:0] _GEN_16524 = state == 3'h1 ? _GEN_16453 : 64'h0; // @[d_cache.scala 210:33]
  wire  _GEN_16525 = state == 3'h1 | _GEN_16511; // @[d_cache.scala 210:33]
  wire  _GEN_16526 = state == 3'h1 & _GEN_16455; // @[d_cache.scala 210:33]
  wire  _GEN_16527 = state == 3'h1 ? 1'h0 : _GEN_16512; // @[d_cache.scala 210:33]
  wire  _GEN_16528 = state == 3'h1 ? 1'h0 : _GEN_16513; // @[d_cache.scala 210:33]
  wire  _GEN_16529 = state == 3'h1 ? 1'h0 : _GEN_16514; // @[d_cache.scala 210:33]
  wire [63:0] _GEN_16541 = state == 3'h0 ? 64'h0 : _GEN_16520; // @[d_cache.scala 194:23 206:25]
  wire [31:0] _GEN_16542 = state == 3'h0 ? 32'h0 : _GEN_16521; // @[d_cache.scala 194:23 207:25]
  wire [41:0] _GEN_17833 = reset ? 42'h0 : _GEN_16192; // @[d_cache.scala 30:{34,34}]
  wire  _GEN_17835 = ~_T_24 & _T_25; // @[d_cache.scala 90:27]
  assign io_to_lsu_arready = state == 3'h0 ? io_from_axi_arready : _GEN_16525; // @[d_cache.scala 194:23 196:27]
  assign io_to_lsu_rdata = state == 3'h0 ? 64'h0 : _GEN_16524; // @[d_cache.scala 194:23 195:25]
  assign io_to_lsu_rvalid = state == 3'h0 ? 1'h0 : _GEN_16526; // @[d_cache.scala 194:23 197:26]
  assign io_to_lsu_awready = state == 3'h0 ? io_from_axi_awready : _GEN_16528; // @[d_cache.scala 194:23 200:27]
  assign io_to_lsu_wready = state == 3'h0 ? 1'h0 : _GEN_16527; // @[d_cache.scala 194:23 198:26]
  assign io_to_lsu_bvalid = state == 3'h0 ? 1'h0 : _GEN_16529; // @[d_cache.scala 194:23 199:26]
  assign io_to_axi_araddr = state == 3'h0 ? io_from_lsu_araddr : _GEN_16516; // @[d_cache.scala 194:23 202:26]
  assign io_to_axi_arvalid = state == 3'h0 ? 1'h0 : _GEN_16515; // @[d_cache.scala 194:23 201:27]
  assign io_to_axi_rready = state == 3'h0 ? io_from_lsu_rready : _GEN_16517; // @[d_cache.scala 194:23 203:26]
  assign io_to_axi_awaddr = state == 3'h0 ? 32'h0 : _GEN_16518; // @[d_cache.scala 194:23 204:26]
  assign io_to_axi_awvalid = state == 3'h0 ? 1'h0 : _GEN_16519; // @[d_cache.scala 194:23 205:27]
  assign io_to_axi_wdata = _GEN_16541[31:0];
  assign io_to_axi_wstrb = _GEN_16542[7:0];
  assign io_to_axi_wvalid = state == 3'h0 ? 1'h0 : _GEN_16522; // @[d_cache.scala 194:23 208:26]
  assign io_to_axi_bready = state == 3'h0 ? io_from_lsu_bready : _GEN_16523; // @[d_cache.scala 194:23 209:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_0 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_0 <= _GEN_2059;
        end else begin
          ram_0_0 <= _GEN_12079;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_1 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_1 <= _GEN_2060;
        end else begin
          ram_0_1 <= _GEN_12080;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_2 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_2 <= _GEN_2061;
        end else begin
          ram_0_2 <= _GEN_12081;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_3 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_3 <= _GEN_2062;
        end else begin
          ram_0_3 <= _GEN_12082;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_4 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_4 <= _GEN_2063;
        end else begin
          ram_0_4 <= _GEN_12083;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_5 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_5 <= _GEN_2064;
        end else begin
          ram_0_5 <= _GEN_12084;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_6 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_6 <= _GEN_2065;
        end else begin
          ram_0_6 <= _GEN_12085;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_7 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_7 <= _GEN_2066;
        end else begin
          ram_0_7 <= _GEN_12086;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_8 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_8 <= _GEN_2067;
        end else begin
          ram_0_8 <= _GEN_12087;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_9 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_9 <= _GEN_2068;
        end else begin
          ram_0_9 <= _GEN_12088;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_10 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_10 <= _GEN_2069;
        end else begin
          ram_0_10 <= _GEN_12089;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_11 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_11 <= _GEN_2070;
        end else begin
          ram_0_11 <= _GEN_12090;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_12 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_12 <= _GEN_2071;
        end else begin
          ram_0_12 <= _GEN_12091;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_13 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_13 <= _GEN_2072;
        end else begin
          ram_0_13 <= _GEN_12092;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_14 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_14 <= _GEN_2073;
        end else begin
          ram_0_14 <= _GEN_12093;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_15 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_15 <= _GEN_2074;
        end else begin
          ram_0_15 <= _GEN_12094;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_16 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_16 <= _GEN_2075;
        end else begin
          ram_0_16 <= _GEN_12095;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_17 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_17 <= _GEN_2076;
        end else begin
          ram_0_17 <= _GEN_12096;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_18 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_18 <= _GEN_2077;
        end else begin
          ram_0_18 <= _GEN_12097;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_19 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_19 <= _GEN_2078;
        end else begin
          ram_0_19 <= _GEN_12098;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_20 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_20 <= _GEN_2079;
        end else begin
          ram_0_20 <= _GEN_12099;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_21 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_21 <= _GEN_2080;
        end else begin
          ram_0_21 <= _GEN_12100;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_22 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_22 <= _GEN_2081;
        end else begin
          ram_0_22 <= _GEN_12101;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_23 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_23 <= _GEN_2082;
        end else begin
          ram_0_23 <= _GEN_12102;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_24 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_24 <= _GEN_2083;
        end else begin
          ram_0_24 <= _GEN_12103;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_25 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_25 <= _GEN_2084;
        end else begin
          ram_0_25 <= _GEN_12104;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_26 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_26 <= _GEN_2085;
        end else begin
          ram_0_26 <= _GEN_12105;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_27 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_27 <= _GEN_2086;
        end else begin
          ram_0_27 <= _GEN_12106;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_28 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_28 <= _GEN_2087;
        end else begin
          ram_0_28 <= _GEN_12107;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_29 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_29 <= _GEN_2088;
        end else begin
          ram_0_29 <= _GEN_12108;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_30 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_30 <= _GEN_2089;
        end else begin
          ram_0_30 <= _GEN_12109;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_31 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_31 <= _GEN_2090;
        end else begin
          ram_0_31 <= _GEN_12110;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_32 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_32 <= _GEN_2091;
        end else begin
          ram_0_32 <= _GEN_12111;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_33 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_33 <= _GEN_2092;
        end else begin
          ram_0_33 <= _GEN_12112;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_34 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_34 <= _GEN_2093;
        end else begin
          ram_0_34 <= _GEN_12113;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_35 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_35 <= _GEN_2094;
        end else begin
          ram_0_35 <= _GEN_12114;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_36 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_36 <= _GEN_2095;
        end else begin
          ram_0_36 <= _GEN_12115;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_37 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_37 <= _GEN_2096;
        end else begin
          ram_0_37 <= _GEN_12116;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_38 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_38 <= _GEN_2097;
        end else begin
          ram_0_38 <= _GEN_12117;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_39 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_39 <= _GEN_2098;
        end else begin
          ram_0_39 <= _GEN_12118;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_40 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_40 <= _GEN_2099;
        end else begin
          ram_0_40 <= _GEN_12119;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_41 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_41 <= _GEN_2100;
        end else begin
          ram_0_41 <= _GEN_12120;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_42 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_42 <= _GEN_2101;
        end else begin
          ram_0_42 <= _GEN_12121;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_43 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_43 <= _GEN_2102;
        end else begin
          ram_0_43 <= _GEN_12122;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_44 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_44 <= _GEN_2103;
        end else begin
          ram_0_44 <= _GEN_12123;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_45 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_45 <= _GEN_2104;
        end else begin
          ram_0_45 <= _GEN_12124;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_46 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_46 <= _GEN_2105;
        end else begin
          ram_0_46 <= _GEN_12125;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_47 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_47 <= _GEN_2106;
        end else begin
          ram_0_47 <= _GEN_12126;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_48 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_48 <= _GEN_2107;
        end else begin
          ram_0_48 <= _GEN_12127;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_49 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_49 <= _GEN_2108;
        end else begin
          ram_0_49 <= _GEN_12128;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_50 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_50 <= _GEN_2109;
        end else begin
          ram_0_50 <= _GEN_12129;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_51 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_51 <= _GEN_2110;
        end else begin
          ram_0_51 <= _GEN_12130;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_52 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_52 <= _GEN_2111;
        end else begin
          ram_0_52 <= _GEN_12131;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_53 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_53 <= _GEN_2112;
        end else begin
          ram_0_53 <= _GEN_12132;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_54 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_54 <= _GEN_2113;
        end else begin
          ram_0_54 <= _GEN_12133;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_55 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_55 <= _GEN_2114;
        end else begin
          ram_0_55 <= _GEN_12134;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_56 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_56 <= _GEN_2115;
        end else begin
          ram_0_56 <= _GEN_12135;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_57 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_57 <= _GEN_2116;
        end else begin
          ram_0_57 <= _GEN_12136;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_58 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_58 <= _GEN_2117;
        end else begin
          ram_0_58 <= _GEN_12137;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_59 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_59 <= _GEN_2118;
        end else begin
          ram_0_59 <= _GEN_12138;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_60 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_60 <= _GEN_2119;
        end else begin
          ram_0_60 <= _GEN_12139;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_61 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_61 <= _GEN_2120;
        end else begin
          ram_0_61 <= _GEN_12140;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_62 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_62 <= _GEN_2121;
        end else begin
          ram_0_62 <= _GEN_12141;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_63 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_63 <= _GEN_2122;
        end else begin
          ram_0_63 <= _GEN_12142;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_64 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_64 <= _GEN_2123;
        end else begin
          ram_0_64 <= _GEN_12143;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_65 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_65 <= _GEN_2124;
        end else begin
          ram_0_65 <= _GEN_12144;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_66 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_66 <= _GEN_2125;
        end else begin
          ram_0_66 <= _GEN_12145;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_67 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_67 <= _GEN_2126;
        end else begin
          ram_0_67 <= _GEN_12146;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_68 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_68 <= _GEN_2127;
        end else begin
          ram_0_68 <= _GEN_12147;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_69 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_69 <= _GEN_2128;
        end else begin
          ram_0_69 <= _GEN_12148;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_70 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_70 <= _GEN_2129;
        end else begin
          ram_0_70 <= _GEN_12149;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_71 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_71 <= _GEN_2130;
        end else begin
          ram_0_71 <= _GEN_12150;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_72 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_72 <= _GEN_2131;
        end else begin
          ram_0_72 <= _GEN_12151;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_73 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_73 <= _GEN_2132;
        end else begin
          ram_0_73 <= _GEN_12152;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_74 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_74 <= _GEN_2133;
        end else begin
          ram_0_74 <= _GEN_12153;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_75 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_75 <= _GEN_2134;
        end else begin
          ram_0_75 <= _GEN_12154;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_76 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_76 <= _GEN_2135;
        end else begin
          ram_0_76 <= _GEN_12155;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_77 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_77 <= _GEN_2136;
        end else begin
          ram_0_77 <= _GEN_12156;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_78 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_78 <= _GEN_2137;
        end else begin
          ram_0_78 <= _GEN_12157;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_79 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_79 <= _GEN_2138;
        end else begin
          ram_0_79 <= _GEN_12158;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_80 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_80 <= _GEN_2139;
        end else begin
          ram_0_80 <= _GEN_12159;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_81 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_81 <= _GEN_2140;
        end else begin
          ram_0_81 <= _GEN_12160;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_82 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_82 <= _GEN_2141;
        end else begin
          ram_0_82 <= _GEN_12161;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_83 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_83 <= _GEN_2142;
        end else begin
          ram_0_83 <= _GEN_12162;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_84 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_84 <= _GEN_2143;
        end else begin
          ram_0_84 <= _GEN_12163;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_85 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_85 <= _GEN_2144;
        end else begin
          ram_0_85 <= _GEN_12164;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_86 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_86 <= _GEN_2145;
        end else begin
          ram_0_86 <= _GEN_12165;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_87 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_87 <= _GEN_2146;
        end else begin
          ram_0_87 <= _GEN_12166;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_88 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_88 <= _GEN_2147;
        end else begin
          ram_0_88 <= _GEN_12167;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_89 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_89 <= _GEN_2148;
        end else begin
          ram_0_89 <= _GEN_12168;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_90 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_90 <= _GEN_2149;
        end else begin
          ram_0_90 <= _GEN_12169;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_91 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_91 <= _GEN_2150;
        end else begin
          ram_0_91 <= _GEN_12170;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_92 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_92 <= _GEN_2151;
        end else begin
          ram_0_92 <= _GEN_12171;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_93 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_93 <= _GEN_2152;
        end else begin
          ram_0_93 <= _GEN_12172;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_94 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_94 <= _GEN_2153;
        end else begin
          ram_0_94 <= _GEN_12173;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_95 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_95 <= _GEN_2154;
        end else begin
          ram_0_95 <= _GEN_12174;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_96 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_96 <= _GEN_2155;
        end else begin
          ram_0_96 <= _GEN_12175;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_97 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_97 <= _GEN_2156;
        end else begin
          ram_0_97 <= _GEN_12176;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_98 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_98 <= _GEN_2157;
        end else begin
          ram_0_98 <= _GEN_12177;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_99 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_99 <= _GEN_2158;
        end else begin
          ram_0_99 <= _GEN_12178;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_100 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_100 <= _GEN_2159;
        end else begin
          ram_0_100 <= _GEN_12179;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_101 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_101 <= _GEN_2160;
        end else begin
          ram_0_101 <= _GEN_12180;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_102 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_102 <= _GEN_2161;
        end else begin
          ram_0_102 <= _GEN_12181;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_103 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_103 <= _GEN_2162;
        end else begin
          ram_0_103 <= _GEN_12182;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_104 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_104 <= _GEN_2163;
        end else begin
          ram_0_104 <= _GEN_12183;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_105 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_105 <= _GEN_2164;
        end else begin
          ram_0_105 <= _GEN_12184;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_106 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_106 <= _GEN_2165;
        end else begin
          ram_0_106 <= _GEN_12185;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_107 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_107 <= _GEN_2166;
        end else begin
          ram_0_107 <= _GEN_12186;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_108 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_108 <= _GEN_2167;
        end else begin
          ram_0_108 <= _GEN_12187;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_109 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_109 <= _GEN_2168;
        end else begin
          ram_0_109 <= _GEN_12188;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_110 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_110 <= _GEN_2169;
        end else begin
          ram_0_110 <= _GEN_12189;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_111 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_111 <= _GEN_2170;
        end else begin
          ram_0_111 <= _GEN_12190;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_112 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_112 <= _GEN_2171;
        end else begin
          ram_0_112 <= _GEN_12191;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_113 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_113 <= _GEN_2172;
        end else begin
          ram_0_113 <= _GEN_12192;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_114 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_114 <= _GEN_2173;
        end else begin
          ram_0_114 <= _GEN_12193;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_115 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_115 <= _GEN_2174;
        end else begin
          ram_0_115 <= _GEN_12194;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_116 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_116 <= _GEN_2175;
        end else begin
          ram_0_116 <= _GEN_12195;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_117 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_117 <= _GEN_2176;
        end else begin
          ram_0_117 <= _GEN_12196;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_118 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_118 <= _GEN_2177;
        end else begin
          ram_0_118 <= _GEN_12197;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_119 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_119 <= _GEN_2178;
        end else begin
          ram_0_119 <= _GEN_12198;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_120 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_120 <= _GEN_2179;
        end else begin
          ram_0_120 <= _GEN_12199;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_121 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_121 <= _GEN_2180;
        end else begin
          ram_0_121 <= _GEN_12200;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_122 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_122 <= _GEN_2181;
        end else begin
          ram_0_122 <= _GEN_12201;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_123 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_123 <= _GEN_2182;
        end else begin
          ram_0_123 <= _GEN_12202;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_124 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_124 <= _GEN_2183;
        end else begin
          ram_0_124 <= _GEN_12203;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_125 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_125 <= _GEN_2184;
        end else begin
          ram_0_125 <= _GEN_12204;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_126 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_126 <= _GEN_2185;
        end else begin
          ram_0_126 <= _GEN_12205;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 18:24]
      ram_0_127 <= 64'h0; // @[d_cache.scala 18:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_0_127 <= _GEN_2186;
        end else begin
          ram_0_127 <= _GEN_12206;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_0 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_0 <= _GEN_2315;
        end else begin
          ram_1_0 <= _GEN_12464;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_1 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_1 <= _GEN_2316;
        end else begin
          ram_1_1 <= _GEN_12465;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_2 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_2 <= _GEN_2317;
        end else begin
          ram_1_2 <= _GEN_12466;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_3 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_3 <= _GEN_2318;
        end else begin
          ram_1_3 <= _GEN_12467;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_4 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_4 <= _GEN_2319;
        end else begin
          ram_1_4 <= _GEN_12468;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_5 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_5 <= _GEN_2320;
        end else begin
          ram_1_5 <= _GEN_12469;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_6 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_6 <= _GEN_2321;
        end else begin
          ram_1_6 <= _GEN_12470;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_7 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_7 <= _GEN_2322;
        end else begin
          ram_1_7 <= _GEN_12471;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_8 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_8 <= _GEN_2323;
        end else begin
          ram_1_8 <= _GEN_12472;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_9 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_9 <= _GEN_2324;
        end else begin
          ram_1_9 <= _GEN_12473;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_10 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_10 <= _GEN_2325;
        end else begin
          ram_1_10 <= _GEN_12474;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_11 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_11 <= _GEN_2326;
        end else begin
          ram_1_11 <= _GEN_12475;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_12 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_12 <= _GEN_2327;
        end else begin
          ram_1_12 <= _GEN_12476;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_13 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_13 <= _GEN_2328;
        end else begin
          ram_1_13 <= _GEN_12477;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_14 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_14 <= _GEN_2329;
        end else begin
          ram_1_14 <= _GEN_12478;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_15 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_15 <= _GEN_2330;
        end else begin
          ram_1_15 <= _GEN_12479;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_16 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_16 <= _GEN_2331;
        end else begin
          ram_1_16 <= _GEN_12480;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_17 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_17 <= _GEN_2332;
        end else begin
          ram_1_17 <= _GEN_12481;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_18 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_18 <= _GEN_2333;
        end else begin
          ram_1_18 <= _GEN_12482;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_19 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_19 <= _GEN_2334;
        end else begin
          ram_1_19 <= _GEN_12483;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_20 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_20 <= _GEN_2335;
        end else begin
          ram_1_20 <= _GEN_12484;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_21 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_21 <= _GEN_2336;
        end else begin
          ram_1_21 <= _GEN_12485;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_22 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_22 <= _GEN_2337;
        end else begin
          ram_1_22 <= _GEN_12486;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_23 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_23 <= _GEN_2338;
        end else begin
          ram_1_23 <= _GEN_12487;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_24 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_24 <= _GEN_2339;
        end else begin
          ram_1_24 <= _GEN_12488;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_25 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_25 <= _GEN_2340;
        end else begin
          ram_1_25 <= _GEN_12489;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_26 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_26 <= _GEN_2341;
        end else begin
          ram_1_26 <= _GEN_12490;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_27 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_27 <= _GEN_2342;
        end else begin
          ram_1_27 <= _GEN_12491;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_28 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_28 <= _GEN_2343;
        end else begin
          ram_1_28 <= _GEN_12492;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_29 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_29 <= _GEN_2344;
        end else begin
          ram_1_29 <= _GEN_12493;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_30 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_30 <= _GEN_2345;
        end else begin
          ram_1_30 <= _GEN_12494;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_31 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_31 <= _GEN_2346;
        end else begin
          ram_1_31 <= _GEN_12495;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_32 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_32 <= _GEN_2347;
        end else begin
          ram_1_32 <= _GEN_12496;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_33 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_33 <= _GEN_2348;
        end else begin
          ram_1_33 <= _GEN_12497;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_34 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_34 <= _GEN_2349;
        end else begin
          ram_1_34 <= _GEN_12498;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_35 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_35 <= _GEN_2350;
        end else begin
          ram_1_35 <= _GEN_12499;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_36 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_36 <= _GEN_2351;
        end else begin
          ram_1_36 <= _GEN_12500;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_37 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_37 <= _GEN_2352;
        end else begin
          ram_1_37 <= _GEN_12501;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_38 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_38 <= _GEN_2353;
        end else begin
          ram_1_38 <= _GEN_12502;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_39 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_39 <= _GEN_2354;
        end else begin
          ram_1_39 <= _GEN_12503;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_40 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_40 <= _GEN_2355;
        end else begin
          ram_1_40 <= _GEN_12504;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_41 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_41 <= _GEN_2356;
        end else begin
          ram_1_41 <= _GEN_12505;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_42 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_42 <= _GEN_2357;
        end else begin
          ram_1_42 <= _GEN_12506;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_43 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_43 <= _GEN_2358;
        end else begin
          ram_1_43 <= _GEN_12507;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_44 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_44 <= _GEN_2359;
        end else begin
          ram_1_44 <= _GEN_12508;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_45 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_45 <= _GEN_2360;
        end else begin
          ram_1_45 <= _GEN_12509;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_46 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_46 <= _GEN_2361;
        end else begin
          ram_1_46 <= _GEN_12510;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_47 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_47 <= _GEN_2362;
        end else begin
          ram_1_47 <= _GEN_12511;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_48 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_48 <= _GEN_2363;
        end else begin
          ram_1_48 <= _GEN_12512;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_49 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_49 <= _GEN_2364;
        end else begin
          ram_1_49 <= _GEN_12513;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_50 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_50 <= _GEN_2365;
        end else begin
          ram_1_50 <= _GEN_12514;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_51 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_51 <= _GEN_2366;
        end else begin
          ram_1_51 <= _GEN_12515;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_52 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_52 <= _GEN_2367;
        end else begin
          ram_1_52 <= _GEN_12516;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_53 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_53 <= _GEN_2368;
        end else begin
          ram_1_53 <= _GEN_12517;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_54 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_54 <= _GEN_2369;
        end else begin
          ram_1_54 <= _GEN_12518;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_55 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_55 <= _GEN_2370;
        end else begin
          ram_1_55 <= _GEN_12519;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_56 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_56 <= _GEN_2371;
        end else begin
          ram_1_56 <= _GEN_12520;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_57 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_57 <= _GEN_2372;
        end else begin
          ram_1_57 <= _GEN_12521;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_58 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_58 <= _GEN_2373;
        end else begin
          ram_1_58 <= _GEN_12522;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_59 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_59 <= _GEN_2374;
        end else begin
          ram_1_59 <= _GEN_12523;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_60 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_60 <= _GEN_2375;
        end else begin
          ram_1_60 <= _GEN_12524;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_61 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_61 <= _GEN_2376;
        end else begin
          ram_1_61 <= _GEN_12525;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_62 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_62 <= _GEN_2377;
        end else begin
          ram_1_62 <= _GEN_12526;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_63 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_63 <= _GEN_2378;
        end else begin
          ram_1_63 <= _GEN_12527;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_64 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_64 <= _GEN_2379;
        end else begin
          ram_1_64 <= _GEN_12528;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_65 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_65 <= _GEN_2380;
        end else begin
          ram_1_65 <= _GEN_12529;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_66 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_66 <= _GEN_2381;
        end else begin
          ram_1_66 <= _GEN_12530;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_67 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_67 <= _GEN_2382;
        end else begin
          ram_1_67 <= _GEN_12531;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_68 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_68 <= _GEN_2383;
        end else begin
          ram_1_68 <= _GEN_12532;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_69 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_69 <= _GEN_2384;
        end else begin
          ram_1_69 <= _GEN_12533;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_70 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_70 <= _GEN_2385;
        end else begin
          ram_1_70 <= _GEN_12534;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_71 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_71 <= _GEN_2386;
        end else begin
          ram_1_71 <= _GEN_12535;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_72 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_72 <= _GEN_2387;
        end else begin
          ram_1_72 <= _GEN_12536;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_73 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_73 <= _GEN_2388;
        end else begin
          ram_1_73 <= _GEN_12537;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_74 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_74 <= _GEN_2389;
        end else begin
          ram_1_74 <= _GEN_12538;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_75 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_75 <= _GEN_2390;
        end else begin
          ram_1_75 <= _GEN_12539;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_76 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_76 <= _GEN_2391;
        end else begin
          ram_1_76 <= _GEN_12540;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_77 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_77 <= _GEN_2392;
        end else begin
          ram_1_77 <= _GEN_12541;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_78 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_78 <= _GEN_2393;
        end else begin
          ram_1_78 <= _GEN_12542;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_79 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_79 <= _GEN_2394;
        end else begin
          ram_1_79 <= _GEN_12543;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_80 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_80 <= _GEN_2395;
        end else begin
          ram_1_80 <= _GEN_12544;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_81 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_81 <= _GEN_2396;
        end else begin
          ram_1_81 <= _GEN_12545;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_82 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_82 <= _GEN_2397;
        end else begin
          ram_1_82 <= _GEN_12546;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_83 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_83 <= _GEN_2398;
        end else begin
          ram_1_83 <= _GEN_12547;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_84 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_84 <= _GEN_2399;
        end else begin
          ram_1_84 <= _GEN_12548;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_85 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_85 <= _GEN_2400;
        end else begin
          ram_1_85 <= _GEN_12549;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_86 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_86 <= _GEN_2401;
        end else begin
          ram_1_86 <= _GEN_12550;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_87 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_87 <= _GEN_2402;
        end else begin
          ram_1_87 <= _GEN_12551;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_88 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_88 <= _GEN_2403;
        end else begin
          ram_1_88 <= _GEN_12552;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_89 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_89 <= _GEN_2404;
        end else begin
          ram_1_89 <= _GEN_12553;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_90 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_90 <= _GEN_2405;
        end else begin
          ram_1_90 <= _GEN_12554;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_91 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_91 <= _GEN_2406;
        end else begin
          ram_1_91 <= _GEN_12555;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_92 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_92 <= _GEN_2407;
        end else begin
          ram_1_92 <= _GEN_12556;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_93 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_93 <= _GEN_2408;
        end else begin
          ram_1_93 <= _GEN_12557;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_94 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_94 <= _GEN_2409;
        end else begin
          ram_1_94 <= _GEN_12558;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_95 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_95 <= _GEN_2410;
        end else begin
          ram_1_95 <= _GEN_12559;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_96 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_96 <= _GEN_2411;
        end else begin
          ram_1_96 <= _GEN_12560;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_97 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_97 <= _GEN_2412;
        end else begin
          ram_1_97 <= _GEN_12561;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_98 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_98 <= _GEN_2413;
        end else begin
          ram_1_98 <= _GEN_12562;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_99 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_99 <= _GEN_2414;
        end else begin
          ram_1_99 <= _GEN_12563;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_100 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_100 <= _GEN_2415;
        end else begin
          ram_1_100 <= _GEN_12564;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_101 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_101 <= _GEN_2416;
        end else begin
          ram_1_101 <= _GEN_12565;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_102 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_102 <= _GEN_2417;
        end else begin
          ram_1_102 <= _GEN_12566;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_103 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_103 <= _GEN_2418;
        end else begin
          ram_1_103 <= _GEN_12567;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_104 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_104 <= _GEN_2419;
        end else begin
          ram_1_104 <= _GEN_12568;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_105 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_105 <= _GEN_2420;
        end else begin
          ram_1_105 <= _GEN_12569;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_106 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_106 <= _GEN_2421;
        end else begin
          ram_1_106 <= _GEN_12570;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_107 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_107 <= _GEN_2422;
        end else begin
          ram_1_107 <= _GEN_12571;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_108 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_108 <= _GEN_2423;
        end else begin
          ram_1_108 <= _GEN_12572;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_109 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_109 <= _GEN_2424;
        end else begin
          ram_1_109 <= _GEN_12573;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_110 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_110 <= _GEN_2425;
        end else begin
          ram_1_110 <= _GEN_12574;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_111 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_111 <= _GEN_2426;
        end else begin
          ram_1_111 <= _GEN_12575;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_112 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_112 <= _GEN_2427;
        end else begin
          ram_1_112 <= _GEN_12576;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_113 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_113 <= _GEN_2428;
        end else begin
          ram_1_113 <= _GEN_12577;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_114 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_114 <= _GEN_2429;
        end else begin
          ram_1_114 <= _GEN_12578;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_115 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_115 <= _GEN_2430;
        end else begin
          ram_1_115 <= _GEN_12579;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_116 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_116 <= _GEN_2431;
        end else begin
          ram_1_116 <= _GEN_12580;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_117 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_117 <= _GEN_2432;
        end else begin
          ram_1_117 <= _GEN_12581;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_118 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_118 <= _GEN_2433;
        end else begin
          ram_1_118 <= _GEN_12582;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_119 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_119 <= _GEN_2434;
        end else begin
          ram_1_119 <= _GEN_12583;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_120 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_120 <= _GEN_2435;
        end else begin
          ram_1_120 <= _GEN_12584;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_121 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_121 <= _GEN_2436;
        end else begin
          ram_1_121 <= _GEN_12585;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_122 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_122 <= _GEN_2437;
        end else begin
          ram_1_122 <= _GEN_12586;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_123 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_123 <= _GEN_2438;
        end else begin
          ram_1_123 <= _GEN_12587;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_124 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_124 <= _GEN_2439;
        end else begin
          ram_1_124 <= _GEN_12588;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_125 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_125 <= _GEN_2440;
        end else begin
          ram_1_125 <= _GEN_12589;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_126 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_126 <= _GEN_2441;
        end else begin
          ram_1_126 <= _GEN_12590;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_1_127 <= 64'h0; // @[d_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          ram_1_127 <= _GEN_2442;
        end else begin
          ram_1_127 <= _GEN_12591;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_0 <= _GEN_12207;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_1 <= _GEN_12208;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_2 <= _GEN_12209;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_3 <= _GEN_12210;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_4 <= _GEN_12211;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_5 <= _GEN_12212;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_6 <= _GEN_12213;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_7 <= _GEN_12214;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_8 <= _GEN_12215;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_9 <= _GEN_12216;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_10 <= _GEN_12217;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_11 <= _GEN_12218;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_12 <= _GEN_12219;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_13 <= _GEN_12220;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_14 <= _GEN_12221;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_15 <= _GEN_12222;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_16 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_16 <= _GEN_12223;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_17 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_17 <= _GEN_12224;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_18 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_18 <= _GEN_12225;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_19 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_19 <= _GEN_12226;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_20 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_20 <= _GEN_12227;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_21 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_21 <= _GEN_12228;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_22 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_22 <= _GEN_12229;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_23 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_23 <= _GEN_12230;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_24 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_24 <= _GEN_12231;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_25 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_25 <= _GEN_12232;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_26 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_26 <= _GEN_12233;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_27 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_27 <= _GEN_12234;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_28 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_28 <= _GEN_12235;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_29 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_29 <= _GEN_12236;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_30 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_30 <= _GEN_12237;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_31 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_31 <= _GEN_12238;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_32 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_32 <= _GEN_12239;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_33 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_33 <= _GEN_12240;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_34 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_34 <= _GEN_12241;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_35 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_35 <= _GEN_12242;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_36 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_36 <= _GEN_12243;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_37 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_37 <= _GEN_12244;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_38 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_38 <= _GEN_12245;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_39 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_39 <= _GEN_12246;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_40 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_40 <= _GEN_12247;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_41 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_41 <= _GEN_12248;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_42 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_42 <= _GEN_12249;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_43 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_43 <= _GEN_12250;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_44 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_44 <= _GEN_12251;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_45 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_45 <= _GEN_12252;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_46 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_46 <= _GEN_12253;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_47 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_47 <= _GEN_12254;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_48 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_48 <= _GEN_12255;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_49 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_49 <= _GEN_12256;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_50 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_50 <= _GEN_12257;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_51 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_51 <= _GEN_12258;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_52 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_52 <= _GEN_12259;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_53 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_53 <= _GEN_12260;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_54 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_54 <= _GEN_12261;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_55 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_55 <= _GEN_12262;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_56 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_56 <= _GEN_12263;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_57 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_57 <= _GEN_12264;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_58 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_58 <= _GEN_12265;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_59 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_59 <= _GEN_12266;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_60 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_60 <= _GEN_12267;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_61 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_61 <= _GEN_12268;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_62 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_62 <= _GEN_12269;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_63 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_63 <= _GEN_12270;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_64 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_64 <= _GEN_12271;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_65 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_65 <= _GEN_12272;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_66 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_66 <= _GEN_12273;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_67 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_67 <= _GEN_12274;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_68 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_68 <= _GEN_12275;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_69 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_69 <= _GEN_12276;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_70 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_70 <= _GEN_12277;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_71 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_71 <= _GEN_12278;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_72 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_72 <= _GEN_12279;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_73 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_73 <= _GEN_12280;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_74 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_74 <= _GEN_12281;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_75 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_75 <= _GEN_12282;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_76 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_76 <= _GEN_12283;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_77 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_77 <= _GEN_12284;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_78 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_78 <= _GEN_12285;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_79 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_79 <= _GEN_12286;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_80 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_80 <= _GEN_12287;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_81 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_81 <= _GEN_12288;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_82 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_82 <= _GEN_12289;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_83 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_83 <= _GEN_12290;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_84 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_84 <= _GEN_12291;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_85 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_85 <= _GEN_12292;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_86 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_86 <= _GEN_12293;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_87 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_87 <= _GEN_12294;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_88 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_88 <= _GEN_12295;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_89 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_89 <= _GEN_12296;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_90 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_90 <= _GEN_12297;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_91 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_91 <= _GEN_12298;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_92 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_92 <= _GEN_12299;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_93 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_93 <= _GEN_12300;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_94 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_94 <= _GEN_12301;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_95 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_95 <= _GEN_12302;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_96 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_96 <= _GEN_12303;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_97 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_97 <= _GEN_12304;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_98 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_98 <= _GEN_12305;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_99 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_99 <= _GEN_12306;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_100 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_100 <= _GEN_12307;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_101 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_101 <= _GEN_12308;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_102 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_102 <= _GEN_12309;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_103 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_103 <= _GEN_12310;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_104 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_104 <= _GEN_12311;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_105 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_105 <= _GEN_12312;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_106 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_106 <= _GEN_12313;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_107 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_107 <= _GEN_12314;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_108 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_108 <= _GEN_12315;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_109 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_109 <= _GEN_12316;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_110 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_110 <= _GEN_12317;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_111 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_111 <= _GEN_12318;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_112 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_112 <= _GEN_12319;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_113 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_113 <= _GEN_12320;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_114 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_114 <= _GEN_12321;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_115 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_115 <= _GEN_12322;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_116 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_116 <= _GEN_12323;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_117 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_117 <= _GEN_12324;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_118 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_118 <= _GEN_12325;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_119 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_119 <= _GEN_12326;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_120 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_120 <= _GEN_12327;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_121 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_121 <= _GEN_12328;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_122 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_122 <= _GEN_12329;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_123 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_123 <= _GEN_12330;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_124 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_124 <= _GEN_12331;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_125 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_125 <= _GEN_12332;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_126 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_126 <= _GEN_12333;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      tag_0_127 <= 32'h0; // @[d_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_0_127 <= _GEN_12334;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_0 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_0 <= _GEN_12592;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_1 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_1 <= _GEN_12593;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_2 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_2 <= _GEN_12594;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_3 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_3 <= _GEN_12595;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_4 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_4 <= _GEN_12596;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_5 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_5 <= _GEN_12597;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_6 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_6 <= _GEN_12598;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_7 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_7 <= _GEN_12599;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_8 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_8 <= _GEN_12600;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_9 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_9 <= _GEN_12601;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_10 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_10 <= _GEN_12602;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_11 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_11 <= _GEN_12603;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_12 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_12 <= _GEN_12604;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_13 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_13 <= _GEN_12605;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_14 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_14 <= _GEN_12606;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_15 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_15 <= _GEN_12607;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_16 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_16 <= _GEN_12608;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_17 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_17 <= _GEN_12609;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_18 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_18 <= _GEN_12610;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_19 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_19 <= _GEN_12611;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_20 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_20 <= _GEN_12612;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_21 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_21 <= _GEN_12613;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_22 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_22 <= _GEN_12614;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_23 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_23 <= _GEN_12615;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_24 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_24 <= _GEN_12616;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_25 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_25 <= _GEN_12617;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_26 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_26 <= _GEN_12618;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_27 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_27 <= _GEN_12619;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_28 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_28 <= _GEN_12620;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_29 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_29 <= _GEN_12621;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_30 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_30 <= _GEN_12622;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_31 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_31 <= _GEN_12623;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_32 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_32 <= _GEN_12624;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_33 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_33 <= _GEN_12625;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_34 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_34 <= _GEN_12626;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_35 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_35 <= _GEN_12627;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_36 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_36 <= _GEN_12628;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_37 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_37 <= _GEN_12629;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_38 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_38 <= _GEN_12630;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_39 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_39 <= _GEN_12631;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_40 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_40 <= _GEN_12632;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_41 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_41 <= _GEN_12633;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_42 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_42 <= _GEN_12634;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_43 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_43 <= _GEN_12635;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_44 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_44 <= _GEN_12636;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_45 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_45 <= _GEN_12637;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_46 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_46 <= _GEN_12638;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_47 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_47 <= _GEN_12639;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_48 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_48 <= _GEN_12640;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_49 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_49 <= _GEN_12641;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_50 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_50 <= _GEN_12642;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_51 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_51 <= _GEN_12643;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_52 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_52 <= _GEN_12644;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_53 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_53 <= _GEN_12645;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_54 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_54 <= _GEN_12646;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_55 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_55 <= _GEN_12647;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_56 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_56 <= _GEN_12648;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_57 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_57 <= _GEN_12649;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_58 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_58 <= _GEN_12650;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_59 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_59 <= _GEN_12651;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_60 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_60 <= _GEN_12652;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_61 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_61 <= _GEN_12653;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_62 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_62 <= _GEN_12654;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_63 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_63 <= _GEN_12655;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_64 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_64 <= _GEN_12656;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_65 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_65 <= _GEN_12657;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_66 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_66 <= _GEN_12658;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_67 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_67 <= _GEN_12659;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_68 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_68 <= _GEN_12660;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_69 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_69 <= _GEN_12661;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_70 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_70 <= _GEN_12662;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_71 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_71 <= _GEN_12663;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_72 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_72 <= _GEN_12664;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_73 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_73 <= _GEN_12665;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_74 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_74 <= _GEN_12666;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_75 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_75 <= _GEN_12667;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_76 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_76 <= _GEN_12668;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_77 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_77 <= _GEN_12669;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_78 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_78 <= _GEN_12670;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_79 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_79 <= _GEN_12671;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_80 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_80 <= _GEN_12672;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_81 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_81 <= _GEN_12673;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_82 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_82 <= _GEN_12674;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_83 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_83 <= _GEN_12675;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_84 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_84 <= _GEN_12676;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_85 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_85 <= _GEN_12677;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_86 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_86 <= _GEN_12678;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_87 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_87 <= _GEN_12679;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_88 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_88 <= _GEN_12680;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_89 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_89 <= _GEN_12681;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_90 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_90 <= _GEN_12682;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_91 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_91 <= _GEN_12683;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_92 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_92 <= _GEN_12684;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_93 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_93 <= _GEN_12685;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_94 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_94 <= _GEN_12686;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_95 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_95 <= _GEN_12687;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_96 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_96 <= _GEN_12688;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_97 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_97 <= _GEN_12689;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_98 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_98 <= _GEN_12690;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_99 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_99 <= _GEN_12691;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_100 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_100 <= _GEN_12692;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_101 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_101 <= _GEN_12693;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_102 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_102 <= _GEN_12694;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_103 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_103 <= _GEN_12695;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_104 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_104 <= _GEN_12696;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_105 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_105 <= _GEN_12697;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_106 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_106 <= _GEN_12698;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_107 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_107 <= _GEN_12699;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_108 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_108 <= _GEN_12700;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_109 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_109 <= _GEN_12701;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_110 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_110 <= _GEN_12702;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_111 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_111 <= _GEN_12703;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_112 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_112 <= _GEN_12704;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_113 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_113 <= _GEN_12705;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_114 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_114 <= _GEN_12706;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_115 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_115 <= _GEN_12707;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_116 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_116 <= _GEN_12708;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_117 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_117 <= _GEN_12709;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_118 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_118 <= _GEN_12710;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_119 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_119 <= _GEN_12711;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_120 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_120 <= _GEN_12712;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_121 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_121 <= _GEN_12713;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_122 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_122 <= _GEN_12714;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_123 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_123 <= _GEN_12715;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_124 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_124 <= _GEN_12716;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_125 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_125 <= _GEN_12717;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_126 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_126 <= _GEN_12718;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      tag_1_127 <= 32'h0; // @[d_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          tag_1_127 <= _GEN_12719;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_0 <= _GEN_12335;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_1 <= _GEN_12336;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_2 <= _GEN_12337;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_3 <= _GEN_12338;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_4 <= _GEN_12339;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_5 <= _GEN_12340;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_6 <= _GEN_12341;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_7 <= _GEN_12342;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_8 <= _GEN_12343;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_9 <= _GEN_12344;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_10 <= _GEN_12345;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_11 <= _GEN_12346;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_12 <= _GEN_12347;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_13 <= _GEN_12348;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_14 <= _GEN_12349;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_15 <= _GEN_12350;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_16 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_16 <= _GEN_12351;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_17 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_17 <= _GEN_12352;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_18 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_18 <= _GEN_12353;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_19 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_19 <= _GEN_12354;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_20 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_20 <= _GEN_12355;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_21 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_21 <= _GEN_12356;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_22 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_22 <= _GEN_12357;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_23 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_23 <= _GEN_12358;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_24 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_24 <= _GEN_12359;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_25 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_25 <= _GEN_12360;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_26 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_26 <= _GEN_12361;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_27 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_27 <= _GEN_12362;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_28 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_28 <= _GEN_12363;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_29 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_29 <= _GEN_12364;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_30 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_30 <= _GEN_12365;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_31 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_31 <= _GEN_12366;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_32 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_32 <= _GEN_12367;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_33 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_33 <= _GEN_12368;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_34 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_34 <= _GEN_12369;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_35 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_35 <= _GEN_12370;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_36 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_36 <= _GEN_12371;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_37 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_37 <= _GEN_12372;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_38 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_38 <= _GEN_12373;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_39 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_39 <= _GEN_12374;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_40 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_40 <= _GEN_12375;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_41 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_41 <= _GEN_12376;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_42 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_42 <= _GEN_12377;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_43 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_43 <= _GEN_12378;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_44 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_44 <= _GEN_12379;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_45 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_45 <= _GEN_12380;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_46 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_46 <= _GEN_12381;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_47 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_47 <= _GEN_12382;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_48 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_48 <= _GEN_12383;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_49 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_49 <= _GEN_12384;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_50 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_50 <= _GEN_12385;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_51 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_51 <= _GEN_12386;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_52 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_52 <= _GEN_12387;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_53 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_53 <= _GEN_12388;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_54 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_54 <= _GEN_12389;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_55 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_55 <= _GEN_12390;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_56 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_56 <= _GEN_12391;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_57 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_57 <= _GEN_12392;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_58 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_58 <= _GEN_12393;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_59 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_59 <= _GEN_12394;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_60 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_60 <= _GEN_12395;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_61 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_61 <= _GEN_12396;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_62 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_62 <= _GEN_12397;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_63 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_63 <= _GEN_12398;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_64 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_64 <= _GEN_12399;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_65 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_65 <= _GEN_12400;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_66 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_66 <= _GEN_12401;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_67 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_67 <= _GEN_12402;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_68 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_68 <= _GEN_12403;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_69 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_69 <= _GEN_12404;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_70 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_70 <= _GEN_12405;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_71 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_71 <= _GEN_12406;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_72 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_72 <= _GEN_12407;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_73 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_73 <= _GEN_12408;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_74 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_74 <= _GEN_12409;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_75 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_75 <= _GEN_12410;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_76 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_76 <= _GEN_12411;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_77 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_77 <= _GEN_12412;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_78 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_78 <= _GEN_12413;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_79 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_79 <= _GEN_12414;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_80 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_80 <= _GEN_12415;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_81 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_81 <= _GEN_12416;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_82 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_82 <= _GEN_12417;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_83 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_83 <= _GEN_12418;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_84 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_84 <= _GEN_12419;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_85 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_85 <= _GEN_12420;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_86 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_86 <= _GEN_12421;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_87 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_87 <= _GEN_12422;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_88 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_88 <= _GEN_12423;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_89 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_89 <= _GEN_12424;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_90 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_90 <= _GEN_12425;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_91 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_91 <= _GEN_12426;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_92 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_92 <= _GEN_12427;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_93 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_93 <= _GEN_12428;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_94 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_94 <= _GEN_12429;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_95 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_95 <= _GEN_12430;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_96 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_96 <= _GEN_12431;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_97 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_97 <= _GEN_12432;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_98 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_98 <= _GEN_12433;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_99 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_99 <= _GEN_12434;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_100 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_100 <= _GEN_12435;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_101 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_101 <= _GEN_12436;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_102 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_102 <= _GEN_12437;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_103 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_103 <= _GEN_12438;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_104 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_104 <= _GEN_12439;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_105 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_105 <= _GEN_12440;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_106 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_106 <= _GEN_12441;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_107 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_107 <= _GEN_12442;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_108 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_108 <= _GEN_12443;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_109 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_109 <= _GEN_12444;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_110 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_110 <= _GEN_12445;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_111 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_111 <= _GEN_12446;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_112 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_112 <= _GEN_12447;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_113 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_113 <= _GEN_12448;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_114 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_114 <= _GEN_12449;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_115 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_115 <= _GEN_12450;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_116 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_116 <= _GEN_12451;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_117 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_117 <= _GEN_12452;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_118 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_118 <= _GEN_12453;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_119 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_119 <= _GEN_12454;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_120 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_120 <= _GEN_12455;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_121 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_121 <= _GEN_12456;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_122 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_122 <= _GEN_12457;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_123 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_123 <= _GEN_12458;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_124 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_124 <= _GEN_12459;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_125 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_125 <= _GEN_12460;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_126 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_126 <= _GEN_12461;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:26]
      valid_0_127 <= 1'h0; // @[d_cache.scala 22:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_0_127 <= _GEN_12462;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_0 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_0 <= _GEN_12720;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_1 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_1 <= _GEN_12721;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_2 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_2 <= _GEN_12722;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_3 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_3 <= _GEN_12723;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_4 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_4 <= _GEN_12724;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_5 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_5 <= _GEN_12725;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_6 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_6 <= _GEN_12726;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_7 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_7 <= _GEN_12727;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_8 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_8 <= _GEN_12728;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_9 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_9 <= _GEN_12729;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_10 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_10 <= _GEN_12730;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_11 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_11 <= _GEN_12731;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_12 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_12 <= _GEN_12732;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_13 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_13 <= _GEN_12733;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_14 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_14 <= _GEN_12734;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_15 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_15 <= _GEN_12735;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_16 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_16 <= _GEN_12736;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_17 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_17 <= _GEN_12737;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_18 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_18 <= _GEN_12738;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_19 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_19 <= _GEN_12739;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_20 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_20 <= _GEN_12740;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_21 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_21 <= _GEN_12741;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_22 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_22 <= _GEN_12742;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_23 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_23 <= _GEN_12743;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_24 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_24 <= _GEN_12744;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_25 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_25 <= _GEN_12745;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_26 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_26 <= _GEN_12746;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_27 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_27 <= _GEN_12747;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_28 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_28 <= _GEN_12748;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_29 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_29 <= _GEN_12749;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_30 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_30 <= _GEN_12750;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_31 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_31 <= _GEN_12751;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_32 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_32 <= _GEN_12752;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_33 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_33 <= _GEN_12753;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_34 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_34 <= _GEN_12754;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_35 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_35 <= _GEN_12755;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_36 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_36 <= _GEN_12756;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_37 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_37 <= _GEN_12757;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_38 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_38 <= _GEN_12758;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_39 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_39 <= _GEN_12759;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_40 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_40 <= _GEN_12760;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_41 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_41 <= _GEN_12761;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_42 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_42 <= _GEN_12762;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_43 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_43 <= _GEN_12763;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_44 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_44 <= _GEN_12764;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_45 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_45 <= _GEN_12765;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_46 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_46 <= _GEN_12766;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_47 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_47 <= _GEN_12767;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_48 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_48 <= _GEN_12768;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_49 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_49 <= _GEN_12769;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_50 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_50 <= _GEN_12770;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_51 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_51 <= _GEN_12771;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_52 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_52 <= _GEN_12772;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_53 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_53 <= _GEN_12773;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_54 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_54 <= _GEN_12774;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_55 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_55 <= _GEN_12775;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_56 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_56 <= _GEN_12776;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_57 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_57 <= _GEN_12777;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_58 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_58 <= _GEN_12778;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_59 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_59 <= _GEN_12779;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_60 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_60 <= _GEN_12780;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_61 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_61 <= _GEN_12781;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_62 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_62 <= _GEN_12782;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_63 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_63 <= _GEN_12783;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_64 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_64 <= _GEN_12784;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_65 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_65 <= _GEN_12785;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_66 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_66 <= _GEN_12786;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_67 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_67 <= _GEN_12787;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_68 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_68 <= _GEN_12788;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_69 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_69 <= _GEN_12789;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_70 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_70 <= _GEN_12790;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_71 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_71 <= _GEN_12791;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_72 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_72 <= _GEN_12792;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_73 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_73 <= _GEN_12793;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_74 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_74 <= _GEN_12794;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_75 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_75 <= _GEN_12795;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_76 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_76 <= _GEN_12796;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_77 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_77 <= _GEN_12797;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_78 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_78 <= _GEN_12798;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_79 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_79 <= _GEN_12799;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_80 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_80 <= _GEN_12800;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_81 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_81 <= _GEN_12801;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_82 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_82 <= _GEN_12802;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_83 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_83 <= _GEN_12803;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_84 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_84 <= _GEN_12804;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_85 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_85 <= _GEN_12805;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_86 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_86 <= _GEN_12806;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_87 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_87 <= _GEN_12807;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_88 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_88 <= _GEN_12808;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_89 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_89 <= _GEN_12809;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_90 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_90 <= _GEN_12810;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_91 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_91 <= _GEN_12811;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_92 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_92 <= _GEN_12812;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_93 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_93 <= _GEN_12813;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_94 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_94 <= _GEN_12814;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_95 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_95 <= _GEN_12815;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_96 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_96 <= _GEN_12816;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_97 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_97 <= _GEN_12817;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_98 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_98 <= _GEN_12818;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_99 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_99 <= _GEN_12819;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_100 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_100 <= _GEN_12820;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_101 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_101 <= _GEN_12821;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_102 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_102 <= _GEN_12822;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_103 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_103 <= _GEN_12823;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_104 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_104 <= _GEN_12824;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_105 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_105 <= _GEN_12825;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_106 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_106 <= _GEN_12826;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_107 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_107 <= _GEN_12827;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_108 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_108 <= _GEN_12828;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_109 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_109 <= _GEN_12829;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_110 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_110 <= _GEN_12830;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_111 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_111 <= _GEN_12831;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_112 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_112 <= _GEN_12832;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_113 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_113 <= _GEN_12833;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_114 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_114 <= _GEN_12834;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_115 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_115 <= _GEN_12835;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_116 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_116 <= _GEN_12836;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_117 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_117 <= _GEN_12837;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_118 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_118 <= _GEN_12838;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_119 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_119 <= _GEN_12839;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_120 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_120 <= _GEN_12840;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_121 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_121 <= _GEN_12841;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_122 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_122 <= _GEN_12842;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_123 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_123 <= _GEN_12843;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_124 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_124 <= _GEN_12844;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_125 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_125 <= _GEN_12845;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_126 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_126 <= _GEN_12846;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:26]
      valid_1_127 <= 1'h0; // @[d_cache.scala 23:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          valid_1_127 <= _GEN_12847;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_0 <= _GEN_2187;
        end else begin
          dirty_0_0 <= _GEN_12850;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_1 <= _GEN_2188;
        end else begin
          dirty_0_1 <= _GEN_12851;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_2 <= _GEN_2189;
        end else begin
          dirty_0_2 <= _GEN_12852;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_3 <= _GEN_2190;
        end else begin
          dirty_0_3 <= _GEN_12853;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_4 <= _GEN_2191;
        end else begin
          dirty_0_4 <= _GEN_12854;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_5 <= _GEN_2192;
        end else begin
          dirty_0_5 <= _GEN_12855;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_6 <= _GEN_2193;
        end else begin
          dirty_0_6 <= _GEN_12856;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_7 <= _GEN_2194;
        end else begin
          dirty_0_7 <= _GEN_12857;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_8 <= _GEN_2195;
        end else begin
          dirty_0_8 <= _GEN_12858;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_9 <= _GEN_2196;
        end else begin
          dirty_0_9 <= _GEN_12859;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_10 <= _GEN_2197;
        end else begin
          dirty_0_10 <= _GEN_12860;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_11 <= _GEN_2198;
        end else begin
          dirty_0_11 <= _GEN_12861;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_12 <= _GEN_2199;
        end else begin
          dirty_0_12 <= _GEN_12862;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_13 <= _GEN_2200;
        end else begin
          dirty_0_13 <= _GEN_12863;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_14 <= _GEN_2201;
        end else begin
          dirty_0_14 <= _GEN_12864;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_15 <= _GEN_2202;
        end else begin
          dirty_0_15 <= _GEN_12865;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_16 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_16 <= _GEN_2203;
        end else begin
          dirty_0_16 <= _GEN_12866;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_17 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_17 <= _GEN_2204;
        end else begin
          dirty_0_17 <= _GEN_12867;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_18 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_18 <= _GEN_2205;
        end else begin
          dirty_0_18 <= _GEN_12868;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_19 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_19 <= _GEN_2206;
        end else begin
          dirty_0_19 <= _GEN_12869;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_20 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_20 <= _GEN_2207;
        end else begin
          dirty_0_20 <= _GEN_12870;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_21 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_21 <= _GEN_2208;
        end else begin
          dirty_0_21 <= _GEN_12871;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_22 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_22 <= _GEN_2209;
        end else begin
          dirty_0_22 <= _GEN_12872;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_23 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_23 <= _GEN_2210;
        end else begin
          dirty_0_23 <= _GEN_12873;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_24 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_24 <= _GEN_2211;
        end else begin
          dirty_0_24 <= _GEN_12874;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_25 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_25 <= _GEN_2212;
        end else begin
          dirty_0_25 <= _GEN_12875;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_26 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_26 <= _GEN_2213;
        end else begin
          dirty_0_26 <= _GEN_12876;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_27 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_27 <= _GEN_2214;
        end else begin
          dirty_0_27 <= _GEN_12877;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_28 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_28 <= _GEN_2215;
        end else begin
          dirty_0_28 <= _GEN_12878;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_29 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_29 <= _GEN_2216;
        end else begin
          dirty_0_29 <= _GEN_12879;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_30 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_30 <= _GEN_2217;
        end else begin
          dirty_0_30 <= _GEN_12880;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_31 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_31 <= _GEN_2218;
        end else begin
          dirty_0_31 <= _GEN_12881;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_32 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_32 <= _GEN_2219;
        end else begin
          dirty_0_32 <= _GEN_12882;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_33 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_33 <= _GEN_2220;
        end else begin
          dirty_0_33 <= _GEN_12883;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_34 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_34 <= _GEN_2221;
        end else begin
          dirty_0_34 <= _GEN_12884;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_35 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_35 <= _GEN_2222;
        end else begin
          dirty_0_35 <= _GEN_12885;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_36 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_36 <= _GEN_2223;
        end else begin
          dirty_0_36 <= _GEN_12886;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_37 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_37 <= _GEN_2224;
        end else begin
          dirty_0_37 <= _GEN_12887;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_38 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_38 <= _GEN_2225;
        end else begin
          dirty_0_38 <= _GEN_12888;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_39 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_39 <= _GEN_2226;
        end else begin
          dirty_0_39 <= _GEN_12889;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_40 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_40 <= _GEN_2227;
        end else begin
          dirty_0_40 <= _GEN_12890;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_41 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_41 <= _GEN_2228;
        end else begin
          dirty_0_41 <= _GEN_12891;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_42 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_42 <= _GEN_2229;
        end else begin
          dirty_0_42 <= _GEN_12892;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_43 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_43 <= _GEN_2230;
        end else begin
          dirty_0_43 <= _GEN_12893;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_44 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_44 <= _GEN_2231;
        end else begin
          dirty_0_44 <= _GEN_12894;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_45 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_45 <= _GEN_2232;
        end else begin
          dirty_0_45 <= _GEN_12895;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_46 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_46 <= _GEN_2233;
        end else begin
          dirty_0_46 <= _GEN_12896;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_47 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_47 <= _GEN_2234;
        end else begin
          dirty_0_47 <= _GEN_12897;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_48 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_48 <= _GEN_2235;
        end else begin
          dirty_0_48 <= _GEN_12898;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_49 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_49 <= _GEN_2236;
        end else begin
          dirty_0_49 <= _GEN_12899;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_50 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_50 <= _GEN_2237;
        end else begin
          dirty_0_50 <= _GEN_12900;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_51 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_51 <= _GEN_2238;
        end else begin
          dirty_0_51 <= _GEN_12901;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_52 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_52 <= _GEN_2239;
        end else begin
          dirty_0_52 <= _GEN_12902;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_53 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_53 <= _GEN_2240;
        end else begin
          dirty_0_53 <= _GEN_12903;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_54 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_54 <= _GEN_2241;
        end else begin
          dirty_0_54 <= _GEN_12904;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_55 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_55 <= _GEN_2242;
        end else begin
          dirty_0_55 <= _GEN_12905;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_56 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_56 <= _GEN_2243;
        end else begin
          dirty_0_56 <= _GEN_12906;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_57 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_57 <= _GEN_2244;
        end else begin
          dirty_0_57 <= _GEN_12907;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_58 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_58 <= _GEN_2245;
        end else begin
          dirty_0_58 <= _GEN_12908;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_59 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_59 <= _GEN_2246;
        end else begin
          dirty_0_59 <= _GEN_12909;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_60 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_60 <= _GEN_2247;
        end else begin
          dirty_0_60 <= _GEN_12910;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_61 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_61 <= _GEN_2248;
        end else begin
          dirty_0_61 <= _GEN_12911;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_62 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_62 <= _GEN_2249;
        end else begin
          dirty_0_62 <= _GEN_12912;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_63 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_63 <= _GEN_2250;
        end else begin
          dirty_0_63 <= _GEN_12913;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_64 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_64 <= _GEN_2251;
        end else begin
          dirty_0_64 <= _GEN_12914;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_65 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_65 <= _GEN_2252;
        end else begin
          dirty_0_65 <= _GEN_12915;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_66 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_66 <= _GEN_2253;
        end else begin
          dirty_0_66 <= _GEN_12916;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_67 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_67 <= _GEN_2254;
        end else begin
          dirty_0_67 <= _GEN_12917;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_68 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_68 <= _GEN_2255;
        end else begin
          dirty_0_68 <= _GEN_12918;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_69 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_69 <= _GEN_2256;
        end else begin
          dirty_0_69 <= _GEN_12919;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_70 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_70 <= _GEN_2257;
        end else begin
          dirty_0_70 <= _GEN_12920;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_71 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_71 <= _GEN_2258;
        end else begin
          dirty_0_71 <= _GEN_12921;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_72 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_72 <= _GEN_2259;
        end else begin
          dirty_0_72 <= _GEN_12922;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_73 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_73 <= _GEN_2260;
        end else begin
          dirty_0_73 <= _GEN_12923;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_74 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_74 <= _GEN_2261;
        end else begin
          dirty_0_74 <= _GEN_12924;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_75 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_75 <= _GEN_2262;
        end else begin
          dirty_0_75 <= _GEN_12925;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_76 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_76 <= _GEN_2263;
        end else begin
          dirty_0_76 <= _GEN_12926;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_77 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_77 <= _GEN_2264;
        end else begin
          dirty_0_77 <= _GEN_12927;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_78 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_78 <= _GEN_2265;
        end else begin
          dirty_0_78 <= _GEN_12928;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_79 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_79 <= _GEN_2266;
        end else begin
          dirty_0_79 <= _GEN_12929;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_80 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_80 <= _GEN_2267;
        end else begin
          dirty_0_80 <= _GEN_12930;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_81 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_81 <= _GEN_2268;
        end else begin
          dirty_0_81 <= _GEN_12931;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_82 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_82 <= _GEN_2269;
        end else begin
          dirty_0_82 <= _GEN_12932;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_83 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_83 <= _GEN_2270;
        end else begin
          dirty_0_83 <= _GEN_12933;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_84 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_84 <= _GEN_2271;
        end else begin
          dirty_0_84 <= _GEN_12934;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_85 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_85 <= _GEN_2272;
        end else begin
          dirty_0_85 <= _GEN_12935;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_86 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_86 <= _GEN_2273;
        end else begin
          dirty_0_86 <= _GEN_12936;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_87 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_87 <= _GEN_2274;
        end else begin
          dirty_0_87 <= _GEN_12937;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_88 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_88 <= _GEN_2275;
        end else begin
          dirty_0_88 <= _GEN_12938;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_89 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_89 <= _GEN_2276;
        end else begin
          dirty_0_89 <= _GEN_12939;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_90 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_90 <= _GEN_2277;
        end else begin
          dirty_0_90 <= _GEN_12940;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_91 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_91 <= _GEN_2278;
        end else begin
          dirty_0_91 <= _GEN_12941;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_92 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_92 <= _GEN_2279;
        end else begin
          dirty_0_92 <= _GEN_12942;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_93 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_93 <= _GEN_2280;
        end else begin
          dirty_0_93 <= _GEN_12943;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_94 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_94 <= _GEN_2281;
        end else begin
          dirty_0_94 <= _GEN_12944;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_95 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_95 <= _GEN_2282;
        end else begin
          dirty_0_95 <= _GEN_12945;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_96 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_96 <= _GEN_2283;
        end else begin
          dirty_0_96 <= _GEN_12946;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_97 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_97 <= _GEN_2284;
        end else begin
          dirty_0_97 <= _GEN_12947;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_98 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_98 <= _GEN_2285;
        end else begin
          dirty_0_98 <= _GEN_12948;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_99 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_99 <= _GEN_2286;
        end else begin
          dirty_0_99 <= _GEN_12949;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_100 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_100 <= _GEN_2287;
        end else begin
          dirty_0_100 <= _GEN_12950;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_101 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_101 <= _GEN_2288;
        end else begin
          dirty_0_101 <= _GEN_12951;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_102 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_102 <= _GEN_2289;
        end else begin
          dirty_0_102 <= _GEN_12952;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_103 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_103 <= _GEN_2290;
        end else begin
          dirty_0_103 <= _GEN_12953;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_104 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_104 <= _GEN_2291;
        end else begin
          dirty_0_104 <= _GEN_12954;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_105 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_105 <= _GEN_2292;
        end else begin
          dirty_0_105 <= _GEN_12955;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_106 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_106 <= _GEN_2293;
        end else begin
          dirty_0_106 <= _GEN_12956;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_107 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_107 <= _GEN_2294;
        end else begin
          dirty_0_107 <= _GEN_12957;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_108 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_108 <= _GEN_2295;
        end else begin
          dirty_0_108 <= _GEN_12958;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_109 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_109 <= _GEN_2296;
        end else begin
          dirty_0_109 <= _GEN_12959;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_110 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_110 <= _GEN_2297;
        end else begin
          dirty_0_110 <= _GEN_12960;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_111 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_111 <= _GEN_2298;
        end else begin
          dirty_0_111 <= _GEN_12961;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_112 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_112 <= _GEN_2299;
        end else begin
          dirty_0_112 <= _GEN_12962;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_113 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_113 <= _GEN_2300;
        end else begin
          dirty_0_113 <= _GEN_12963;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_114 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_114 <= _GEN_2301;
        end else begin
          dirty_0_114 <= _GEN_12964;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_115 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_115 <= _GEN_2302;
        end else begin
          dirty_0_115 <= _GEN_12965;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_116 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_116 <= _GEN_2303;
        end else begin
          dirty_0_116 <= _GEN_12966;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_117 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_117 <= _GEN_2304;
        end else begin
          dirty_0_117 <= _GEN_12967;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_118 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_118 <= _GEN_2305;
        end else begin
          dirty_0_118 <= _GEN_12968;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_119 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_119 <= _GEN_2306;
        end else begin
          dirty_0_119 <= _GEN_12969;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_120 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_120 <= _GEN_2307;
        end else begin
          dirty_0_120 <= _GEN_12970;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_121 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_121 <= _GEN_2308;
        end else begin
          dirty_0_121 <= _GEN_12971;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_122 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_122 <= _GEN_2309;
        end else begin
          dirty_0_122 <= _GEN_12972;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_123 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_123 <= _GEN_2310;
        end else begin
          dirty_0_123 <= _GEN_12973;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_124 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_124 <= _GEN_2311;
        end else begin
          dirty_0_124 <= _GEN_12974;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_125 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_125 <= _GEN_2312;
        end else begin
          dirty_0_125 <= _GEN_12975;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_126 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_126 <= _GEN_2313;
        end else begin
          dirty_0_126 <= _GEN_12976;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      dirty_0_127 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_0_127 <= _GEN_2314;
        end else begin
          dirty_0_127 <= _GEN_12977;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_0 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_0 <= _GEN_2443;
        end else begin
          dirty_1_0 <= _GEN_12978;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_1 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_1 <= _GEN_2444;
        end else begin
          dirty_1_1 <= _GEN_12979;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_2 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_2 <= _GEN_2445;
        end else begin
          dirty_1_2 <= _GEN_12980;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_3 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_3 <= _GEN_2446;
        end else begin
          dirty_1_3 <= _GEN_12981;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_4 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_4 <= _GEN_2447;
        end else begin
          dirty_1_4 <= _GEN_12982;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_5 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_5 <= _GEN_2448;
        end else begin
          dirty_1_5 <= _GEN_12983;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_6 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_6 <= _GEN_2449;
        end else begin
          dirty_1_6 <= _GEN_12984;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_7 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_7 <= _GEN_2450;
        end else begin
          dirty_1_7 <= _GEN_12985;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_8 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_8 <= _GEN_2451;
        end else begin
          dirty_1_8 <= _GEN_12986;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_9 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_9 <= _GEN_2452;
        end else begin
          dirty_1_9 <= _GEN_12987;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_10 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_10 <= _GEN_2453;
        end else begin
          dirty_1_10 <= _GEN_12988;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_11 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_11 <= _GEN_2454;
        end else begin
          dirty_1_11 <= _GEN_12989;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_12 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_12 <= _GEN_2455;
        end else begin
          dirty_1_12 <= _GEN_12990;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_13 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_13 <= _GEN_2456;
        end else begin
          dirty_1_13 <= _GEN_12991;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_14 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_14 <= _GEN_2457;
        end else begin
          dirty_1_14 <= _GEN_12992;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_15 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_15 <= _GEN_2458;
        end else begin
          dirty_1_15 <= _GEN_12993;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_16 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_16 <= _GEN_2459;
        end else begin
          dirty_1_16 <= _GEN_12994;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_17 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_17 <= _GEN_2460;
        end else begin
          dirty_1_17 <= _GEN_12995;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_18 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_18 <= _GEN_2461;
        end else begin
          dirty_1_18 <= _GEN_12996;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_19 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_19 <= _GEN_2462;
        end else begin
          dirty_1_19 <= _GEN_12997;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_20 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_20 <= _GEN_2463;
        end else begin
          dirty_1_20 <= _GEN_12998;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_21 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_21 <= _GEN_2464;
        end else begin
          dirty_1_21 <= _GEN_12999;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_22 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_22 <= _GEN_2465;
        end else begin
          dirty_1_22 <= _GEN_13000;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_23 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_23 <= _GEN_2466;
        end else begin
          dirty_1_23 <= _GEN_13001;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_24 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_24 <= _GEN_2467;
        end else begin
          dirty_1_24 <= _GEN_13002;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_25 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_25 <= _GEN_2468;
        end else begin
          dirty_1_25 <= _GEN_13003;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_26 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_26 <= _GEN_2469;
        end else begin
          dirty_1_26 <= _GEN_13004;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_27 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_27 <= _GEN_2470;
        end else begin
          dirty_1_27 <= _GEN_13005;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_28 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_28 <= _GEN_2471;
        end else begin
          dirty_1_28 <= _GEN_13006;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_29 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_29 <= _GEN_2472;
        end else begin
          dirty_1_29 <= _GEN_13007;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_30 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_30 <= _GEN_2473;
        end else begin
          dirty_1_30 <= _GEN_13008;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_31 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_31 <= _GEN_2474;
        end else begin
          dirty_1_31 <= _GEN_13009;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_32 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_32 <= _GEN_2475;
        end else begin
          dirty_1_32 <= _GEN_13010;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_33 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_33 <= _GEN_2476;
        end else begin
          dirty_1_33 <= _GEN_13011;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_34 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_34 <= _GEN_2477;
        end else begin
          dirty_1_34 <= _GEN_13012;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_35 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_35 <= _GEN_2478;
        end else begin
          dirty_1_35 <= _GEN_13013;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_36 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_36 <= _GEN_2479;
        end else begin
          dirty_1_36 <= _GEN_13014;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_37 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_37 <= _GEN_2480;
        end else begin
          dirty_1_37 <= _GEN_13015;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_38 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_38 <= _GEN_2481;
        end else begin
          dirty_1_38 <= _GEN_13016;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_39 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_39 <= _GEN_2482;
        end else begin
          dirty_1_39 <= _GEN_13017;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_40 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_40 <= _GEN_2483;
        end else begin
          dirty_1_40 <= _GEN_13018;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_41 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_41 <= _GEN_2484;
        end else begin
          dirty_1_41 <= _GEN_13019;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_42 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_42 <= _GEN_2485;
        end else begin
          dirty_1_42 <= _GEN_13020;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_43 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_43 <= _GEN_2486;
        end else begin
          dirty_1_43 <= _GEN_13021;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_44 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_44 <= _GEN_2487;
        end else begin
          dirty_1_44 <= _GEN_13022;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_45 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_45 <= _GEN_2488;
        end else begin
          dirty_1_45 <= _GEN_13023;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_46 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_46 <= _GEN_2489;
        end else begin
          dirty_1_46 <= _GEN_13024;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_47 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_47 <= _GEN_2490;
        end else begin
          dirty_1_47 <= _GEN_13025;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_48 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_48 <= _GEN_2491;
        end else begin
          dirty_1_48 <= _GEN_13026;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_49 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_49 <= _GEN_2492;
        end else begin
          dirty_1_49 <= _GEN_13027;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_50 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_50 <= _GEN_2493;
        end else begin
          dirty_1_50 <= _GEN_13028;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_51 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_51 <= _GEN_2494;
        end else begin
          dirty_1_51 <= _GEN_13029;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_52 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_52 <= _GEN_2495;
        end else begin
          dirty_1_52 <= _GEN_13030;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_53 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_53 <= _GEN_2496;
        end else begin
          dirty_1_53 <= _GEN_13031;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_54 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_54 <= _GEN_2497;
        end else begin
          dirty_1_54 <= _GEN_13032;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_55 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_55 <= _GEN_2498;
        end else begin
          dirty_1_55 <= _GEN_13033;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_56 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_56 <= _GEN_2499;
        end else begin
          dirty_1_56 <= _GEN_13034;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_57 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_57 <= _GEN_2500;
        end else begin
          dirty_1_57 <= _GEN_13035;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_58 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_58 <= _GEN_2501;
        end else begin
          dirty_1_58 <= _GEN_13036;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_59 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_59 <= _GEN_2502;
        end else begin
          dirty_1_59 <= _GEN_13037;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_60 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_60 <= _GEN_2503;
        end else begin
          dirty_1_60 <= _GEN_13038;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_61 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_61 <= _GEN_2504;
        end else begin
          dirty_1_61 <= _GEN_13039;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_62 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_62 <= _GEN_2505;
        end else begin
          dirty_1_62 <= _GEN_13040;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_63 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_63 <= _GEN_2506;
        end else begin
          dirty_1_63 <= _GEN_13041;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_64 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_64 <= _GEN_2507;
        end else begin
          dirty_1_64 <= _GEN_13042;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_65 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_65 <= _GEN_2508;
        end else begin
          dirty_1_65 <= _GEN_13043;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_66 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_66 <= _GEN_2509;
        end else begin
          dirty_1_66 <= _GEN_13044;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_67 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_67 <= _GEN_2510;
        end else begin
          dirty_1_67 <= _GEN_13045;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_68 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_68 <= _GEN_2511;
        end else begin
          dirty_1_68 <= _GEN_13046;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_69 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_69 <= _GEN_2512;
        end else begin
          dirty_1_69 <= _GEN_13047;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_70 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_70 <= _GEN_2513;
        end else begin
          dirty_1_70 <= _GEN_13048;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_71 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_71 <= _GEN_2514;
        end else begin
          dirty_1_71 <= _GEN_13049;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_72 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_72 <= _GEN_2515;
        end else begin
          dirty_1_72 <= _GEN_13050;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_73 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_73 <= _GEN_2516;
        end else begin
          dirty_1_73 <= _GEN_13051;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_74 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_74 <= _GEN_2517;
        end else begin
          dirty_1_74 <= _GEN_13052;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_75 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_75 <= _GEN_2518;
        end else begin
          dirty_1_75 <= _GEN_13053;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_76 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_76 <= _GEN_2519;
        end else begin
          dirty_1_76 <= _GEN_13054;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_77 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_77 <= _GEN_2520;
        end else begin
          dirty_1_77 <= _GEN_13055;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_78 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_78 <= _GEN_2521;
        end else begin
          dirty_1_78 <= _GEN_13056;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_79 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_79 <= _GEN_2522;
        end else begin
          dirty_1_79 <= _GEN_13057;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_80 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_80 <= _GEN_2523;
        end else begin
          dirty_1_80 <= _GEN_13058;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_81 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_81 <= _GEN_2524;
        end else begin
          dirty_1_81 <= _GEN_13059;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_82 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_82 <= _GEN_2525;
        end else begin
          dirty_1_82 <= _GEN_13060;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_83 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_83 <= _GEN_2526;
        end else begin
          dirty_1_83 <= _GEN_13061;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_84 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_84 <= _GEN_2527;
        end else begin
          dirty_1_84 <= _GEN_13062;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_85 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_85 <= _GEN_2528;
        end else begin
          dirty_1_85 <= _GEN_13063;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_86 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_86 <= _GEN_2529;
        end else begin
          dirty_1_86 <= _GEN_13064;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_87 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_87 <= _GEN_2530;
        end else begin
          dirty_1_87 <= _GEN_13065;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_88 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_88 <= _GEN_2531;
        end else begin
          dirty_1_88 <= _GEN_13066;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_89 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_89 <= _GEN_2532;
        end else begin
          dirty_1_89 <= _GEN_13067;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_90 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_90 <= _GEN_2533;
        end else begin
          dirty_1_90 <= _GEN_13068;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_91 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_91 <= _GEN_2534;
        end else begin
          dirty_1_91 <= _GEN_13069;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_92 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_92 <= _GEN_2535;
        end else begin
          dirty_1_92 <= _GEN_13070;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_93 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_93 <= _GEN_2536;
        end else begin
          dirty_1_93 <= _GEN_13071;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_94 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_94 <= _GEN_2537;
        end else begin
          dirty_1_94 <= _GEN_13072;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_95 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_95 <= _GEN_2538;
        end else begin
          dirty_1_95 <= _GEN_13073;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_96 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_96 <= _GEN_2539;
        end else begin
          dirty_1_96 <= _GEN_13074;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_97 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_97 <= _GEN_2540;
        end else begin
          dirty_1_97 <= _GEN_13075;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_98 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_98 <= _GEN_2541;
        end else begin
          dirty_1_98 <= _GEN_13076;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_99 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_99 <= _GEN_2542;
        end else begin
          dirty_1_99 <= _GEN_13077;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_100 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_100 <= _GEN_2543;
        end else begin
          dirty_1_100 <= _GEN_13078;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_101 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_101 <= _GEN_2544;
        end else begin
          dirty_1_101 <= _GEN_13079;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_102 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_102 <= _GEN_2545;
        end else begin
          dirty_1_102 <= _GEN_13080;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_103 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_103 <= _GEN_2546;
        end else begin
          dirty_1_103 <= _GEN_13081;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_104 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_104 <= _GEN_2547;
        end else begin
          dirty_1_104 <= _GEN_13082;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_105 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_105 <= _GEN_2548;
        end else begin
          dirty_1_105 <= _GEN_13083;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_106 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_106 <= _GEN_2549;
        end else begin
          dirty_1_106 <= _GEN_13084;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_107 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_107 <= _GEN_2550;
        end else begin
          dirty_1_107 <= _GEN_13085;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_108 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_108 <= _GEN_2551;
        end else begin
          dirty_1_108 <= _GEN_13086;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_109 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_109 <= _GEN_2552;
        end else begin
          dirty_1_109 <= _GEN_13087;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_110 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_110 <= _GEN_2553;
        end else begin
          dirty_1_110 <= _GEN_13088;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_111 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_111 <= _GEN_2554;
        end else begin
          dirty_1_111 <= _GEN_13089;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_112 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_112 <= _GEN_2555;
        end else begin
          dirty_1_112 <= _GEN_13090;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_113 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_113 <= _GEN_2556;
        end else begin
          dirty_1_113 <= _GEN_13091;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_114 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_114 <= _GEN_2557;
        end else begin
          dirty_1_114 <= _GEN_13092;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_115 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_115 <= _GEN_2558;
        end else begin
          dirty_1_115 <= _GEN_13093;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_116 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_116 <= _GEN_2559;
        end else begin
          dirty_1_116 <= _GEN_13094;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_117 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_117 <= _GEN_2560;
        end else begin
          dirty_1_117 <= _GEN_13095;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_118 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_118 <= _GEN_2561;
        end else begin
          dirty_1_118 <= _GEN_13096;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_119 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_119 <= _GEN_2562;
        end else begin
          dirty_1_119 <= _GEN_13097;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_120 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_120 <= _GEN_2563;
        end else begin
          dirty_1_120 <= _GEN_13098;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_121 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_121 <= _GEN_2564;
        end else begin
          dirty_1_121 <= _GEN_13099;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_122 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_122 <= _GEN_2565;
        end else begin
          dirty_1_122 <= _GEN_13100;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_123 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_123 <= _GEN_2566;
        end else begin
          dirty_1_123 <= _GEN_13101;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_124 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_124 <= _GEN_2567;
        end else begin
          dirty_1_124 <= _GEN_13102;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_125 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_125 <= _GEN_2568;
        end else begin
          dirty_1_125 <= _GEN_13103;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_126 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_126 <= _GEN_2569;
        end else begin
          dirty_1_126 <= _GEN_13104;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      dirty_1_127 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (3'h2 == state) begin // @[d_cache.scala 78:18]
          dirty_1_127 <= _GEN_2570;
        end else begin
          dirty_1_127 <= _GEN_13105;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:27]
      way0_hit <= 1'h0; // @[d_cache.scala 26:27]
    end else begin
      way0_hit <= _T_6;
    end
    if (reset) begin // @[d_cache.scala 27:27]
      way1_hit <= 1'h0; // @[d_cache.scala 27:27]
    end else begin
      way1_hit <= _T_11;
    end
    if (reset) begin // @[d_cache.scala 29:34]
      write_back_data <= 64'h0; // @[d_cache.scala 29:34]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          write_back_data <= _GEN_12848;
        end
      end
    end
    write_back_addr <= _GEN_17833[31:0]; // @[d_cache.scala 30:{34,34}]
    if (reset) begin // @[d_cache.scala 33:28]
      unuse_way <= 2'h0; // @[d_cache.scala 33:28]
    end else if (~_GEN_255) begin // @[d_cache.scala 65:31]
      unuse_way <= 2'h1; // @[d_cache.scala 66:19]
    end else if (~_GEN_512) begin // @[d_cache.scala 67:37]
      unuse_way <= 2'h2; // @[d_cache.scala 68:19]
    end else begin
      unuse_way <= 2'h0; // @[d_cache.scala 70:19]
    end
    if (reset) begin // @[d_cache.scala 34:31]
      receive_data <= 64'h0; // @[d_cache.scala 34:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          receive_data <= _GEN_12078;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:24]
      quene <= 1'h0; // @[d_cache.scala 35:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 78:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 78:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 78:18]
          quene <= _GEN_12463;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 73:24]
      state <= 3'h0; // @[d_cache.scala 73:24]
    end else if (3'h0 == state) begin // @[d_cache.scala 78:18]
      if (io_from_lsu_arvalid) begin // @[d_cache.scala 80:38]
        state <= 3'h1; // @[d_cache.scala 81:23]
      end else if (io_from_lsu_awvalid) begin // @[d_cache.scala 82:44]
        state <= 3'h2; // @[d_cache.scala 83:23]
      end
    end else if (3'h1 == state) begin // @[d_cache.scala 78:18]
      if (way0_hit) begin // @[d_cache.scala 88:27]
        state <= _GEN_902;
      end else begin
        state <= _GEN_1031;
      end
    end else if (3'h2 == state) begin // @[d_cache.scala 78:18]
      state <= _GEN_2058;
    end else begin
      state <= _GEN_12077;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"read addr : %x  write addr : %x\n",io_from_lsu_araddr,io_from_lsu_awaddr); // @[d_cache.scala 15:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"d_cache state:%d\n",state); // @[d_cache.scala 74:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"bvalid:%d\n",io_from_axi_bvalid); // @[d_cache.scala 75:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"receive data:%x\n",receive_data); // @[d_cache.scala 76:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"wstrb:%x\n",io_from_lsu_wstrb); // @[d_cache.scala 77:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_24 & _T_25 & way0_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_0:%d\n",7'h7f == index[6:0] ? dirty_0_127 : _GEN_900); // @[d_cache.scala 90:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17835 & ~way0_hit & way1_hit & io_from_lsu_rready & _T_1) begin
          $fwrite(32'h80000002,"dirty_1:%d\n",7'h7f == index[6:0] ? dirty_1_127 : _GEN_1029); // @[d_cache.scala 96:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"to lsu rdata:%x\n",io_to_lsu_rdata); // @[d_cache.scala 356:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"cacheline0:%x   cacheline1:%x\n",_GEN_1160,_GEN_5393); // @[d_cache.scala 357:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  ram_0_64 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  ram_0_65 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  ram_0_66 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  ram_0_67 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  ram_0_68 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  ram_0_69 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  ram_0_70 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  ram_0_71 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  ram_0_72 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  ram_0_73 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  ram_0_74 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  ram_0_75 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  ram_0_76 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  ram_0_77 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  ram_0_78 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  ram_0_79 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  ram_0_80 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  ram_0_81 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  ram_0_82 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  ram_0_83 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  ram_0_84 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  ram_0_85 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  ram_0_86 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  ram_0_87 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  ram_0_88 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  ram_0_89 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  ram_0_90 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  ram_0_91 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  ram_0_92 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  ram_0_93 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  ram_0_94 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  ram_0_95 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  ram_0_96 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  ram_0_97 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  ram_0_98 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  ram_0_99 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  ram_0_100 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  ram_0_101 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  ram_0_102 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  ram_0_103 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  ram_0_104 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  ram_0_105 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  ram_0_106 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  ram_0_107 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  ram_0_108 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  ram_0_109 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  ram_0_110 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  ram_0_111 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  ram_0_112 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  ram_0_113 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  ram_0_114 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  ram_0_115 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  ram_0_116 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  ram_0_117 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  ram_0_118 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  ram_0_119 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  ram_0_120 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  ram_0_121 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  ram_0_122 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  ram_0_123 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  ram_0_124 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  ram_0_125 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  ram_0_126 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  ram_0_127 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  ram_1_0 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  ram_1_1 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  ram_1_2 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  ram_1_3 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  ram_1_4 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  ram_1_5 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  ram_1_6 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  ram_1_7 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  ram_1_8 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  ram_1_9 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  ram_1_10 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  ram_1_11 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  ram_1_12 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  ram_1_13 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  ram_1_14 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  ram_1_15 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  ram_1_16 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  ram_1_17 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  ram_1_18 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  ram_1_19 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  ram_1_20 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  ram_1_21 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  ram_1_22 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  ram_1_23 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  ram_1_24 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  ram_1_25 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  ram_1_26 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  ram_1_27 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  ram_1_28 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  ram_1_29 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  ram_1_30 = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  ram_1_31 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  ram_1_32 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  ram_1_33 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  ram_1_34 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  ram_1_35 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  ram_1_36 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  ram_1_37 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  ram_1_38 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  ram_1_39 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  ram_1_40 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  ram_1_41 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  ram_1_42 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  ram_1_43 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  ram_1_44 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  ram_1_45 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  ram_1_46 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  ram_1_47 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  ram_1_48 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  ram_1_49 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  ram_1_50 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  ram_1_51 = _RAND_179[63:0];
  _RAND_180 = {2{`RANDOM}};
  ram_1_52 = _RAND_180[63:0];
  _RAND_181 = {2{`RANDOM}};
  ram_1_53 = _RAND_181[63:0];
  _RAND_182 = {2{`RANDOM}};
  ram_1_54 = _RAND_182[63:0];
  _RAND_183 = {2{`RANDOM}};
  ram_1_55 = _RAND_183[63:0];
  _RAND_184 = {2{`RANDOM}};
  ram_1_56 = _RAND_184[63:0];
  _RAND_185 = {2{`RANDOM}};
  ram_1_57 = _RAND_185[63:0];
  _RAND_186 = {2{`RANDOM}};
  ram_1_58 = _RAND_186[63:0];
  _RAND_187 = {2{`RANDOM}};
  ram_1_59 = _RAND_187[63:0];
  _RAND_188 = {2{`RANDOM}};
  ram_1_60 = _RAND_188[63:0];
  _RAND_189 = {2{`RANDOM}};
  ram_1_61 = _RAND_189[63:0];
  _RAND_190 = {2{`RANDOM}};
  ram_1_62 = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  ram_1_63 = _RAND_191[63:0];
  _RAND_192 = {2{`RANDOM}};
  ram_1_64 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  ram_1_65 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  ram_1_66 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  ram_1_67 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  ram_1_68 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  ram_1_69 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  ram_1_70 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  ram_1_71 = _RAND_199[63:0];
  _RAND_200 = {2{`RANDOM}};
  ram_1_72 = _RAND_200[63:0];
  _RAND_201 = {2{`RANDOM}};
  ram_1_73 = _RAND_201[63:0];
  _RAND_202 = {2{`RANDOM}};
  ram_1_74 = _RAND_202[63:0];
  _RAND_203 = {2{`RANDOM}};
  ram_1_75 = _RAND_203[63:0];
  _RAND_204 = {2{`RANDOM}};
  ram_1_76 = _RAND_204[63:0];
  _RAND_205 = {2{`RANDOM}};
  ram_1_77 = _RAND_205[63:0];
  _RAND_206 = {2{`RANDOM}};
  ram_1_78 = _RAND_206[63:0];
  _RAND_207 = {2{`RANDOM}};
  ram_1_79 = _RAND_207[63:0];
  _RAND_208 = {2{`RANDOM}};
  ram_1_80 = _RAND_208[63:0];
  _RAND_209 = {2{`RANDOM}};
  ram_1_81 = _RAND_209[63:0];
  _RAND_210 = {2{`RANDOM}};
  ram_1_82 = _RAND_210[63:0];
  _RAND_211 = {2{`RANDOM}};
  ram_1_83 = _RAND_211[63:0];
  _RAND_212 = {2{`RANDOM}};
  ram_1_84 = _RAND_212[63:0];
  _RAND_213 = {2{`RANDOM}};
  ram_1_85 = _RAND_213[63:0];
  _RAND_214 = {2{`RANDOM}};
  ram_1_86 = _RAND_214[63:0];
  _RAND_215 = {2{`RANDOM}};
  ram_1_87 = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  ram_1_88 = _RAND_216[63:0];
  _RAND_217 = {2{`RANDOM}};
  ram_1_89 = _RAND_217[63:0];
  _RAND_218 = {2{`RANDOM}};
  ram_1_90 = _RAND_218[63:0];
  _RAND_219 = {2{`RANDOM}};
  ram_1_91 = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  ram_1_92 = _RAND_220[63:0];
  _RAND_221 = {2{`RANDOM}};
  ram_1_93 = _RAND_221[63:0];
  _RAND_222 = {2{`RANDOM}};
  ram_1_94 = _RAND_222[63:0];
  _RAND_223 = {2{`RANDOM}};
  ram_1_95 = _RAND_223[63:0];
  _RAND_224 = {2{`RANDOM}};
  ram_1_96 = _RAND_224[63:0];
  _RAND_225 = {2{`RANDOM}};
  ram_1_97 = _RAND_225[63:0];
  _RAND_226 = {2{`RANDOM}};
  ram_1_98 = _RAND_226[63:0];
  _RAND_227 = {2{`RANDOM}};
  ram_1_99 = _RAND_227[63:0];
  _RAND_228 = {2{`RANDOM}};
  ram_1_100 = _RAND_228[63:0];
  _RAND_229 = {2{`RANDOM}};
  ram_1_101 = _RAND_229[63:0];
  _RAND_230 = {2{`RANDOM}};
  ram_1_102 = _RAND_230[63:0];
  _RAND_231 = {2{`RANDOM}};
  ram_1_103 = _RAND_231[63:0];
  _RAND_232 = {2{`RANDOM}};
  ram_1_104 = _RAND_232[63:0];
  _RAND_233 = {2{`RANDOM}};
  ram_1_105 = _RAND_233[63:0];
  _RAND_234 = {2{`RANDOM}};
  ram_1_106 = _RAND_234[63:0];
  _RAND_235 = {2{`RANDOM}};
  ram_1_107 = _RAND_235[63:0];
  _RAND_236 = {2{`RANDOM}};
  ram_1_108 = _RAND_236[63:0];
  _RAND_237 = {2{`RANDOM}};
  ram_1_109 = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  ram_1_110 = _RAND_238[63:0];
  _RAND_239 = {2{`RANDOM}};
  ram_1_111 = _RAND_239[63:0];
  _RAND_240 = {2{`RANDOM}};
  ram_1_112 = _RAND_240[63:0];
  _RAND_241 = {2{`RANDOM}};
  ram_1_113 = _RAND_241[63:0];
  _RAND_242 = {2{`RANDOM}};
  ram_1_114 = _RAND_242[63:0];
  _RAND_243 = {2{`RANDOM}};
  ram_1_115 = _RAND_243[63:0];
  _RAND_244 = {2{`RANDOM}};
  ram_1_116 = _RAND_244[63:0];
  _RAND_245 = {2{`RANDOM}};
  ram_1_117 = _RAND_245[63:0];
  _RAND_246 = {2{`RANDOM}};
  ram_1_118 = _RAND_246[63:0];
  _RAND_247 = {2{`RANDOM}};
  ram_1_119 = _RAND_247[63:0];
  _RAND_248 = {2{`RANDOM}};
  ram_1_120 = _RAND_248[63:0];
  _RAND_249 = {2{`RANDOM}};
  ram_1_121 = _RAND_249[63:0];
  _RAND_250 = {2{`RANDOM}};
  ram_1_122 = _RAND_250[63:0];
  _RAND_251 = {2{`RANDOM}};
  ram_1_123 = _RAND_251[63:0];
  _RAND_252 = {2{`RANDOM}};
  ram_1_124 = _RAND_252[63:0];
  _RAND_253 = {2{`RANDOM}};
  ram_1_125 = _RAND_253[63:0];
  _RAND_254 = {2{`RANDOM}};
  ram_1_126 = _RAND_254[63:0];
  _RAND_255 = {2{`RANDOM}};
  ram_1_127 = _RAND_255[63:0];
  _RAND_256 = {1{`RANDOM}};
  tag_0_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  tag_0_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  tag_0_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  tag_0_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  tag_0_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  tag_0_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  tag_0_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  tag_0_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  tag_0_8 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  tag_0_9 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  tag_0_10 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  tag_0_11 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  tag_0_12 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  tag_0_13 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  tag_0_14 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  tag_0_15 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  tag_0_16 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  tag_0_17 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  tag_0_18 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  tag_0_19 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  tag_0_20 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  tag_0_21 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  tag_0_22 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  tag_0_23 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  tag_0_24 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  tag_0_25 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  tag_0_26 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  tag_0_27 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  tag_0_28 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  tag_0_29 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  tag_0_30 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  tag_0_31 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  tag_0_32 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  tag_0_33 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  tag_0_34 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  tag_0_35 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  tag_0_36 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  tag_0_37 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  tag_0_38 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  tag_0_39 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  tag_0_40 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  tag_0_41 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  tag_0_42 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  tag_0_43 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  tag_0_44 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  tag_0_45 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  tag_0_46 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  tag_0_47 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  tag_0_48 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  tag_0_49 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  tag_0_50 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  tag_0_51 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  tag_0_52 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  tag_0_53 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  tag_0_54 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  tag_0_55 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  tag_0_56 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  tag_0_57 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  tag_0_58 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  tag_0_59 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  tag_0_60 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  tag_0_61 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  tag_0_62 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  tag_0_63 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  tag_0_64 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  tag_0_65 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  tag_0_66 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  tag_0_67 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  tag_0_68 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  tag_0_69 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  tag_0_70 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  tag_0_71 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  tag_0_72 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  tag_0_73 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  tag_0_74 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  tag_0_75 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  tag_0_76 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  tag_0_77 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  tag_0_78 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  tag_0_79 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  tag_0_80 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  tag_0_81 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  tag_0_82 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  tag_0_83 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  tag_0_84 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  tag_0_85 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  tag_0_86 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  tag_0_87 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  tag_0_88 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  tag_0_89 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  tag_0_90 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  tag_0_91 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  tag_0_92 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  tag_0_93 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  tag_0_94 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  tag_0_95 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  tag_0_96 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  tag_0_97 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  tag_0_98 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  tag_0_99 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  tag_0_100 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  tag_0_101 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  tag_0_102 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  tag_0_103 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  tag_0_104 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  tag_0_105 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  tag_0_106 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  tag_0_107 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  tag_0_108 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  tag_0_109 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  tag_0_110 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  tag_0_111 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  tag_0_112 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  tag_0_113 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  tag_0_114 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  tag_0_115 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  tag_0_116 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  tag_0_117 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  tag_0_118 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  tag_0_119 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  tag_0_120 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  tag_0_121 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  tag_0_122 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  tag_0_123 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  tag_0_124 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  tag_0_125 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  tag_0_126 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  tag_0_127 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  tag_1_0 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  tag_1_1 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  tag_1_2 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  tag_1_3 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  tag_1_4 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  tag_1_5 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  tag_1_6 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  tag_1_7 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  tag_1_8 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  tag_1_9 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  tag_1_10 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  tag_1_11 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  tag_1_12 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  tag_1_13 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  tag_1_14 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  tag_1_15 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  tag_1_16 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  tag_1_17 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  tag_1_18 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  tag_1_19 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  tag_1_20 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  tag_1_21 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  tag_1_22 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  tag_1_23 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  tag_1_24 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  tag_1_25 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  tag_1_26 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  tag_1_27 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  tag_1_28 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  tag_1_29 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  tag_1_30 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  tag_1_31 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  tag_1_32 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  tag_1_33 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  tag_1_34 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  tag_1_35 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  tag_1_36 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  tag_1_37 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  tag_1_38 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  tag_1_39 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  tag_1_40 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  tag_1_41 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  tag_1_42 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  tag_1_43 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  tag_1_44 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  tag_1_45 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  tag_1_46 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  tag_1_47 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  tag_1_48 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  tag_1_49 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  tag_1_50 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  tag_1_51 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  tag_1_52 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  tag_1_53 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  tag_1_54 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  tag_1_55 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  tag_1_56 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  tag_1_57 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  tag_1_58 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  tag_1_59 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  tag_1_60 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  tag_1_61 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  tag_1_62 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  tag_1_63 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  tag_1_64 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  tag_1_65 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  tag_1_66 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  tag_1_67 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  tag_1_68 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  tag_1_69 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  tag_1_70 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  tag_1_71 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  tag_1_72 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  tag_1_73 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  tag_1_74 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  tag_1_75 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  tag_1_76 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  tag_1_77 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  tag_1_78 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  tag_1_79 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  tag_1_80 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  tag_1_81 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  tag_1_82 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  tag_1_83 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  tag_1_84 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  tag_1_85 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  tag_1_86 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  tag_1_87 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  tag_1_88 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  tag_1_89 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  tag_1_90 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  tag_1_91 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  tag_1_92 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  tag_1_93 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  tag_1_94 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  tag_1_95 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  tag_1_96 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  tag_1_97 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  tag_1_98 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  tag_1_99 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  tag_1_100 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  tag_1_101 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  tag_1_102 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  tag_1_103 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  tag_1_104 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  tag_1_105 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  tag_1_106 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  tag_1_107 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  tag_1_108 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  tag_1_109 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  tag_1_110 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  tag_1_111 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  tag_1_112 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  tag_1_113 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  tag_1_114 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  tag_1_115 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  tag_1_116 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  tag_1_117 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  tag_1_118 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  tag_1_119 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  tag_1_120 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  tag_1_121 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  tag_1_122 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  tag_1_123 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  tag_1_124 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  tag_1_125 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  tag_1_126 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  tag_1_127 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  valid_0_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_0_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_0_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_0_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_0_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_0_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_0_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_0_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_0_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_0_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_0_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_0_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_0_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_0_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_0_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_0_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  valid_0_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  valid_0_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  valid_0_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  valid_0_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  valid_0_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  valid_0_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  valid_0_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  valid_0_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  valid_0_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  valid_0_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  valid_0_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  valid_0_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  valid_0_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  valid_0_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  valid_0_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  valid_0_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  valid_0_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  valid_0_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  valid_0_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  valid_0_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  valid_0_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  valid_0_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  valid_0_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  valid_0_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  valid_0_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  valid_0_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  valid_0_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  valid_0_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  valid_0_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  valid_0_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  valid_0_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  valid_0_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  valid_0_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  valid_0_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  valid_0_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  valid_0_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  valid_0_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  valid_0_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  valid_0_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  valid_0_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  valid_0_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  valid_0_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  valid_0_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  valid_0_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  valid_0_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  valid_0_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  valid_0_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  valid_0_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  valid_0_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_0_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_0_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_0_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_0_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_0_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_0_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_0_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_0_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_0_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_0_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_0_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_0_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_0_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_0_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_0_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_0_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_0_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_0_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_0_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_0_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_0_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_0_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_0_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_0_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_0_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_0_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_0_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_0_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_0_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_0_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_0_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_0_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_0_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_0_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_0_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_0_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_0_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_0_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_0_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_0_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_0_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_0_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_0_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_0_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_0_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_0_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_0_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_0_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_0_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_0_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_0_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_0_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_0_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_0_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_0_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_0_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_0_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_0_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_0_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_0_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_0_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_0_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_0_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  valid_1_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  valid_1_1 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  valid_1_2 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  valid_1_3 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  valid_1_4 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  valid_1_5 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  valid_1_6 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  valid_1_7 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  valid_1_8 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  valid_1_9 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  valid_1_10 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  valid_1_11 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  valid_1_12 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  valid_1_13 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  valid_1_14 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  valid_1_15 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  valid_1_16 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  valid_1_17 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  valid_1_18 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  valid_1_19 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  valid_1_20 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  valid_1_21 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  valid_1_22 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  valid_1_23 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  valid_1_24 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  valid_1_25 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  valid_1_26 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  valid_1_27 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  valid_1_28 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  valid_1_29 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  valid_1_30 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  valid_1_31 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  valid_1_32 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  valid_1_33 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  valid_1_34 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  valid_1_35 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  valid_1_36 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  valid_1_37 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  valid_1_38 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  valid_1_39 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  valid_1_40 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  valid_1_41 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  valid_1_42 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  valid_1_43 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  valid_1_44 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  valid_1_45 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  valid_1_46 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  valid_1_47 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  valid_1_48 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  valid_1_49 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  valid_1_50 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  valid_1_51 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  valid_1_52 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  valid_1_53 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  valid_1_54 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  valid_1_55 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  valid_1_56 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  valid_1_57 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  valid_1_58 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  valid_1_59 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  valid_1_60 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  valid_1_61 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  valid_1_62 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  valid_1_63 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  valid_1_64 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  valid_1_65 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  valid_1_66 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  valid_1_67 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  valid_1_68 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  valid_1_69 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  valid_1_70 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  valid_1_71 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  valid_1_72 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  valid_1_73 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  valid_1_74 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  valid_1_75 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  valid_1_76 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  valid_1_77 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  valid_1_78 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  valid_1_79 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  valid_1_80 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  valid_1_81 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  valid_1_82 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  valid_1_83 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  valid_1_84 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  valid_1_85 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  valid_1_86 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  valid_1_87 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  valid_1_88 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  valid_1_89 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  valid_1_90 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  valid_1_91 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  valid_1_92 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  valid_1_93 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  valid_1_94 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  valid_1_95 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  valid_1_96 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  valid_1_97 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  valid_1_98 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  valid_1_99 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  valid_1_100 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  valid_1_101 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  valid_1_102 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  valid_1_103 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  valid_1_104 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  valid_1_105 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  valid_1_106 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  valid_1_107 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  valid_1_108 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  valid_1_109 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  valid_1_110 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  valid_1_111 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  valid_1_112 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  valid_1_113 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  valid_1_114 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  valid_1_115 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  valid_1_116 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  valid_1_117 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  valid_1_118 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  valid_1_119 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  valid_1_120 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  valid_1_121 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  valid_1_122 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  valid_1_123 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  valid_1_124 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  valid_1_125 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  valid_1_126 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  valid_1_127 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  dirty_0_0 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  dirty_0_1 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  dirty_0_2 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  dirty_0_3 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  dirty_0_4 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  dirty_0_5 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  dirty_0_6 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  dirty_0_7 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  dirty_0_8 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  dirty_0_9 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  dirty_0_10 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  dirty_0_11 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  dirty_0_12 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  dirty_0_13 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  dirty_0_14 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  dirty_0_15 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  dirty_0_16 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  dirty_0_17 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  dirty_0_18 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  dirty_0_19 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  dirty_0_20 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  dirty_0_21 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  dirty_0_22 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  dirty_0_23 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  dirty_0_24 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  dirty_0_25 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  dirty_0_26 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  dirty_0_27 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  dirty_0_28 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  dirty_0_29 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  dirty_0_30 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  dirty_0_31 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  dirty_0_32 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  dirty_0_33 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  dirty_0_34 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  dirty_0_35 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  dirty_0_36 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  dirty_0_37 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  dirty_0_38 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  dirty_0_39 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  dirty_0_40 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  dirty_0_41 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  dirty_0_42 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  dirty_0_43 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  dirty_0_44 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  dirty_0_45 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  dirty_0_46 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  dirty_0_47 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  dirty_0_48 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  dirty_0_49 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  dirty_0_50 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  dirty_0_51 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  dirty_0_52 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  dirty_0_53 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  dirty_0_54 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  dirty_0_55 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  dirty_0_56 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  dirty_0_57 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  dirty_0_58 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  dirty_0_59 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  dirty_0_60 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  dirty_0_61 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  dirty_0_62 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  dirty_0_63 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  dirty_0_64 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  dirty_0_65 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  dirty_0_66 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  dirty_0_67 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  dirty_0_68 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  dirty_0_69 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  dirty_0_70 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  dirty_0_71 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  dirty_0_72 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  dirty_0_73 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  dirty_0_74 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  dirty_0_75 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  dirty_0_76 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  dirty_0_77 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  dirty_0_78 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  dirty_0_79 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  dirty_0_80 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  dirty_0_81 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  dirty_0_82 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  dirty_0_83 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  dirty_0_84 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  dirty_0_85 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  dirty_0_86 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  dirty_0_87 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  dirty_0_88 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  dirty_0_89 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  dirty_0_90 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  dirty_0_91 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  dirty_0_92 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  dirty_0_93 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  dirty_0_94 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  dirty_0_95 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  dirty_0_96 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  dirty_0_97 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  dirty_0_98 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  dirty_0_99 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  dirty_0_100 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  dirty_0_101 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  dirty_0_102 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  dirty_0_103 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  dirty_0_104 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  dirty_0_105 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  dirty_0_106 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  dirty_0_107 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  dirty_0_108 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  dirty_0_109 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  dirty_0_110 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  dirty_0_111 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  dirty_0_112 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  dirty_0_113 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  dirty_0_114 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  dirty_0_115 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  dirty_0_116 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  dirty_0_117 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  dirty_0_118 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  dirty_0_119 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  dirty_0_120 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  dirty_0_121 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  dirty_0_122 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  dirty_0_123 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  dirty_0_124 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  dirty_0_125 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  dirty_0_126 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  dirty_0_127 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  dirty_1_0 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  dirty_1_1 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  dirty_1_2 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  dirty_1_3 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  dirty_1_4 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  dirty_1_5 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  dirty_1_6 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  dirty_1_7 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  dirty_1_8 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  dirty_1_9 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  dirty_1_10 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  dirty_1_11 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  dirty_1_12 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  dirty_1_13 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  dirty_1_14 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  dirty_1_15 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  dirty_1_16 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  dirty_1_17 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  dirty_1_18 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  dirty_1_19 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  dirty_1_20 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  dirty_1_21 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  dirty_1_22 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  dirty_1_23 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  dirty_1_24 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  dirty_1_25 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  dirty_1_26 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  dirty_1_27 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  dirty_1_28 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  dirty_1_29 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  dirty_1_30 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  dirty_1_31 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  dirty_1_32 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  dirty_1_33 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  dirty_1_34 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  dirty_1_35 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  dirty_1_36 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  dirty_1_37 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  dirty_1_38 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  dirty_1_39 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  dirty_1_40 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  dirty_1_41 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  dirty_1_42 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  dirty_1_43 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  dirty_1_44 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  dirty_1_45 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  dirty_1_46 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  dirty_1_47 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  dirty_1_48 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  dirty_1_49 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  dirty_1_50 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  dirty_1_51 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  dirty_1_52 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  dirty_1_53 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  dirty_1_54 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  dirty_1_55 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  dirty_1_56 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  dirty_1_57 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  dirty_1_58 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  dirty_1_59 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  dirty_1_60 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  dirty_1_61 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  dirty_1_62 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  dirty_1_63 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  dirty_1_64 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  dirty_1_65 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  dirty_1_66 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  dirty_1_67 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  dirty_1_68 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  dirty_1_69 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  dirty_1_70 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  dirty_1_71 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  dirty_1_72 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  dirty_1_73 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  dirty_1_74 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  dirty_1_75 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  dirty_1_76 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  dirty_1_77 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  dirty_1_78 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  dirty_1_79 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  dirty_1_80 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  dirty_1_81 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  dirty_1_82 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  dirty_1_83 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  dirty_1_84 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  dirty_1_85 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  dirty_1_86 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  dirty_1_87 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  dirty_1_88 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  dirty_1_89 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  dirty_1_90 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  dirty_1_91 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  dirty_1_92 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  dirty_1_93 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  dirty_1_94 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  dirty_1_95 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  dirty_1_96 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  dirty_1_97 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  dirty_1_98 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  dirty_1_99 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  dirty_1_100 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  dirty_1_101 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  dirty_1_102 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  dirty_1_103 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  dirty_1_104 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  dirty_1_105 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  dirty_1_106 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  dirty_1_107 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  dirty_1_108 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  dirty_1_109 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  dirty_1_110 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  dirty_1_111 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  dirty_1_112 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  dirty_1_113 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  dirty_1_114 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  dirty_1_115 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  dirty_1_116 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  dirty_1_117 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  dirty_1_118 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  dirty_1_119 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  dirty_1_120 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  dirty_1_121 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  dirty_1_122 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  dirty_1_123 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  dirty_1_124 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  dirty_1_125 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  dirty_1_126 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  dirty_1_127 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  way0_hit = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  way1_hit = _RAND_1025[0:0];
  _RAND_1026 = {2{`RANDOM}};
  write_back_data = _RAND_1026[63:0];
  _RAND_1027 = {1{`RANDOM}};
  write_back_addr = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  unuse_way = _RAND_1028[1:0];
  _RAND_1029 = {2{`RANDOM}};
  receive_data = _RAND_1029[63:0];
  _RAND_1030 = {1{`RANDOM}};
  quene = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  state = _RAND_1031[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
