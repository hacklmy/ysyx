/* verilator lint_off WIDTH */
module ALU(
  input  [63:0] io_src1_value,
  input  [63:0] io_src2_value,
  input  [31:0] io_ALUop,
  output [63:0] io_alu_res
);
  wire [63:0] add_res = io_src1_value + io_src2_value; // @[ALU.scala 25:30]
  wire [63:0] sub_res = io_src1_value - io_src2_value; // @[ALU.scala 26:30]
  wire [63:0] sra_res = $signed(io_src1_value) >>> io_src2_value[5:0]; // @[ALU.scala 27:60]
  wire [63:0] srl_res = io_src1_value >> io_src2_value[5:0]; // @[ALU.scala 28:30]
  wire [126:0] _GEN_0 = {{63'd0}, io_src1_value}; // @[ALU.scala 29:30]
  wire [126:0] sll_res = _GEN_0 << io_src2_value[5:0]; // @[ALU.scala 29:30]
  wire [31:0] _sraw_res_T_1 = io_src1_value[31:0]; // @[ALU.scala 30:43]
  wire [31:0] sraw_res = $signed(_sraw_res_T_1) >>> io_src2_value[4:0]; // @[ALU.scala 30:46]
  wire [31:0] srlw_res = io_src1_value[31:0] >> io_src2_value[4:0]; // @[ALU.scala 31:37]
  wire [62:0] _GEN_1 = {{31'd0}, io_src1_value[31:0]}; // @[ALU.scala 32:37]
  wire [62:0] sllw_res = _GEN_1 << io_src2_value[4:0]; // @[ALU.scala 32:37]
  wire [63:0] or_res = io_src1_value | io_src2_value; // @[ALU.scala 33:29]
  wire [63:0] xor_res = io_src1_value ^ io_src2_value; // @[ALU.scala 34:30]
  wire [63:0] and_res = io_src1_value & io_src2_value; // @[ALU.scala 35:30]
  wire [127:0] _mlu_res_T = io_src1_value * io_src2_value; // @[ALU.scala 36:31]
  wire [63:0] mlu_res = _mlu_res_T[63:0]; // @[ALU.scala 36:44]
  wire [63:0] _mluw_res_T_2 = io_src1_value[31:0] * io_src2_value[31:0]; // @[ALU.scala 37:38]
  wire [31:0] mluw_res = _mluw_res_T_2[31:0]; // @[ALU.scala 37:57]
  wire [31:0] _divw_res_T_3 = io_src2_value[31:0]; // @[ALU.scala 38:64]
  wire [32:0] _divw_res_T_4 = $signed(_sraw_res_T_1) / $signed(_divw_res_T_3); // @[ALU.scala 38:45]
  wire [31:0] divw_res = _divw_res_T_4[31:0]; // @[ALU.scala 38:71]
  wire [31:0] divuw_res = io_src1_value[31:0] / io_src2_value[31:0]; // @[ALU.scala 39:39]
  wire [31:0] remw_res = $signed(_sraw_res_T_1) % $signed(_divw_res_T_3); // @[ALU.scala 40:71]
  wire [31:0] remuw_res = io_src1_value[31:0] % io_src2_value[31:0]; // @[ALU.scala 41:39]
  wire [64:0] div_res = $signed(io_src1_value) / $signed(io_src2_value); // @[ALU.scala 42:59]
  wire [63:0] divu_res = io_src1_value / io_src2_value; // @[ALU.scala 43:31]
  wire [63:0] rem_res = $signed(io_src1_value) % $signed(io_src2_value); // @[ALU.scala 44:59]
  wire [63:0] remu_res = io_src1_value % io_src2_value; // @[ALU.scala 45:31]
  wire [63:0] _alu_res_T_1 = io_src1_value + 64'h4; // @[ALU.scala 62:29]
  wire  _alu_res_T_4 = io_src1_value < io_src2_value; // @[ALU.scala 65:33]
  wire  _alu_res_T_8 = $signed(io_src1_value) < $signed(io_src2_value); // @[ALU.scala 67:41]
  wire [31:0] _alu_res_T_12 = add_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_14 = {_alu_res_T_12,add_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_17 = sub_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_19 = {_alu_res_T_17,sub_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_22 = sllw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_24 = {_alu_res_T_22,sllw_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_27 = sraw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _alu_res_T_28 = $signed(_sraw_res_T_1) >>> io_src2_value[4:0]; // @[ALU.scala 86:55]
  wire [63:0] _alu_res_T_29 = {_alu_res_T_27,_alu_res_T_28}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_32 = srlw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_34 = {_alu_res_T_32,srlw_res}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_37 = mluw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_38 = {_alu_res_T_37,mluw_res}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_41 = divw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_42 = {_alu_res_T_41,divw_res}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_45 = divuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_46 = {_alu_res_T_45,divuw_res}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_49 = remw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_50 = {_alu_res_T_49,remw_res}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_53 = remuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_54 = {_alu_res_T_53,remuw_res}; // @[Cat.scala 31:58]
  wire [63:0] _alu_res_T_56 = 32'hf == io_ALUop ? add_res : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_58 = 32'h4 == io_ALUop ? io_src2_value : _alu_res_T_56; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_60 = 32'h5 == io_ALUop ? _alu_res_T_1 : _alu_res_T_58; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_62 = 32'h6 == io_ALUop ? _alu_res_T_1 : _alu_res_T_60; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_64 = 32'h1e == io_ALUop ? {{63'd0}, _alu_res_T_4} : _alu_res_T_62; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_66 = 32'h1f == io_ALUop ? {{63'd0}, _alu_res_T_8} : _alu_res_T_64; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_68 = 32'hc == io_ALUop ? _alu_res_T_14 : _alu_res_T_66; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_70 = 32'he == io_ALUop ? sub_res : _alu_res_T_68; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_72 = 32'h15 == io_ALUop ? sra_res : _alu_res_T_70; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_74 = 32'hb == io_ALUop ? or_res : _alu_res_T_72; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_76 = 32'h2e == io_ALUop ? xor_res : _alu_res_T_74; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_78 = 32'h8 == io_ALUop ? and_res : _alu_res_T_76; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_80 = 32'hd == io_ALUop ? _alu_res_T_19 : _alu_res_T_78; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_82 = 32'h16 == io_ALUop ? _alu_res_T_24 : _alu_res_T_80; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_84 = 32'h1c == io_ALUop ? _alu_res_T_29 : _alu_res_T_82; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_86 = 32'h1d == io_ALUop ? _alu_res_T_34 : _alu_res_T_84; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_88 = 32'h11 == io_ALUop ? mlu_res : _alu_res_T_86; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_90 = 32'h12 == io_ALUop ? _alu_res_T_38 : _alu_res_T_88; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_92 = 32'h13 == io_ALUop ? _alu_res_T_42 : _alu_res_T_90; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_94 = 32'h30 == io_ALUop ? divu_res : _alu_res_T_92; // @[Mux.scala 81:58]
  wire [64:0] _alu_res_T_96 = 32'h31 == io_ALUop ? div_res : {{1'd0}, _alu_res_T_94}; // @[Mux.scala 81:58]
  wire [64:0] _alu_res_T_98 = 32'h35 == io_ALUop ? {{1'd0}, _alu_res_T_46} : _alu_res_T_96; // @[Mux.scala 81:58]
  wire [64:0] _alu_res_T_100 = 32'h14 == io_ALUop ? {{1'd0}, _alu_res_T_50} : _alu_res_T_98; // @[Mux.scala 81:58]
  wire [64:0] _alu_res_T_102 = 32'h32 == io_ALUop ? {{1'd0}, _alu_res_T_54} : _alu_res_T_100; // @[Mux.scala 81:58]
  wire [64:0] _alu_res_T_104 = 32'h33 == io_ALUop ? {{1'd0}, remu_res} : _alu_res_T_102; // @[Mux.scala 81:58]
  wire [64:0] _alu_res_T_106 = 32'h34 == io_ALUop ? {{1'd0}, rem_res} : _alu_res_T_104; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_108 = 32'h37 == io_ALUop ? sll_res : {{62'd0}, _alu_res_T_106}; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_110 = 32'h39 == io_ALUop ? {{63'd0}, sra_res} : _alu_res_T_108; // @[Mux.scala 81:58]
  wire [126:0] alu_res = 32'h38 == io_ALUop ? {{63'd0}, srl_res} : _alu_res_T_110; // @[Mux.scala 81:58]
  assign io_alu_res = alu_res[63:0]; // @[ALU.scala 108:16]
endmodule
/* verilator lint_on WIDTH */
