module Register(
  input         clock,
  input  [4:0]  io_raddr1,
  input  [4:0]  io_raddr2,
  output [63:0] io_rdata1,
  output [63:0] io_rdata2,
  input         io_we,
  input  [4:0]  io_waddr,
  input  [63:0] io_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [63:0] Reg [0:31]; // @[register.scala 18:18]
  wire  Reg_io_rdata1_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_io_rdata1_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_io_rdata1_MPORT_data; // @[register.scala 18:18]
  wire  Reg_io_rdata2_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_io_rdata2_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_io_rdata2_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_0_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_0_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_0_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_1_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_1_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_1_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_2_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_2_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_2_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_3_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_3_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_3_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_4_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_4_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_4_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_5_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_5_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_5_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_6_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_6_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_6_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_7_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_7_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_7_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_8_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_8_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_8_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_9_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_9_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_9_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_10_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_10_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_10_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_11_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_11_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_11_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_12_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_12_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_12_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_13_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_13_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_13_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_14_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_14_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_14_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_15_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_15_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_15_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_16_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_16_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_16_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_17_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_17_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_17_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_18_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_18_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_18_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_19_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_19_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_19_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_20_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_20_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_20_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_21_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_21_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_21_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_22_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_22_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_22_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_23_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_23_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_23_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_24_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_24_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_24_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_25_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_25_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_25_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_26_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_26_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_26_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_27_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_27_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_27_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_28_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_28_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_28_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_29_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_29_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_29_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_30_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_30_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_30_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_31_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_31_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_31_MPORT_data; // @[register.scala 18:18]
  wire [63:0] Reg_MPORT_data; // @[register.scala 18:18]
  wire [4:0] Reg_MPORT_addr; // @[register.scala 18:18]
  wire  Reg_MPORT_mask; // @[register.scala 18:18]
  wire  Reg_MPORT_en; // @[register.scala 18:18]
  wire [63:0] reg_trace_input_reg_0; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_1; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_2; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_3; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_4; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_5; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_6; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_7; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_8; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_9; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_10; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_11; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_12; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_13; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_14; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_15; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_16; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_17; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_18; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_19; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_20; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_21; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_22; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_23; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_24; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_25; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_26; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_27; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_28; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_29; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_30; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_31; // @[register.scala 24:27]
  wire  _T = io_waddr != 5'h0; // @[register.scala 19:25]
  traceregs reg_trace ( // @[register.scala 24:27]
    .input_reg_0(reg_trace_input_reg_0),
    .input_reg_1(reg_trace_input_reg_1),
    .input_reg_2(reg_trace_input_reg_2),
    .input_reg_3(reg_trace_input_reg_3),
    .input_reg_4(reg_trace_input_reg_4),
    .input_reg_5(reg_trace_input_reg_5),
    .input_reg_6(reg_trace_input_reg_6),
    .input_reg_7(reg_trace_input_reg_7),
    .input_reg_8(reg_trace_input_reg_8),
    .input_reg_9(reg_trace_input_reg_9),
    .input_reg_10(reg_trace_input_reg_10),
    .input_reg_11(reg_trace_input_reg_11),
    .input_reg_12(reg_trace_input_reg_12),
    .input_reg_13(reg_trace_input_reg_13),
    .input_reg_14(reg_trace_input_reg_14),
    .input_reg_15(reg_trace_input_reg_15),
    .input_reg_16(reg_trace_input_reg_16),
    .input_reg_17(reg_trace_input_reg_17),
    .input_reg_18(reg_trace_input_reg_18),
    .input_reg_19(reg_trace_input_reg_19),
    .input_reg_20(reg_trace_input_reg_20),
    .input_reg_21(reg_trace_input_reg_21),
    .input_reg_22(reg_trace_input_reg_22),
    .input_reg_23(reg_trace_input_reg_23),
    .input_reg_24(reg_trace_input_reg_24),
    .input_reg_25(reg_trace_input_reg_25),
    .input_reg_26(reg_trace_input_reg_26),
    .input_reg_27(reg_trace_input_reg_27),
    .input_reg_28(reg_trace_input_reg_28),
    .input_reg_29(reg_trace_input_reg_29),
    .input_reg_30(reg_trace_input_reg_30),
    .input_reg_31(reg_trace_input_reg_31)
  );
  assign Reg_io_rdata1_MPORT_en = 1'h1;
  assign Reg_io_rdata1_MPORT_addr = io_raddr1;
  assign Reg_io_rdata1_MPORT_data = Reg[Reg_io_rdata1_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_io_rdata2_MPORT_en = 1'h1;
  assign Reg_io_rdata2_MPORT_addr = io_raddr2;
  assign Reg_io_rdata2_MPORT_data = Reg[Reg_io_rdata2_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_0_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_0_MPORT_addr = 5'h0;
  assign Reg_reg_trace_io_input_reg_0_MPORT_data = Reg[Reg_reg_trace_io_input_reg_0_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_1_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_1_MPORT_addr = 5'h1;
  assign Reg_reg_trace_io_input_reg_1_MPORT_data = Reg[Reg_reg_trace_io_input_reg_1_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_2_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_2_MPORT_addr = 5'h2;
  assign Reg_reg_trace_io_input_reg_2_MPORT_data = Reg[Reg_reg_trace_io_input_reg_2_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_3_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_3_MPORT_addr = 5'h3;
  assign Reg_reg_trace_io_input_reg_3_MPORT_data = Reg[Reg_reg_trace_io_input_reg_3_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_4_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_4_MPORT_addr = 5'h4;
  assign Reg_reg_trace_io_input_reg_4_MPORT_data = Reg[Reg_reg_trace_io_input_reg_4_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_5_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_5_MPORT_addr = 5'h5;
  assign Reg_reg_trace_io_input_reg_5_MPORT_data = Reg[Reg_reg_trace_io_input_reg_5_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_6_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_6_MPORT_addr = 5'h6;
  assign Reg_reg_trace_io_input_reg_6_MPORT_data = Reg[Reg_reg_trace_io_input_reg_6_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_7_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_7_MPORT_addr = 5'h7;
  assign Reg_reg_trace_io_input_reg_7_MPORT_data = Reg[Reg_reg_trace_io_input_reg_7_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_8_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_8_MPORT_addr = 5'h8;
  assign Reg_reg_trace_io_input_reg_8_MPORT_data = Reg[Reg_reg_trace_io_input_reg_8_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_9_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_9_MPORT_addr = 5'h9;
  assign Reg_reg_trace_io_input_reg_9_MPORT_data = Reg[Reg_reg_trace_io_input_reg_9_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_10_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_10_MPORT_addr = 5'ha;
  assign Reg_reg_trace_io_input_reg_10_MPORT_data = Reg[Reg_reg_trace_io_input_reg_10_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_11_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_11_MPORT_addr = 5'hb;
  assign Reg_reg_trace_io_input_reg_11_MPORT_data = Reg[Reg_reg_trace_io_input_reg_11_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_12_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_12_MPORT_addr = 5'hc;
  assign Reg_reg_trace_io_input_reg_12_MPORT_data = Reg[Reg_reg_trace_io_input_reg_12_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_13_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_13_MPORT_addr = 5'hd;
  assign Reg_reg_trace_io_input_reg_13_MPORT_data = Reg[Reg_reg_trace_io_input_reg_13_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_14_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_14_MPORT_addr = 5'he;
  assign Reg_reg_trace_io_input_reg_14_MPORT_data = Reg[Reg_reg_trace_io_input_reg_14_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_15_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_15_MPORT_addr = 5'hf;
  assign Reg_reg_trace_io_input_reg_15_MPORT_data = Reg[Reg_reg_trace_io_input_reg_15_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_16_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_16_MPORT_addr = 5'h10;
  assign Reg_reg_trace_io_input_reg_16_MPORT_data = Reg[Reg_reg_trace_io_input_reg_16_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_17_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_17_MPORT_addr = 5'h11;
  assign Reg_reg_trace_io_input_reg_17_MPORT_data = Reg[Reg_reg_trace_io_input_reg_17_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_18_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_18_MPORT_addr = 5'h12;
  assign Reg_reg_trace_io_input_reg_18_MPORT_data = Reg[Reg_reg_trace_io_input_reg_18_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_19_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_19_MPORT_addr = 5'h13;
  assign Reg_reg_trace_io_input_reg_19_MPORT_data = Reg[Reg_reg_trace_io_input_reg_19_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_20_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_20_MPORT_addr = 5'h14;
  assign Reg_reg_trace_io_input_reg_20_MPORT_data = Reg[Reg_reg_trace_io_input_reg_20_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_21_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_21_MPORT_addr = 5'h15;
  assign Reg_reg_trace_io_input_reg_21_MPORT_data = Reg[Reg_reg_trace_io_input_reg_21_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_22_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_22_MPORT_addr = 5'h16;
  assign Reg_reg_trace_io_input_reg_22_MPORT_data = Reg[Reg_reg_trace_io_input_reg_22_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_23_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_23_MPORT_addr = 5'h17;
  assign Reg_reg_trace_io_input_reg_23_MPORT_data = Reg[Reg_reg_trace_io_input_reg_23_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_24_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_24_MPORT_addr = 5'h18;
  assign Reg_reg_trace_io_input_reg_24_MPORT_data = Reg[Reg_reg_trace_io_input_reg_24_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_25_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_25_MPORT_addr = 5'h19;
  assign Reg_reg_trace_io_input_reg_25_MPORT_data = Reg[Reg_reg_trace_io_input_reg_25_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_26_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_26_MPORT_addr = 5'h1a;
  assign Reg_reg_trace_io_input_reg_26_MPORT_data = Reg[Reg_reg_trace_io_input_reg_26_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_27_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_27_MPORT_addr = 5'h1b;
  assign Reg_reg_trace_io_input_reg_27_MPORT_data = Reg[Reg_reg_trace_io_input_reg_27_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_28_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_28_MPORT_addr = 5'h1c;
  assign Reg_reg_trace_io_input_reg_28_MPORT_data = Reg[Reg_reg_trace_io_input_reg_28_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_29_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_29_MPORT_addr = 5'h1d;
  assign Reg_reg_trace_io_input_reg_29_MPORT_data = Reg[Reg_reg_trace_io_input_reg_29_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_30_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_30_MPORT_addr = 5'h1e;
  assign Reg_reg_trace_io_input_reg_30_MPORT_data = Reg[Reg_reg_trace_io_input_reg_30_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_31_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_31_MPORT_addr = 5'h1f;
  assign Reg_reg_trace_io_input_reg_31_MPORT_data = Reg[Reg_reg_trace_io_input_reg_31_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_MPORT_data = io_wdata;
  assign Reg_MPORT_addr = io_waddr;
  assign Reg_MPORT_mask = 1'h1;
  assign Reg_MPORT_en = io_we & _T;
  assign io_rdata1 = io_raddr1 == 5'h0 ? 64'h0 : Reg_io_rdata1_MPORT_data; // @[register.scala 22:21]
  assign io_rdata2 = io_raddr2 == 5'h0 ? 64'h0 : Reg_io_rdata2_MPORT_data; // @[register.scala 23:21]
  assign reg_trace_input_reg_0 = Reg_reg_trace_io_input_reg_0_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_1 = Reg_reg_trace_io_input_reg_1_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_2 = Reg_reg_trace_io_input_reg_2_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_3 = Reg_reg_trace_io_input_reg_3_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_4 = Reg_reg_trace_io_input_reg_4_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_5 = Reg_reg_trace_io_input_reg_5_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_6 = Reg_reg_trace_io_input_reg_6_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_7 = Reg_reg_trace_io_input_reg_7_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_8 = Reg_reg_trace_io_input_reg_8_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_9 = Reg_reg_trace_io_input_reg_9_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_10 = Reg_reg_trace_io_input_reg_10_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_11 = Reg_reg_trace_io_input_reg_11_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_12 = Reg_reg_trace_io_input_reg_12_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_13 = Reg_reg_trace_io_input_reg_13_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_14 = Reg_reg_trace_io_input_reg_14_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_15 = Reg_reg_trace_io_input_reg_15_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_16 = Reg_reg_trace_io_input_reg_16_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_17 = Reg_reg_trace_io_input_reg_17_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_18 = Reg_reg_trace_io_input_reg_18_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_19 = Reg_reg_trace_io_input_reg_19_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_20 = Reg_reg_trace_io_input_reg_20_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_21 = Reg_reg_trace_io_input_reg_21_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_22 = Reg_reg_trace_io_input_reg_22_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_23 = Reg_reg_trace_io_input_reg_23_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_24 = Reg_reg_trace_io_input_reg_24_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_25 = Reg_reg_trace_io_input_reg_25_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_26 = Reg_reg_trace_io_input_reg_26_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_27 = Reg_reg_trace_io_input_reg_27_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_28 = Reg_reg_trace_io_input_reg_28_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_29 = Reg_reg_trace_io_input_reg_29_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_30 = Reg_reg_trace_io_input_reg_30_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_31 = Reg_reg_trace_io_input_reg_31_MPORT_data; // @[register.scala 26:57]
  always @(posedge clock) begin
    if (Reg_MPORT_en & Reg_MPORT_mask) begin
      Reg[Reg_MPORT_addr] <= Reg_MPORT_data; // @[register.scala 18:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    Reg[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU(
  input         clock,
  input         reset,
  input         io_ds_allowin,
  input         io_br_taken,
  input  [63:0] io_br_target,
  output [63:0] io_to_ds_pc,
  output        io_fs_to_ds_valid,
  output [31:0] io_inst,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rlast,
  input         io_axi_in_rvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  input         io_fence,
  output        io_clear_cache,
  input         io_cache_init
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  fs_valid; // @[IFU.scala 29:27]
  reg  fs_ready_go; // @[IFU.scala 30:30]
  reg  cache_init; // @[IFU.scala 35:29]
  wire  fs_to_ds_valid = fs_valid & fs_ready_go; // @[IFU.scala 71:33]
  wire  _T = fs_to_ds_valid & io_ds_allowin; // @[IFU.scala 38:31]
  wire  _GEN_0 = fs_to_ds_valid & io_ds_allowin & cache_init ? 1'h0 : cache_init; // @[IFU.scala 38:60 39:20 35:29]
  wire  _GEN_1 = io_cache_init | _GEN_0; // @[IFU.scala 36:24 37:20]
  reg [63:0] fs_pc; // @[IFU.scala 42:24]
  reg [31:0] fs_inst; // @[IFU.scala 43:26]
  wire  _GEN_3 = io_axi_in_rvalid | fs_ready_go; // @[IFU.scala 56:27 58:21 30:30]
  wire [63:0] seq_pc = fs_pc + 64'h4; // @[IFU.scala 67:24]
  wire  fs_allowin = ~fs_valid | fs_ready_go & io_ds_allowin; // @[IFU.scala 72:29]
  wire  _GEN_5 = fs_allowin | fs_valid; // @[IFU.scala 74:36 75:18 29:27]
  reg  inst_ready; // @[IFU.scala 85:29]
  wire  _GEN_7 = io_axi_in_rvalid & inst_ready & io_axi_in_rlast ? 1'h0 : 1'h1; // @[IFU.scala 86:60 87:20 89:20]
  assign io_to_ds_pc = fs_pc; // @[IFU.scala 82:17]
  assign io_fs_to_ds_valid = fs_valid & fs_ready_go; // @[IFU.scala 71:33]
  assign io_inst = fs_inst; // @[IFU.scala 108:13]
  assign io_axi_out_araddr = fs_pc[31:0]; // @[IFU.scala 92:31]
  assign io_axi_out_arvalid = fs_valid & ~fs_ready_go; // @[IFU.scala 93:36]
  assign io_axi_out_rready = inst_ready; // @[IFU.scala 97:23]
  assign io_clear_cache = io_fence & ~cache_init; // @[IFU.scala 54:32]
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 29:27]
      fs_valid <= 1'h0; // @[IFU.scala 29:27]
    end else begin
      fs_valid <= _GEN_5;
    end
    if (reset) begin // @[IFU.scala 30:30]
      fs_ready_go <= 1'h0; // @[IFU.scala 30:30]
    end else if (_T) begin // @[IFU.scala 60:42]
      fs_ready_go <= 1'h0; // @[IFU.scala 61:21]
    end else begin
      fs_ready_go <= _GEN_3;
    end
    if (reset) begin // @[IFU.scala 35:29]
      cache_init <= 1'h0; // @[IFU.scala 35:29]
    end else begin
      cache_init <= _GEN_1;
    end
    if (reset) begin // @[IFU.scala 42:24]
      fs_pc <= 64'h7ffffffc; // @[IFU.scala 42:24]
    end else if (fs_allowin) begin // @[IFU.scala 74:36]
      if (io_br_taken) begin // @[IFU.scala 68:19]
        fs_pc <= io_br_target;
      end else begin
        fs_pc <= seq_pc;
      end
    end
    if (reset) begin // @[IFU.scala 43:26]
      fs_inst <= 32'h0; // @[IFU.scala 43:26]
    end else if (io_axi_in_rvalid) begin // @[IFU.scala 56:27]
      fs_inst <= io_axi_in_rdata[31:0]; // @[IFU.scala 57:17]
    end
    inst_ready <= reset | _GEN_7; // @[IFU.scala 85:{29,29}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fs_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  fs_ready_go = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cache_init = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  fs_pc = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  fs_inst = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  inst_ready = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module csr_reg(
  input         clock,
  input         io_wen1,
  input         io_wen2,
  input  [1:0]  io_waddr1,
  input  [63:0] io_wdata1,
  input  [63:0] io_wdata2,
  input  [1:0]  io_raddr,
  output [63:0] io_rdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [63:0] CSR_Reg [0:3]; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_io_rdata_MPORT_en; // @[csr_reg.scala 19:22]
  wire [1:0] CSR_Reg_io_rdata_MPORT_addr; // @[csr_reg.scala 19:22]
  wire [63:0] CSR_Reg_io_rdata_MPORT_data; // @[csr_reg.scala 19:22]
  wire [63:0] CSR_Reg_MPORT_data; // @[csr_reg.scala 19:22]
  wire [1:0] CSR_Reg_MPORT_addr; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_MPORT_mask; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_MPORT_en; // @[csr_reg.scala 19:22]
  wire [63:0] CSR_Reg_MPORT_1_data; // @[csr_reg.scala 19:22]
  wire [1:0] CSR_Reg_MPORT_1_addr; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_MPORT_1_mask; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_MPORT_1_en; // @[csr_reg.scala 19:22]
  assign CSR_Reg_io_rdata_MPORT_en = 1'h1;
  assign CSR_Reg_io_rdata_MPORT_addr = io_raddr;
  assign CSR_Reg_io_rdata_MPORT_data = CSR_Reg[CSR_Reg_io_rdata_MPORT_addr]; // @[csr_reg.scala 19:22]
  assign CSR_Reg_MPORT_data = io_wdata1;
  assign CSR_Reg_MPORT_addr = io_waddr1;
  assign CSR_Reg_MPORT_mask = 1'h1;
  assign CSR_Reg_MPORT_en = io_wen1;
  assign CSR_Reg_MPORT_1_data = io_wdata2;
  assign CSR_Reg_MPORT_1_addr = 2'h3;
  assign CSR_Reg_MPORT_1_mask = 1'h1;
  assign CSR_Reg_MPORT_1_en = io_wen2;
  assign io_rdata = CSR_Reg_io_rdata_MPORT_data; // @[csr_reg.scala 26:14]
  always @(posedge clock) begin
    if (CSR_Reg_MPORT_en & CSR_Reg_MPORT_mask) begin
      CSR_Reg[CSR_Reg_MPORT_addr] <= CSR_Reg_MPORT_data; // @[csr_reg.scala 19:22]
    end
    if (CSR_Reg_MPORT_1_en & CSR_Reg_MPORT_1_mask) begin
      CSR_Reg[CSR_Reg_MPORT_1_addr] <= CSR_Reg_MPORT_1_data; // @[csr_reg.scala 19:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    CSR_Reg[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_fs_to_ds_valid,
  output        io_ds_to_es_valid,
  input         io_es_allowin,
  input  [31:0] io_from_fs_inst,
  output        io_br_taken,
  output [63:0] io_br_target,
  output        io_ds_allowin,
  output        io_fence,
  output [4:0]  io_raddr1,
  output [4:0]  io_raddr2,
  input  [63:0] io_rdata1,
  input  [63:0] io_rdata2,
  output [63:0] io_to_es_pc,
  output [31:0] io_ALUop,
  output [63:0] io_src1,
  output [63:0] io_src2,
  output [4:0]  io_rf_dst,
  output [63:0] io_store_data,
  output        io_ctrl_sign_reg_write,
  output        io_ctrl_sign_Writemem_en,
  output        io_ctrl_sign_Readmem_en,
  output [7:0]  io_ctrl_sign_Wmask,
  output [2:0]  io_load_type,
  input         io_es_ld,
  input  [63:0] io_es_fwd_res,
  input  [63:0] io_ms_fwd_res,
  input  [63:0] io_ws_fwd_res,
  input         io_es_fwd_ready,
  input         io_ms_fwd_ready,
  input         io_es_rf_we,
  input         io_ms_rf_we,
  input         io_ws_rf_we,
  input         io_es_valid,
  input         io_ms_valid,
  input         io_ws_valid,
  input  [4:0]  io_es_rf_dst,
  input  [4:0]  io_ms_rf_dst,
  input  [4:0]  io_ws_rf_dst,
  output        io_ds_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  csr_reg_clock; // @[IDU.scala 448:21]
  wire  csr_reg_io_wen1; // @[IDU.scala 448:21]
  wire  csr_reg_io_wen2; // @[IDU.scala 448:21]
  wire [1:0] csr_reg_io_waddr1; // @[IDU.scala 448:21]
  wire [63:0] csr_reg_io_wdata1; // @[IDU.scala 448:21]
  wire [63:0] csr_reg_io_wdata2; // @[IDU.scala 448:21]
  wire [1:0] csr_reg_io_raddr; // @[IDU.scala 448:21]
  wire [63:0] csr_reg_io_rdata; // @[IDU.scala 448:21]
  reg  ds_valid; // @[IDU.scala 111:27]
  reg [63:0] ds_pc; // @[IDU.scala 115:24]
  reg [31:0] inst; // @[IDU.scala 117:23]
  reg  br_taken_cancel; // @[IDU.scala 121:34]
  wire [31:0] _src1_is_pc_T = inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_1 = 32'h6f == _src1_is_pc_T; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_3 = 32'h17 == _src1_is_pc_T; // @[Lookup.scala 31:38]
  wire [31:0] _src1_is_pc_T_4 = inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_5 = 32'h1063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_7 = 32'h63 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_9 = 32'h5063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_11 = 32'h4063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_13 = 32'h6063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_15 = 32'h7063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  src1_is_pc = _src1_is_pc_T_1 | (_src1_is_pc_T_3 | (_src1_is_pc_T_5 | (_src1_is_pc_T_7 | (_src1_is_pc_T_9 | (
    _src1_is_pc_T_11 | (_src1_is_pc_T_13 | _src1_is_pc_T_15)))))); // @[Lookup.scala 34:39]
  wire  _inst_type_T_1 = 32'h13 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_5 = 32'h37 == _src1_is_pc_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_9 = 32'h67 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_11 = 32'h3023 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_13 = 32'h3013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_15 = 32'h2003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_16 = inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_17 = 32'h3b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_19 = 32'h40000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_25 = 32'h3003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_27 = 32'h1b == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_29 = 32'h33 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_30 = inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_31 = 32'h40005013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_33 = 32'h4003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_35 = 32'h1023 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_37 = 32'h23 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_39 = 32'h6033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_41 = 32'h4013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_43 = 32'h7033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_45 = 32'h7013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_47 = 32'h4000003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_49 = 32'h103b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_51 = 32'h1013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_53 = 32'h5013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_55 = 32'h101b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_57 = 32'h4000501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_59 = 32'h501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_61 = 32'h4000503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_63 = 32'h503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_65 = 32'h3033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_67 = 32'h2033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_75 = 32'h2023 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_77 = 32'h1003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_79 = 32'h5003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_81 = 32'h2000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_83 = 32'h200003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_85 = 32'h200403b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_87 = 32'h200603b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_89 = 32'h4033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_91 = 32'h6013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_93 = 32'h2005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_95 = 32'h2004033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_97 = 32'h200503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_99 = 32'h200703b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_101 = 32'h2007033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_103 = 32'h2006033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_105 = 32'h1033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_107 = 32'h5033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_109 = 32'h40005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_111 = 32'h2013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_113 = 32'h6003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_115 = 32'h3 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_119 = 32'h73 == inst; // @[Lookup.scala 31:38]
  wire  _inst_type_T_121 = 32'h1073 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_123 = 32'h2073 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_125 = 32'h3073 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire [6:0] _inst_type_T_126 = _inst_type_T_125 ? 7'h40 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_127 = _inst_type_T_123 ? 7'h40 : _inst_type_T_126; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_128 = _inst_type_T_121 ? 7'h40 : _inst_type_T_127; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_129 = _inst_type_T_119 ? 7'h40 : _inst_type_T_128; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_130 = _src1_is_pc_T_15 ? 7'h45 : _inst_type_T_129; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_131 = _inst_type_T_115 ? 7'h40 : _inst_type_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_132 = _inst_type_T_113 ? 7'h40 : _inst_type_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_133 = _inst_type_T_111 ? 7'h40 : _inst_type_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_134 = _inst_type_T_109 ? 7'h41 : _inst_type_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_135 = _inst_type_T_107 ? 7'h41 : _inst_type_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_136 = _inst_type_T_105 ? 7'h41 : _inst_type_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_137 = _inst_type_T_103 ? 7'h41 : _inst_type_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_138 = _inst_type_T_101 ? 7'h41 : _inst_type_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_139 = _inst_type_T_99 ? 7'h41 : _inst_type_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_140 = _inst_type_T_97 ? 7'h41 : _inst_type_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_141 = _inst_type_T_95 ? 7'h41 : _inst_type_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_142 = _inst_type_T_93 ? 7'h41 : _inst_type_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_143 = _inst_type_T_91 ? 7'h40 : _inst_type_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_144 = _inst_type_T_89 ? 7'h41 : _inst_type_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_145 = _inst_type_T_87 ? 7'h41 : _inst_type_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_146 = _inst_type_T_85 ? 7'h41 : _inst_type_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_147 = _inst_type_T_83 ? 7'h41 : _inst_type_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_148 = _inst_type_T_81 ? 7'h41 : _inst_type_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_149 = _inst_type_T_79 ? 7'h40 : _inst_type_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_150 = _inst_type_T_77 ? 7'h40 : _inst_type_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_151 = _inst_type_T_75 ? 7'h44 : _inst_type_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_152 = _src1_is_pc_T_13 ? 7'h45 : _inst_type_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_153 = _src1_is_pc_T_11 ? 7'h45 : _inst_type_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_154 = _src1_is_pc_T_9 ? 7'h45 : _inst_type_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_155 = _inst_type_T_67 ? 7'h41 : _inst_type_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_156 = _inst_type_T_65 ? 7'h41 : _inst_type_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_157 = _inst_type_T_63 ? 7'h41 : _inst_type_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_158 = _inst_type_T_61 ? 7'h41 : _inst_type_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_159 = _inst_type_T_59 ? 7'h40 : _inst_type_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_160 = _inst_type_T_57 ? 7'h40 : _inst_type_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_161 = _inst_type_T_55 ? 7'h40 : _inst_type_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_162 = _inst_type_T_53 ? 7'h40 : _inst_type_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_163 = _inst_type_T_51 ? 7'h40 : _inst_type_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_164 = _inst_type_T_49 ? 7'h41 : _inst_type_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_165 = _inst_type_T_47 ? 7'h41 : _inst_type_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_166 = _inst_type_T_45 ? 7'h40 : _inst_type_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_167 = _inst_type_T_43 ? 7'h41 : _inst_type_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_168 = _inst_type_T_41 ? 7'h40 : _inst_type_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_169 = _inst_type_T_39 ? 7'h41 : _inst_type_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_170 = _inst_type_T_37 ? 7'h44 : _inst_type_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_171 = _inst_type_T_35 ? 7'h44 : _inst_type_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_172 = _inst_type_T_33 ? 7'h40 : _inst_type_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_173 = _inst_type_T_31 ? 7'h40 : _inst_type_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_174 = _inst_type_T_29 ? 7'h41 : _inst_type_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_175 = _inst_type_T_27 ? 7'h40 : _inst_type_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_176 = _inst_type_T_25 ? 7'h40 : _inst_type_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_177 = _src1_is_pc_T_7 ? 7'h45 : _inst_type_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_178 = _src1_is_pc_T_5 ? 7'h45 : _inst_type_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_179 = _inst_type_T_19 ? 7'h41 : _inst_type_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_180 = _inst_type_T_17 ? 7'h41 : _inst_type_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_181 = _inst_type_T_15 ? 7'h40 : _inst_type_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_182 = _inst_type_T_13 ? 7'h40 : _inst_type_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_183 = _inst_type_T_11 ? 7'h44 : _inst_type_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_184 = _inst_type_T_9 ? 7'h40 : _inst_type_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_185 = _src1_is_pc_T_1 ? 7'h43 : _inst_type_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_186 = _inst_type_T_5 ? 7'h42 : _inst_type_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_187 = _src1_is_pc_T_3 ? 7'h42 : _inst_type_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_188 = _inst_type_T_1 ? 7'h40 : _inst_type_T_187; // @[Lookup.scala 34:39]
  wire [31:0] inst_type = {{25'd0}, _inst_type_T_188}; // @[IDU.scala 236:15 65:25]
  wire  _conflict_es_rs1_T_1 = inst_type == 32'h45; // @[IDU.scala 491:47]
  wire  _csr_write_T_10 = _inst_type_T_121 | (_inst_type_T_123 | _inst_type_T_125); // @[Lookup.scala 34:39]
  wire [1:0] csr_write = _inst_type_T_119 ? 2'h3 : {{1'd0}, _csr_write_T_10}; // @[Lookup.scala 34:39]
  wire  _conflict_es_rs1_T_3 = csr_write == 2'h1; // @[IDU.scala 491:72]
  wire  _conflict_es_rs1_T_4 = ~src1_is_pc | inst_type == 32'h45 | csr_write == 2'h1; // @[IDU.scala 491:59]
  wire [4:0] rs1 = inst[19:15]; // @[IDU.scala 226:16]
  wire  _conflict_es_rs1_T_6 = rs1 != 5'h0; // @[IDU.scala 491:111]
  wire  conflict_es_rs1 = (~src1_is_pc | inst_type == 32'h45 | csr_write == 2'h1) & (rs1 == io_es_rf_dst & rs1 != 5'h0
     & io_es_rf_we & io_es_valid); // @[IDU.scala 491:81]
  wire  src2_is_imm = 32'h45 == inst_type | (32'h43 == inst_type | (32'h44 == inst_type | (32'h42 == inst_type | 32'h40
     == inst_type))); // @[Mux.scala 81:58]
  wire  _conflict_es_rs2_T_5 = csr_write == 2'h3; // @[IDU.scala 494:92]
  wire  _conflict_es_rs2_T_6 = ~src2_is_imm | inst_type == 32'h44 | _conflict_es_rs1_T_1 | csr_write == 2'h3; // @[IDU.scala 494:81]
  wire [4:0] rs2 = csr_write[0] ? 5'h11 : inst[24:20]; // @[IDU.scala 225:15]
  wire  _conflict_es_rs2_T_8 = rs2 != 5'h0; // @[IDU.scala 494:130]
  wire  conflict_es_rs2 = (~src2_is_imm | inst_type == 32'h44 | _conflict_es_rs1_T_1 | csr_write == 2'h3) & (rs2 ==
    io_es_rf_dst & rs2 != 5'h0 & io_es_rf_we & io_es_valid); // @[IDU.scala 494:100]
  wire  conflict_ms_rs1 = _conflict_es_rs1_T_4 & (rs1 == io_ms_rf_dst & _conflict_es_rs1_T_6 & io_ms_rf_we & io_ms_valid
    ); // @[IDU.scala 492:81]
  wire  conflict_ms_rs2 = _conflict_es_rs2_T_6 & (rs2 == io_ms_rf_dst & _conflict_es_rs2_T_8 & io_ms_rf_we & io_ms_valid
    ); // @[IDU.scala 495:100]
  wire  conflict_ws_rs1 = _conflict_es_rs1_T_4 & (rs1 == io_ws_rf_dst & _conflict_es_rs1_T_6 & io_ws_rf_we & io_ws_valid
    ); // @[IDU.scala 493:81]
  wire  conflict_ws_rs2 = _conflict_es_rs2_T_6 & (rs2 == io_ws_rf_dst & _conflict_es_rs2_T_8 & io_ws_rf_we & io_ws_valid
    ); // @[IDU.scala 496:100]
  wire  _ALUop_T_3 = 32'h100073 == inst; // @[Lookup.scala 31:38]
  wire  _ALUop_T_111 = 32'h30200073 == inst; // @[Lookup.scala 31:38]
  wire [6:0] _ALUop_T_118 = _inst_type_T_125 ? 7'h47 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_119 = _inst_type_T_123 ? 7'h46 : _ALUop_T_118; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_120 = _inst_type_T_121 ? 7'h3f : _ALUop_T_119; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_121 = _ALUop_T_111 ? 7'h3e : _ALUop_T_120; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_122 = _inst_type_T_119 ? 7'h3d : _ALUop_T_121; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_123 = _inst_type_T_115 ? 7'hf : _ALUop_T_122; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_124 = _inst_type_T_113 ? 7'hf : _ALUop_T_123; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_125 = _inst_type_T_111 ? 7'h1f : _ALUop_T_124; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_126 = _inst_type_T_109 ? 7'h39 : _ALUop_T_125; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_127 = _inst_type_T_107 ? 7'h38 : _ALUop_T_126; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_128 = _inst_type_T_105 ? 7'h37 : _ALUop_T_127; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_129 = _inst_type_T_103 ? 7'h34 : _ALUop_T_128; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_130 = _inst_type_T_101 ? 7'h33 : _ALUop_T_129; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_131 = _inst_type_T_99 ? 7'h32 : _ALUop_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_132 = _inst_type_T_97 ? 7'h35 : _ALUop_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_133 = _inst_type_T_95 ? 7'h31 : _ALUop_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_134 = _inst_type_T_93 ? 7'h30 : _ALUop_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_135 = _inst_type_T_91 ? 7'hb : _ALUop_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_136 = _inst_type_T_89 ? 7'h2e : _ALUop_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_137 = _inst_type_T_87 ? 7'h14 : _ALUop_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_138 = _inst_type_T_85 ? 7'h13 : _ALUop_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_139 = _inst_type_T_83 ? 7'h12 : _ALUop_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_140 = _inst_type_T_81 ? 7'h11 : _ALUop_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_141 = _inst_type_T_79 ? 7'hf : _ALUop_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_142 = _inst_type_T_77 ? 7'hf : _ALUop_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_143 = _inst_type_T_75 ? 7'hf : _ALUop_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_144 = _inst_type_T_67 ? 7'h1f : _ALUop_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_145 = _inst_type_T_65 ? 7'h1e : _ALUop_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_146 = _inst_type_T_63 ? 7'h1d : _ALUop_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_147 = _inst_type_T_61 ? 7'h1c : _ALUop_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_148 = _inst_type_T_59 ? 7'h1d : _ALUop_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_149 = _inst_type_T_57 ? 7'h1c : _ALUop_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_150 = _inst_type_T_55 ? 7'h16 : _ALUop_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_151 = _inst_type_T_53 ? 7'h38 : _ALUop_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_152 = _inst_type_T_51 ? 7'h37 : _ALUop_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_153 = _inst_type_T_49 ? 7'h16 : _ALUop_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_154 = _inst_type_T_47 ? 7'hd : _ALUop_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_155 = _inst_type_T_45 ? 7'h8 : _ALUop_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_156 = _inst_type_T_43 ? 7'h8 : _ALUop_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_157 = _inst_type_T_41 ? 7'h2e : _ALUop_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_158 = _inst_type_T_39 ? 7'hb : _ALUop_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_159 = _inst_type_T_37 ? 7'hf : _ALUop_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_160 = _inst_type_T_35 ? 7'hf : _ALUop_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_161 = _inst_type_T_33 ? 7'hf : _ALUop_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_162 = _inst_type_T_31 ? 7'h15 : _ALUop_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_163 = _inst_type_T_29 ? 7'hf : _ALUop_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_164 = _inst_type_T_27 ? 7'hc : _ALUop_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_165 = _inst_type_T_25 ? 7'hf : _ALUop_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_166 = _inst_type_T_19 ? 7'he : _ALUop_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_167 = _inst_type_T_17 ? 7'hc : _ALUop_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_168 = _inst_type_T_15 ? 7'hf : _ALUop_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_169 = _inst_type_T_13 ? 7'h1e : _ALUop_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_170 = _inst_type_T_11 ? 7'hf : _ALUop_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_171 = _inst_type_T_9 ? 7'h6 : _ALUop_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_172 = _src1_is_pc_T_1 ? 7'h5 : _ALUop_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_173 = _inst_type_T_5 ? 7'h4 : _ALUop_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_174 = _src1_is_pc_T_3 ? 7'hf : _ALUop_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_175 = _ALUop_T_3 ? 7'h2 : _ALUop_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_176 = _inst_type_T_1 ? 7'hf : _ALUop_T_175; // @[Lookup.scala 34:39]
  wire [31:0] ALUop = {{25'd0}, _ALUop_T_176}; // @[IDU.scala 310:11 64:21]
  wire  _ds_ready_go_T_30 = ALUop == 32'h6 & io_fs_to_ds_valid & ds_valid | ALUop != 32'h6; // @[IDU.scala 150:473]
  wire  ds_ready_go = ((conflict_es_rs1 | conflict_es_rs2) & (io_es_fwd_ready & ~io_es_ld) | ~(conflict_es_rs1 |
    conflict_es_rs2) & (conflict_ms_rs1 | conflict_ms_rs2) & io_ms_fwd_ready | ~(conflict_es_rs1 | conflict_es_rs2) & ~(
    conflict_ms_rs1 | conflict_ms_rs2) & (conflict_ws_rs1 | conflict_ws_rs2) | ~(conflict_es_rs1 | conflict_es_rs2 |
    conflict_ms_rs1 | conflict_ms_rs2 | conflict_ws_rs1 | conflict_ws_rs2)) & _ds_ready_go_T_30; // @[IDU.scala 150:419]
  wire  ds_allowin = ~ds_valid | ds_ready_go & io_es_allowin; // @[IDU.scala 152:29]
  wire  _T_1 = ~br_taken_cancel; // @[IDU.scala 133:26]
  wire [63:0] _rdata1_T = conflict_ws_rs1 ? io_ws_fwd_res : io_rdata1; // @[IDU.scala 497:86]
  wire [63:0] _rdata1_T_1 = conflict_ms_rs1 ? io_ms_fwd_res : _rdata1_T; // @[IDU.scala 497:52]
  wire [63:0] rdata1 = conflict_es_rs1 ? io_es_fwd_res : _rdata1_T_1; // @[IDU.scala 497:18]
  wire [63:0] _br_taken_T = conflict_es_rs1 ? io_es_fwd_res : _rdata1_T_1; // @[IDU.scala 482:27]
  wire [63:0] _rdata2_T = conflict_ws_rs2 ? io_ws_fwd_res : io_rdata2; // @[IDU.scala 498:86]
  wire [63:0] _rdata2_T_1 = conflict_ms_rs2 ? io_ms_fwd_res : _rdata2_T; // @[IDU.scala 498:52]
  wire [63:0] rdata2 = conflict_es_rs2 ? io_es_fwd_res : _rdata2_T_1; // @[IDU.scala 498:18]
  wire [63:0] _br_taken_T_1 = conflict_es_rs2 ? io_es_fwd_res : _rdata2_T_1; // @[IDU.scala 482:45]
  wire  _br_taken_T_2 = $signed(_br_taken_T) != $signed(_br_taken_T_1); // @[IDU.scala 482:34]
  wire  _br_taken_T_6 = $signed(_br_taken_T) == $signed(_br_taken_T_1); // @[IDU.scala 483:34]
  wire  _br_taken_T_10 = $signed(_br_taken_T) >= $signed(_br_taken_T_1); // @[IDU.scala 484:34]
  wire  _br_taken_T_14 = $signed(_br_taken_T) < $signed(_br_taken_T_1); // @[IDU.scala 485:34]
  wire  _br_taken_T_16 = rdata1 < rdata2; // @[IDU.scala 486:28]
  wire  _br_taken_T_18 = rdata1 >= rdata2; // @[IDU.scala 487:28]
  wire  _br_taken_T_42 = _src1_is_pc_T_15 ? _br_taken_T_18 : _inst_type_T_119 | _ALUop_T_111; // @[Lookup.scala 34:39]
  wire  _br_taken_T_43 = _src1_is_pc_T_13 ? _br_taken_T_16 : _br_taken_T_42; // @[Lookup.scala 34:39]
  wire  _br_taken_T_44 = _src1_is_pc_T_11 ? _br_taken_T_14 : _br_taken_T_43; // @[Lookup.scala 34:39]
  wire  _br_taken_T_45 = _src1_is_pc_T_9 ? _br_taken_T_10 : _br_taken_T_44; // @[Lookup.scala 34:39]
  wire  _br_taken_T_46 = _src1_is_pc_T_7 ? _br_taken_T_6 : _br_taken_T_45; // @[Lookup.scala 34:39]
  wire  _br_taken_T_47 = _src1_is_pc_T_5 ? _br_taken_T_2 : _br_taken_T_46; // @[Lookup.scala 34:39]
  wire  br_taken = _src1_is_pc_T_1 | (_inst_type_T_9 | _br_taken_T_47); // @[Lookup.scala 34:39]
  wire  _T_2 = br_taken & ~br_taken_cancel; // @[IDU.scala 133:23]
  wire [4:0] rd = inst[11:7]; // @[IDU.scala 227:15]
  wire  fence = 32'h100f == inst; // @[Lookup.scala 31:38]
  wire [11:0] imm_imm = inst[31:20]; // @[IDU.scala 82:23]
  wire [51:0] _imm_T_2 = imm_imm[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_3 = {_imm_T_2,imm_imm}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_1 = {inst[31],inst[19:12],inst[20],inst[30:21]}; // @[Cat.scala 31:58]
  wire [42:0] _imm_T_6 = imm_imm_1[19] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_7 = {_imm_T_6,inst[31],inst[19:12],inst[20],inst[30:21],1'h0}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_2 = inst[31:12]; // @[IDU.scala 86:23]
  wire [31:0] _imm_T_10 = imm_imm_2[19] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_12 = {_imm_T_10,imm_imm_2,12'h0}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_3 = {inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [51:0] _imm_T_15 = imm_imm_3[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_16 = {_imm_T_15,inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_4 = {inst[31],inst[7],inst[30:25],inst[11:8]}; // @[Cat.scala 31:58]
  wire [50:0] _imm_T_19 = imm_imm_4[11] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_20 = {_imm_T_19,inst[31],inst[7],inst[30:25],inst[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [63:0] _imm_T_22 = 32'h40 == inst_type ? _imm_T_3 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_24 = 32'h43 == inst_type ? _imm_T_7 : _imm_T_22; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_26 = 32'h42 == inst_type ? _imm_T_12 : _imm_T_24; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_28 = 32'h44 == inst_type ? _imm_T_16 : _imm_T_26; // @[Mux.scala 81:58]
  wire [63:0] imm = 32'h45 == inst_type ? _imm_T_20 : _imm_T_28; // @[Mux.scala 81:58]
  wire  _reg_write_T_28 = fence ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _reg_write_T_29 = _ALUop_T_111 ? 1'h0 : _reg_write_T_28; // @[Lookup.scala 34:39]
  wire  _reg_write_T_30 = _inst_type_T_119 ? 1'h0 : _reg_write_T_29; // @[Lookup.scala 34:39]
  wire  _reg_write_T_31 = _src1_is_pc_T_15 ? 1'h0 : _reg_write_T_30; // @[Lookup.scala 34:39]
  wire  _reg_write_T_32 = _src1_is_pc_T_13 ? 1'h0 : _reg_write_T_31; // @[Lookup.scala 34:39]
  wire  _reg_write_T_33 = _src1_is_pc_T_11 ? 1'h0 : _reg_write_T_32; // @[Lookup.scala 34:39]
  wire  _reg_write_T_34 = _src1_is_pc_T_9 ? 1'h0 : _reg_write_T_33; // @[Lookup.scala 34:39]
  wire  _reg_write_T_35 = _src1_is_pc_T_7 ? 1'h0 : _reg_write_T_34; // @[Lookup.scala 34:39]
  wire  _reg_write_T_36 = _src1_is_pc_T_5 ? 1'h0 : _reg_write_T_35; // @[Lookup.scala 34:39]
  wire  _reg_write_T_37 = _inst_type_T_75 ? 1'h0 : _reg_write_T_36; // @[Lookup.scala 34:39]
  wire  _reg_write_T_38 = _inst_type_T_37 ? 1'h0 : _reg_write_T_37; // @[Lookup.scala 34:39]
  wire  _reg_write_T_39 = _inst_type_T_35 ? 1'h0 : _reg_write_T_38; // @[Lookup.scala 34:39]
  wire  _reg_write_T_40 = _inst_type_T_11 ? 1'h0 : _reg_write_T_39; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_14 = _inst_type_T_79 ? 3'h7 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_15 = _inst_type_T_115 ? 3'h6 : _load_type_T_14; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_16 = _inst_type_T_77 ? 3'h5 : _load_type_T_15; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_17 = _inst_type_T_113 ? 3'h4 : _load_type_T_16; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_18 = _inst_type_T_33 ? 3'h3 : _load_type_T_17; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_19 = _inst_type_T_25 ? 3'h2 : _load_type_T_18; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_8 = _inst_type_T_75 ? 4'hf : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_9 = _inst_type_T_37 ? 4'h1 : _Wmask_T_8; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_10 = _inst_type_T_35 ? 4'h3 : _Wmask_T_9; // @[Lookup.scala 34:39]
  wire [1:0] _csr_index_T_6 = 12'h300 == imm[11:0] ? 2'h2 : {{1'd0}, 12'h341 == imm[11:0]}; // @[Mux.scala 81:58]
  wire [1:0] csr_index = 12'h342 == imm[11:0] ? 2'h3 : _csr_index_T_6; // @[Mux.scala 81:58]
  wire [63:0] _csr_wdata_T = rdata1 | csr_reg_io_rdata; // @[IDU.scala 457:26]
  wire [63:0] _csr_wdata_T_1 = ~csr_reg_io_rdata; // @[IDU.scala 458:29]
  wire [63:0] _csr_wdata_T_2 = rdata1 & _csr_wdata_T_1; // @[IDU.scala 458:26]
  wire [63:0] _csr_wdata_T_9 = _inst_type_T_125 ? _csr_wdata_T_2 : 64'h0; // @[Lookup.scala 34:39]
  wire [63:0] _csr_wdata_T_10 = _inst_type_T_123 ? _csr_wdata_T : _csr_wdata_T_9; // @[Lookup.scala 34:39]
  wire [63:0] csr_wdata = _inst_type_T_121 ? rdata1 : _csr_wdata_T_10; // @[Lookup.scala 34:39]
  wire [1:0] _T_11 = ALUop == 32'h3e ? 2'h1 : csr_index; // @[IDU.scala 461:48]
  wire [1:0] _T_18 = _conflict_es_rs1_T_3 ? csr_index : 2'h0; // @[IDU.scala 463:46]
  wire [63:0] _T_22 = _conflict_es_rs1_T_3 ? csr_wdata : 64'h0; // @[IDU.scala 464:48]
  wire [63:0] src1 = src1_is_pc ? ds_pc : rdata1; // @[IDU.scala 470:16]
  wire [63:0] src2 = src2_is_imm ? imm : rdata2; // @[IDU.scala 471:16]
  wire [63:0] _br_target_T_1 = src1 + src2; // @[IDU.scala 474:35]
  wire [63:0] _br_target_T_4 = _br_target_T_1 & 64'hfffffffffffffffe; // @[IDU.scala 475:31]
  wire [63:0] _br_target_T_6 = csr_reg_io_rdata + 64'h4; // @[IDU.scala 477:28]
  wire [63:0] _br_target_T_13 = _ALUop_T_111 ? _br_target_T_6 : _br_target_T_1; // @[Lookup.scala 34:39]
  wire [63:0] _br_target_T_14 = _inst_type_T_119 ? csr_reg_io_rdata : _br_target_T_13; // @[Lookup.scala 34:39]
  wire [31:0] _io_store_data_T_11 = _inst_type_T_75 ? rdata2[31:0] : 32'h0; // @[Lookup.scala 34:39]
  wire [31:0] _io_store_data_T_12 = _inst_type_T_37 ? {{24'd0}, rdata2[7:0]} : _io_store_data_T_11; // @[Lookup.scala 34:39]
  wire [31:0] _io_store_data_T_13 = _inst_type_T_35 ? {{16'd0}, rdata2[15:0]} : _io_store_data_T_12; // @[Lookup.scala 34:39]
  csr_reg csr_reg ( // @[IDU.scala 448:21]
    .clock(csr_reg_clock),
    .io_wen1(csr_reg_io_wen1),
    .io_wen2(csr_reg_io_wen2),
    .io_waddr1(csr_reg_io_waddr1),
    .io_wdata1(csr_reg_io_wdata1),
    .io_wdata2(csr_reg_io_wdata2),
    .io_raddr(csr_reg_io_raddr),
    .io_rdata(csr_reg_io_rdata)
  );
  assign io_ds_to_es_valid = ds_valid & ds_ready_go; // @[IDU.scala 151:32]
  assign io_br_taken = br_taken & _T_1; // @[IDU.scala 502:29]
  assign io_br_target = _inst_type_T_9 ? _br_target_T_4 : _br_target_T_14; // @[Lookup.scala 34:39]
  assign io_ds_allowin = ~ds_valid | ds_ready_go & io_es_allowin; // @[IDU.scala 152:29]
  assign io_fence = 32'h100f == inst; // @[Lookup.scala 31:38]
  assign io_raddr1 = inst[19:15]; // @[IDU.scala 226:16]
  assign io_raddr2 = csr_write[0] ? 5'h11 : inst[24:20]; // @[IDU.scala 225:15]
  assign io_to_es_pc = ds_pc; // @[IDU.scala 525:17]
  assign io_ALUop = {{25'd0}, _ALUop_T_176}; // @[IDU.scala 310:11 64:21]
  assign io_src1 = csr_write[0] ? csr_reg_io_rdata : src1; // @[IDU.scala 514:19]
  assign io_src2 = src2_is_imm ? imm : rdata2; // @[IDU.scala 471:16]
  assign io_rf_dst = inst[11:7]; // @[IDU.scala 227:15]
  assign io_store_data = _inst_type_T_11 ? rdata2 : {{32'd0}, _io_store_data_T_13}; // @[Lookup.scala 34:39]
  assign io_ctrl_sign_reg_write = _ALUop_T_3 ? 1'h0 : _reg_write_T_40; // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Writemem_en = 32'h44 == inst_type; // @[Mux.scala 81:61]
  assign io_ctrl_sign_Readmem_en = _inst_type_T_25 | (_inst_type_T_15 | (_inst_type_T_113 | (_inst_type_T_77 | (
    _inst_type_T_79 | (_inst_type_T_115 | _inst_type_T_33))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Wmask = _inst_type_T_11 ? 8'hff : {{4'd0}, _Wmask_T_10}; // @[Lookup.scala 34:39]
  assign io_load_type = _inst_type_T_15 ? 3'h1 : _load_type_T_19; // @[Lookup.scala 34:39]
  assign io_ds_valid = ds_valid; // @[IDU.scala 527:17]
  assign csr_reg_clock = clock;
  assign csr_reg_io_wen1 = csr_write[0] & ds_valid; // @[IDU.scala 462:38]
  assign csr_reg_io_wen2 = csr_write[1] & ds_valid; // @[IDU.scala 465:38]
  assign csr_reg_io_waddr1 = _conflict_es_rs2_T_5 ? 2'h1 : _T_18; // @[IDU.scala 463:22]
  assign csr_reg_io_wdata1 = _conflict_es_rs2_T_5 ? ds_pc : _T_22; // @[IDU.scala 464:22]
  assign csr_reg_io_wdata2 = conflict_es_rs2 ? io_es_fwd_res : _rdata2_T_1; // @[IDU.scala 498:18]
  assign csr_reg_io_raddr = csr_write[1] ? 2'h0 : _T_11; // @[IDU.scala 461:21]
  always @(posedge clock) begin
    if (reset) begin // @[IDU.scala 111:27]
      ds_valid <= 1'h0; // @[IDU.scala 111:27]
    end else if (br_taken & ds_allowin & io_fs_to_ds_valid & _T_1) begin // @[IDU.scala 141:74]
      ds_valid <= 1'h0; // @[IDU.scala 142:18]
    end else if (ds_allowin) begin // @[IDU.scala 143:27]
      ds_valid <= io_fs_to_ds_valid; // @[IDU.scala 144:18]
    end
    if (reset) begin // @[IDU.scala 115:24]
      ds_pc <= 64'h0; // @[IDU.scala 115:24]
    end else if (io_fs_to_ds_valid & ds_allowin) begin // @[IDU.scala 146:40]
      ds_pc <= io_pc; // @[IDU.scala 147:15]
    end
    if (reset) begin // @[IDU.scala 117:23]
      inst <= 32'h0; // @[IDU.scala 117:23]
    end else if (io_fs_to_ds_valid & ds_allowin) begin // @[IDU.scala 146:40]
      inst <= io_from_fs_inst; // @[IDU.scala 148:14]
    end
    if (reset) begin // @[IDU.scala 121:34]
      br_taken_cancel <= 1'h0; // @[IDU.scala 121:34]
    end else if (ds_allowin & io_fs_to_ds_valid) begin // @[IDU.scala 132:42]
      br_taken_cancel <= _T_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ds_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  ds_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  br_taken_cancel = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module partial_product(
  input  [2:0]  io_y,
  input  [63:0] io_x,
  output        io_c,
  output [63:0] io_p
);
  wire [64:0] _io_p_T = {io_x, 1'h0}; // @[Mul.scala 24:18]
  wire [64:0] _io_p_T_2 = ~_io_p_T; // @[Mul.scala 25:12]
  wire [63:0] _io_p_T_3 = ~io_x; // @[Mul.scala 26:12]
  wire [63:0] _io_p_T_6 = 3'h1 == io_y ? io_x : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_p_T_8 = 3'h2 == io_y ? io_x : _io_p_T_6; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_10 = 3'h3 == io_y ? _io_p_T : {{1'd0}, _io_p_T_8}; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_12 = 3'h4 == io_y ? _io_p_T_2 : _io_p_T_10; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_14 = 3'h5 == io_y ? {{1'd0}, _io_p_T_3} : _io_p_T_12; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_16 = 3'h6 == io_y ? {{1'd0}, _io_p_T_3} : _io_p_T_14; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_18 = 3'h7 == io_y ? 65'h0 : _io_p_T_16; // @[Mux.scala 81:58]
  assign io_c = 3'h6 == io_y | (3'h5 == io_y | 3'h4 == io_y); // @[Mux.scala 81:58]
  assign io_p = _io_p_T_18[63:0]; // @[Mul.scala 20:8]
endmodule
module Mul(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input         io_mulw,
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output        io_out_valid,
  output [31:0] io_result_hi,
  output [31:0] io_result_lo
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [95:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] booth_partial_io_y; // @[Mul.scala 91:43]
  wire [63:0] booth_partial_io_x; // @[Mul.scala 91:43]
  wire  booth_partial_io_c; // @[Mul.scala 91:43]
  wire [63:0] booth_partial_io_p; // @[Mul.scala 91:43]
  wire  sign = io_multiplicand[63] ^ io_multiplier[63]; // @[Mul.scala 51:33]
  reg [63:0] res; // @[Mul.scala 53:22]
  reg [1:0] state; // @[Mul.scala 55:24]
  reg [127:0] src1; // @[Mul.scala 57:23]
  reg [64:0] src2; // @[Mul.scala 58:23]
  wire [31:0] _src1_32_T_2 = io_multiplicand[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _src1_32_T_4 = {_src1_32_T_2,io_multiplicand[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] src1_32 = io_mulw ? _src1_32_T_4 : io_multiplicand; // @[Mul.scala 65:19]
  wire [31:0] _src2_32_T_2 = io_multiplier[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _src2_32_T_4 = {_src2_32_T_2,io_multiplier[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] src2_32 = io_mulw ? _src2_32_T_4 : io_multiplier; // @[Mul.scala 66:19]
  wire [63:0] _real_cand_T_5 = src1_32[63] ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 74:12]
  wire [127:0] real_cand = {_real_cand_T_5,src1_32}; // @[Cat.scala 31:58]
  wire [64:0] _real_er_T = {src2_32,1'h0}; // @[Cat.scala 31:58]
  wire [127:0] _GEN_1 = io_mul_valid ? real_cand : src1; // @[Mul.scala 77:44 79:22 57:23]
  wire [63:0] real_er = _real_er_T[63:0]; // @[Mul.scala 61:23 69:13]
  wire [63:0] _res_T_1 = res + booth_partial_io_p; // @[Mul.scala 95:32]
  wire [63:0] _GEN_25 = {{63'd0}, booth_partial_io_c}; // @[Mul.scala 95:53]
  wire [63:0] _res_T_3 = _res_T_1 + _GEN_25; // @[Mul.scala 95:53]
  wire [129:0] _src1_T = {src1, 2'h0}; // @[Mul.scala 97:34]
  wire [63:0] _GEN_3 = src2 != 65'h0 ? _res_T_3 : res; // @[Mul.scala 53:22 94:33 95:25]
  wire [129:0] _GEN_5 = src2 != 65'h0 ? _src1_T : {{2'd0}, src1}; // @[Mul.scala 57:23 94:33 97:26]
  wire [63:0] _GEN_14 = 2'h1 == state ? _GEN_3 : res; // @[Mul.scala 71:18 53:22]
  wire [129:0] _GEN_16 = 2'h1 == state ? _GEN_5 : {{2'd0}, src1}; // @[Mul.scala 71:18 57:23]
  wire [129:0] _GEN_18 = 2'h0 == state ? {{2'd0}, _GEN_1} : _GEN_16; // @[Mul.scala 71:18]
  wire [63:0] _GEN_20 = 2'h0 == state ? res : _GEN_14; // @[Mul.scala 71:18 53:22]
  wire  _T_8 = state == 2'h2; // @[Mul.scala 132:21]
  wire [31:0] _io_result_hi_T_1 = {sign,res[62:32]}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_27 = state == 2'h2 ? _io_result_hi_T_1 : 32'h0; // @[Mul.scala 132:35 149:22]
  wire [31:0] _GEN_28 = state == 2'h2 ? res[31:0] : 32'h0; // @[Mul.scala 132:35 150:22]
  wire  _GEN_31 = state == 2'h1 ? 1'h0 : _T_8; // @[Mul.scala 127:33 129:22]
  wire [31:0] _GEN_32 = state == 2'h1 ? 32'h0 : _GEN_27; // @[Mul.scala 127:33 130:22]
  wire [31:0] _GEN_33 = state == 2'h1 ? 32'h0 : _GEN_28; // @[Mul.scala 127:33 131:22]
  wire [129:0] _GEN_30 = reset ? 130'h0 : _GEN_18; // @[Mul.scala 57:{23,23}]
  partial_product booth_partial ( // @[Mul.scala 91:43]
    .io_y(booth_partial_io_y),
    .io_x(booth_partial_io_x),
    .io_c(booth_partial_io_c),
    .io_p(booth_partial_io_p)
  );
  assign io_out_valid = state == 2'h0 ? 1'h0 : _GEN_31; // @[Mul.scala 122:23 124:22]
  assign io_result_hi = state == 2'h0 ? 32'h0 : _GEN_32; // @[Mul.scala 122:23 125:22]
  assign io_result_lo = state == 2'h0 ? 32'h0 : _GEN_33; // @[Mul.scala 122:23 126:22]
  assign booth_partial_io_y = src2[2:0]; // @[Mul.scala 92:43]
  assign booth_partial_io_x = src1[63:0]; // @[Mul.scala 93:36]
  always @(posedge clock) begin
    if (reset) begin // @[Mul.scala 53:22]
      res <= 64'h0; // @[Mul.scala 53:22]
    end else if (state == 2'h0) begin // @[Mul.scala 122:23]
      res <= _GEN_20;
    end else if (state == 2'h1) begin // @[Mul.scala 127:33]
      res <= _GEN_20;
    end else if (state == 2'h2) begin // @[Mul.scala 132:35]
      res <= 64'h0;
    end else begin
      res <= _GEN_20;
    end
    if (reset) begin // @[Mul.scala 55:24]
      state <= 2'h0; // @[Mul.scala 55:24]
    end else if (2'h0 == state) begin // @[Mul.scala 71:18]
      if (io_mul_valid) begin // @[Mul.scala 77:44]
        state <= 2'h1; // @[Mul.scala 78:23]
      end
    end else if (2'h1 == state) begin // @[Mul.scala 71:18]
      if (!(src2 != 65'h0)) begin // @[Mul.scala 94:33]
        state <= 2'h2; // @[Mul.scala 99:27]
      end
    end else if (2'h2 == state) begin // @[Mul.scala 71:18]
      state <= 2'h0;
    end
    src1 <= _GEN_30[127:0]; // @[Mul.scala 57:{23,23}]
    if (reset) begin // @[Mul.scala 58:23]
      src2 <= 65'h0; // @[Mul.scala 58:23]
    end else if (2'h0 == state) begin // @[Mul.scala 71:18]
      if (io_mul_valid) begin // @[Mul.scala 77:44]
        src2 <= {{1'd0}, real_er}; // @[Mul.scala 80:22]
      end
    end else if (2'h1 == state) begin // @[Mul.scala 71:18]
      if (src2 != 65'h0) begin // @[Mul.scala 94:33]
        src2 <= {{2'd0}, src2[64:2]}; // @[Mul.scala 96:26]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  res = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  _RAND_2 = {4{`RANDOM}};
  src1 = _RAND_2[127:0];
  _RAND_3 = {3{`RANDOM}};
  src2 = _RAND_3[64:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Div(
  input         clock,
  input         reset,
  input  [63:0] io_dividend,
  input  [63:0] io_divisor,
  input         io_div_valid,
  input         io_divw,
  input         io_div_signed,
  output        io_out_valid,
  output [63:0] io_quotient,
  output [63:0] io_remainder
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  dend_neg = io_divw ? io_dividend[31] : io_dividend[63]; // @[Div.scala 25:20]
  wire  sor_neg = io_divw ? io_divisor[31] : io_divisor[63]; // @[Div.scala 26:19]
  wire  quotient_neg = dend_neg & ~sor_neg | ~dend_neg & sor_neg; // @[Div.scala 27:43]
  wire [31:0] _src1_32_s_T_2 = io_dividend[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _src1_32_s_T_4 = {_src1_32_s_T_2,io_dividend[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] src1_32_s = io_divw ? _src1_32_s_T_4 : io_dividend; // @[Div.scala 35:21]
  wire [31:0] _src2_32_s_T_2 = io_divisor[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _src2_32_s_T_4 = {_src2_32_s_T_2,io_divisor[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] src2_32_s = io_divw ? _src2_32_s_T_4 : io_divisor; // @[Div.scala 36:21]
  wire [63:0] src1_32 = io_divw ? {{32'd0}, io_dividend[31:0]} : io_dividend; // @[Div.scala 37:19]
  wire [63:0] src2_32 = io_divw ? {{32'd0}, io_divisor[31:0]} : io_divisor; // @[Div.scala 38:19]
  wire [63:0] _real_cand_T_2 = ~src1_32_s; // @[Div.scala 42:61]
  wire [63:0] _real_cand_T_4 = _real_cand_T_2 + 64'h1; // @[Div.scala 42:71]
  wire [63:0] _real_cand_T_5 = dend_neg ? _real_cand_T_4 : src1_32_s; // @[Div.scala 42:45]
  wire [63:0] real_cand = io_div_signed ? _real_cand_T_5 : src1_32; // @[Div.scala 42:21]
  wire [63:0] _real_er_T_2 = ~src2_32_s; // @[Div.scala 43:58]
  wire [63:0] _real_er_T_4 = _real_er_T_2 + 64'h1; // @[Div.scala 43:68]
  wire [63:0] _real_er_T_5 = sor_neg ? _real_er_T_4 : src2_32_s; // @[Div.scala 43:43]
  wire [63:0] real_er = io_div_signed ? _real_er_T_5 : src2_32; // @[Div.scala 43:19]
  wire [95:0] _src1_T_1 = {32'h0,real_cand}; // @[Cat.scala 31:58]
  wire [64:0] src2 = {1'h0,real_er}; // @[Cat.scala 31:58]
  reg [127:0] div_cand; // @[Div.scala 50:27]
  reg  div_start; // @[Div.scala 51:28]
  reg [63:0] quotient; // @[Div.scala 53:27]
  reg [31:0] step_num; // @[Div.scala 55:27]
  wire  _GEN_0 = io_div_valid | div_start; // @[Div.scala 62:27 63:23 51:28]
  wire [127:0] src1 = {{32'd0}, _src1_T_1}; // @[Div.scala 45:20 47:10]
  wire [127:0] _GEN_1 = io_div_valid ? src1 : div_cand; // @[Div.scala 62:27 64:22 50:27]
  wire [63:0] _GEN_2 = io_div_valid ? 64'h0 : quotient; // @[Div.scala 62:27 65:22 53:27]
  wire [31:0] _GEN_3 = io_div_valid ? 32'h40 : step_num; // @[Div.scala 62:27 67:22 55:27]
  wire [64:0] sub_res = div_cand[127:63] - src2; // @[Div.scala 75:41]
  wire [64:0] _quotient_T_2 = {quotient, 1'h0}; // @[Div.scala 77:57]
  wire [64:0] _quotient_T_4 = _quotient_T_2 | 65'h1; // @[Div.scala 77:81]
  wire [64:0] _quotient_T_5 = sub_res[64] ? _quotient_T_2 : _quotient_T_4; // @[Div.scala 77:28]
  wire [127:0] update_cand = {sub_res, 63'h0}; // @[Div.scala 78:36]
  wire [127:0] _new_cand_T_2 = div_cand & 128'h7fffffffffffffff; // @[Div.scala 79:68]
  wire [127:0] _new_cand_T_3 = _new_cand_T_2 | update_cand; // @[Div.scala 79:93]
  wire [127:0] new_cand = sub_res[64] ? div_cand : _new_cand_T_3; // @[Div.scala 79:28]
  wire [128:0] _div_cand_T = {new_cand, 1'h0}; // @[Div.scala 80:34]
  wire [31:0] _step_num_T_1 = step_num - 32'h1; // @[Div.scala 81:34]
  wire [63:0] _io_remainder_T_3 = ~div_cand[127:64]; // @[Div.scala 87:77]
  wire [63:0] _io_remainder_T_5 = _io_remainder_T_3 + 64'h1; // @[Div.scala 87:94]
  wire [63:0] _io_remainder_T_7 = dend_neg ? _io_remainder_T_5 : div_cand[127:64]; // @[Div.scala 87:56]
  wire [63:0] _io_remainder_T_9 = io_div_signed ? _io_remainder_T_7 : div_cand[127:64]; // @[Div.scala 87:32]
  wire [63:0] _io_quotient_T_2 = ~quotient; // @[Div.scala 89:75]
  wire [63:0] _io_quotient_T_4 = _io_quotient_T_2 + 64'h1; // @[Div.scala 89:84]
  wire [63:0] _io_quotient_T_5 = quotient_neg ? _io_quotient_T_4 : quotient; // @[Div.scala 89:55]
  wire [63:0] _io_quotient_T_6 = io_div_signed ? _io_quotient_T_5 : quotient; // @[Div.scala 89:31]
  wire [64:0] _GEN_8 = $signed(step_num) > 32'sh0 ? _quotient_T_5 : {{1'd0}, _GEN_2}; // @[Div.scala 71:36 77:22]
  wire [128:0] _GEN_9 = $signed(step_num) > 32'sh0 ? _div_cand_T : {{1'd0}, _GEN_1}; // @[Div.scala 71:36 80:22]
  wire [63:0] _GEN_11 = $signed(step_num) > 32'sh0 ? 64'h0 : _io_remainder_T_9; // @[Div.scala 71:36 82:26 87:26]
  wire  _GEN_12 = $signed(step_num) > 32'sh0 ? 1'h0 : 1'h1; // @[Div.scala 71:36 83:26 88:26]
  wire [63:0] _GEN_13 = $signed(step_num) > 32'sh0 ? 64'h0 : _io_quotient_T_6; // @[Div.scala 71:36 84:25 89:25]
  wire  _GEN_14 = $signed(step_num) > 32'sh0 & _GEN_0; // @[Div.scala 71:36 86:23]
  wire [64:0] _GEN_15 = div_start ? _GEN_8 : {{1'd0}, _GEN_2}; // @[Div.scala 70:20]
  wire [128:0] _GEN_16 = div_start ? _GEN_9 : {{1'd0}, _GEN_1}; // @[Div.scala 70:20]
  wire [128:0] _GEN_22 = reset ? 129'h0 : _GEN_16; // @[Div.scala 50:{27,27}]
  wire [64:0] _GEN_23 = reset ? 65'h0 : _GEN_15; // @[Div.scala 53:{27,27}]
  assign io_out_valid = div_start & _GEN_12; // @[Div.scala 70:20 93:22]
  assign io_quotient = div_start ? _GEN_13 : 64'h0; // @[Div.scala 70:20 94:21]
  assign io_remainder = div_start ? _GEN_11 : 64'h0; // @[Div.scala 70:20 92:22]
  always @(posedge clock) begin
    div_cand <= _GEN_22[127:0]; // @[Div.scala 50:{27,27}]
    if (reset) begin // @[Div.scala 51:28]
      div_start <= 1'h0; // @[Div.scala 51:28]
    end else if (div_start) begin // @[Div.scala 70:20]
      div_start <= _GEN_14;
    end else begin
      div_start <= _GEN_0;
    end
    quotient <= _GEN_23[63:0]; // @[Div.scala 53:{27,27}]
    if (reset) begin // @[Div.scala 55:27]
      step_num <= 32'h0; // @[Div.scala 55:27]
    end else if (div_start) begin // @[Div.scala 70:20]
      if ($signed(step_num) > 32'sh0) begin // @[Div.scala 71:36]
        step_num <= _step_num_T_1; // @[Div.scala 81:22]
      end else begin
        step_num <= _GEN_3;
      end
    end else begin
      step_num <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  div_cand = _RAND_0[127:0];
  _RAND_1 = {1{`RANDOM}};
  div_start = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  quotient = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  step_num = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [63:0] io_src1_value,
  input  [63:0] io_src2_value,
  input  [31:0] io_ALUop,
  input         io_src_valid,
  output        io_alu_busy,
  output [63:0] io_alu_res
);
  wire  Mul_clock; // @[ALU.scala 60:28]
  wire  Mul_reset; // @[ALU.scala 60:28]
  wire  Mul_io_mul_valid; // @[ALU.scala 60:28]
  wire  Mul_io_mulw; // @[ALU.scala 60:28]
  wire [63:0] Mul_io_multiplicand; // @[ALU.scala 60:28]
  wire [63:0] Mul_io_multiplier; // @[ALU.scala 60:28]
  wire  Mul_io_out_valid; // @[ALU.scala 60:28]
  wire [31:0] Mul_io_result_hi; // @[ALU.scala 60:28]
  wire [31:0] Mul_io_result_lo; // @[ALU.scala 60:28]
  wire  Div_clock; // @[ALU.scala 61:28]
  wire  Div_reset; // @[ALU.scala 61:28]
  wire [63:0] Div_io_dividend; // @[ALU.scala 61:28]
  wire [63:0] Div_io_divisor; // @[ALU.scala 61:28]
  wire  Div_io_div_valid; // @[ALU.scala 61:28]
  wire  Div_io_divw; // @[ALU.scala 61:28]
  wire  Div_io_div_signed; // @[ALU.scala 61:28]
  wire  Div_io_out_valid; // @[ALU.scala 61:28]
  wire [63:0] Div_io_quotient; // @[ALU.scala 61:28]
  wire [63:0] Div_io_remainder; // @[ALU.scala 61:28]
  wire  mul_valid = 32'h12 == io_ALUop | 32'h11 == io_ALUop; // @[Mux.scala 81:58]
  wire  div_valid = 32'h32 == io_ALUop | (32'h14 == io_ALUop | (32'h33 == io_ALUop | (32'h34 == io_ALUop | (32'h35 ==
    io_ALUop | (32'h13 == io_ALUop | (32'h30 == io_ALUop | 32'h31 == io_ALUop)))))); // @[Mux.scala 81:58]
  wire [63:0] add_res = io_src1_value + io_src2_value; // @[ALU.scala 77:30]
  wire [63:0] sub_res = io_src1_value - io_src2_value; // @[ALU.scala 78:30]
  wire [63:0] sra_res = $signed(io_src1_value) >>> io_src2_value[5:0]; // @[ALU.scala 79:60]
  wire [63:0] srl_res = io_src1_value >> io_src2_value[5:0]; // @[ALU.scala 80:30]
  wire [126:0] _GEN_0 = {{63'd0}, io_src1_value}; // @[ALU.scala 81:30]
  wire [126:0] sll_res = _GEN_0 << io_src2_value[5:0]; // @[ALU.scala 81:30]
  wire [31:0] _sraw_res_T_1 = io_src1_value[31:0]; // @[ALU.scala 82:43]
  wire [31:0] sraw_res = $signed(_sraw_res_T_1) >>> io_src2_value[4:0]; // @[ALU.scala 82:46]
  wire [31:0] srlw_res = io_src1_value[31:0] >> io_src2_value[4:0]; // @[ALU.scala 83:37]
  wire [62:0] _GEN_1 = {{31'd0}, io_src1_value[31:0]}; // @[ALU.scala 84:37]
  wire [62:0] sllw_res = _GEN_1 << io_src2_value[4:0]; // @[ALU.scala 84:37]
  wire [63:0] or_res = io_src1_value | io_src2_value; // @[ALU.scala 85:29]
  wire [63:0] xor_res = io_src1_value ^ io_src2_value; // @[ALU.scala 86:30]
  wire [63:0] and_res = io_src1_value & io_src2_value; // @[ALU.scala 87:30]
  wire [63:0] mlu_res = {Mul_io_result_hi,Mul_io_result_lo}; // @[Cat.scala 31:58]
  wire [31:0] divw_res = Div_io_quotient[31:0]; // @[ALU.scala 90:39]
  wire [31:0] remw_res = Div_io_remainder[31:0]; // @[ALU.scala 92:40]
  wire [63:0] _alu_res_T_1 = io_src1_value + 64'h4; // @[ALU.scala 115:29]
  wire  _alu_res_T_4 = io_src1_value < io_src2_value; // @[ALU.scala 118:33]
  wire  _alu_res_T_8 = $signed(io_src1_value) < $signed(io_src2_value); // @[ALU.scala 120:41]
  wire [31:0] _alu_res_T_12 = add_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_14 = {_alu_res_T_12,add_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_17 = sub_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_19 = {_alu_res_T_17,sub_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_22 = sllw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_24 = {_alu_res_T_22,sllw_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_27 = sraw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _alu_res_T_28 = $signed(_sraw_res_T_1) >>> io_src2_value[4:0]; // @[ALU.scala 139:55]
  wire [63:0] _alu_res_T_29 = {_alu_res_T_27,_alu_res_T_28}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_32 = srlw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_34 = {_alu_res_T_32,srlw_res}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_37 = Mul_io_result_lo[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_38 = {_alu_res_T_37,Mul_io_result_lo}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_41 = divw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_42 = {_alu_res_T_41,divw_res}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_49 = remw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_50 = {_alu_res_T_49,remw_res}; // @[Cat.scala 31:58]
  wire [63:0] _alu_res_T_56 = 32'hf == io_ALUop ? add_res : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_58 = 32'h4 == io_ALUop ? io_src2_value : _alu_res_T_56; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_60 = 32'h5 == io_ALUop ? _alu_res_T_1 : _alu_res_T_58; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_62 = 32'h6 == io_ALUop ? _alu_res_T_1 : _alu_res_T_60; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_64 = 32'h1e == io_ALUop ? {{63'd0}, _alu_res_T_4} : _alu_res_T_62; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_66 = 32'h1f == io_ALUop ? {{63'd0}, _alu_res_T_8} : _alu_res_T_64; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_68 = 32'hc == io_ALUop ? _alu_res_T_14 : _alu_res_T_66; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_70 = 32'he == io_ALUop ? sub_res : _alu_res_T_68; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_72 = 32'h15 == io_ALUop ? sra_res : _alu_res_T_70; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_74 = 32'hb == io_ALUop ? or_res : _alu_res_T_72; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_76 = 32'h2e == io_ALUop ? xor_res : _alu_res_T_74; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_78 = 32'h8 == io_ALUop ? and_res : _alu_res_T_76; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_80 = 32'hd == io_ALUop ? _alu_res_T_19 : _alu_res_T_78; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_82 = 32'h16 == io_ALUop ? _alu_res_T_24 : _alu_res_T_80; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_84 = 32'h1c == io_ALUop ? _alu_res_T_29 : _alu_res_T_82; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_86 = 32'h1d == io_ALUop ? _alu_res_T_34 : _alu_res_T_84; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_88 = 32'h11 == io_ALUop ? mlu_res : _alu_res_T_86; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_90 = 32'h12 == io_ALUop ? _alu_res_T_38 : _alu_res_T_88; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_92 = 32'h13 == io_ALUop ? _alu_res_T_42 : _alu_res_T_90; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_94 = 32'h30 == io_ALUop ? Div_io_quotient : _alu_res_T_92; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_96 = 32'h31 == io_ALUop ? Div_io_quotient : _alu_res_T_94; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_98 = 32'h35 == io_ALUop ? _alu_res_T_42 : _alu_res_T_96; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_100 = 32'h14 == io_ALUop ? _alu_res_T_50 : _alu_res_T_98; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_102 = 32'h32 == io_ALUop ? _alu_res_T_50 : _alu_res_T_100; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_104 = 32'h33 == io_ALUop ? Div_io_remainder : _alu_res_T_102; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_106 = 32'h34 == io_ALUop ? Div_io_remainder : _alu_res_T_104; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_108 = 32'h37 == io_ALUop ? sll_res : {{63'd0}, _alu_res_T_106}; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_110 = 32'h39 == io_ALUop ? {{63'd0}, sra_res} : _alu_res_T_108; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_112 = 32'h38 == io_ALUop ? {{63'd0}, srl_res} : _alu_res_T_110; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_114 = 32'h3f == io_ALUop ? {{63'd0}, io_src1_value} : _alu_res_T_112; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_116 = 32'h46 == io_ALUop ? {{63'd0}, io_src1_value} : _alu_res_T_114; // @[Mux.scala 81:58]
  wire [126:0] alu_res = 32'h47 == io_ALUop ? {{63'd0}, io_src1_value} : _alu_res_T_116; // @[Mux.scala 81:58]
  Mul Mul ( // @[ALU.scala 60:28]
    .clock(Mul_clock),
    .reset(Mul_reset),
    .io_mul_valid(Mul_io_mul_valid),
    .io_mulw(Mul_io_mulw),
    .io_multiplicand(Mul_io_multiplicand),
    .io_multiplier(Mul_io_multiplier),
    .io_out_valid(Mul_io_out_valid),
    .io_result_hi(Mul_io_result_hi),
    .io_result_lo(Mul_io_result_lo)
  );
  Div Div ( // @[ALU.scala 61:28]
    .clock(Div_clock),
    .reset(Div_reset),
    .io_dividend(Div_io_dividend),
    .io_divisor(Div_io_divisor),
    .io_div_valid(Div_io_div_valid),
    .io_divw(Div_io_divw),
    .io_div_signed(Div_io_div_signed),
    .io_out_valid(Div_io_out_valid),
    .io_quotient(Div_io_quotient),
    .io_remainder(Div_io_remainder)
  );
  assign io_alu_busy = mul_valid ? ~Mul_io_out_valid : div_valid & ~Div_io_out_valid; // @[ALU.scala 161:23]
  assign io_alu_res = alu_res[63:0]; // @[ALU.scala 162:16]
  assign Mul_clock = clock;
  assign Mul_reset = reset;
  assign Mul_io_mul_valid = mul_valid & io_src_valid; // @[ALU.scala 62:39]
  assign Mul_io_mulw = io_ALUop == 32'h12; // @[ALU.scala 45:22]
  assign Mul_io_multiplicand = io_src1_value; // @[ALU.scala 66:29]
  assign Mul_io_multiplier = io_src2_value; // @[ALU.scala 67:27]
  assign Div_clock = clock;
  assign Div_reset = reset;
  assign Div_io_dividend = io_src1_value; // @[ALU.scala 69:25]
  assign Div_io_divisor = io_src2_value; // @[ALU.scala 70:24]
  assign Div_io_div_valid = div_valid & io_src_valid; // @[ALU.scala 71:39]
  assign Div_io_divw = 32'h32 == io_ALUop | (32'h14 == io_ALUop | (32'h35 == io_ALUop | 32'h13 == io_ALUop)); // @[Mux.scala 81:58]
  assign Div_io_div_signed = 32'h14 == io_ALUop | (32'h34 == io_ALUop | (32'h13 == io_ALUop | 32'h31 == io_ALUop)); // @[Mux.scala 81:58]
endmodule
module EXU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_ds_to_es_valid,
  input         io_ms_allowin,
  output        io_es_allowin,
  input  [31:0] io_ALUop,
  input  [63:0] io_src1_value,
  input  [63:0] io_src2_value,
  input  [4:0]  io_rf_dst,
  input  [63:0] io_store_data,
  output        io_es_to_ms_valid,
  input  [2:0]  io_load_type,
  output [63:0] io_to_ms_pc,
  output [63:0] io_to_ms_alures,
  output [63:0] io_to_ms_store_data,
  output        io_to_ms_wen,
  output [7:0]  io_to_ms_wstrb,
  output        io_to_ms_ren,
  output [63:0] io_to_ms_maddr,
  output [4:0]  io_to_ms_rf_dst,
  output        io_to_ms_rf_we,
  output [2:0]  io_to_ms_load_type,
  input         io_ctrl_sign_reg_write,
  input         io_ctrl_sign_Writemem_en,
  input         io_ctrl_sign_Readmem_en,
  input  [7:0]  io_ctrl_sign_Wmask,
  output        io_es_valid,
  output        io_es_rf_we,
  output [4:0]  io_es_rf_dst,
  output        io_es_fwd_ready,
  output [63:0] io_es_fwd_res,
  output        io_es_ld
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  ALU_clock; // @[EXU.scala 40:21]
  wire  ALU_reset; // @[EXU.scala 40:21]
  wire [63:0] ALU_io_src1_value; // @[EXU.scala 40:21]
  wire [63:0] ALU_io_src2_value; // @[EXU.scala 40:21]
  wire [31:0] ALU_io_ALUop; // @[EXU.scala 40:21]
  wire  ALU_io_src_valid; // @[EXU.scala 40:21]
  wire  ALU_io_alu_busy; // @[EXU.scala 40:21]
  wire [63:0] ALU_io_alu_res; // @[EXU.scala 40:21]
  reg [63:0] es_pc; // @[EXU.scala 42:24]
  reg  es_valid; // @[EXU.scala 43:27]
  reg [4:0] es_rd; // @[EXU.scala 47:24]
  reg  es_rf_we; // @[EXU.scala 48:27]
  reg [63:0] src1_value; // @[EXU.scala 50:29]
  reg [63:0] src2_value; // @[EXU.scala 51:29]
  reg [63:0] store_data; // @[EXU.scala 52:29]
  reg [7:0] st_wstrb; // @[EXU.scala 53:27]
  reg  st_we; // @[EXU.scala 54:24]
  reg  ld_we; // @[EXU.scala 55:24]
  reg [31:0] ALUop; // @[EXU.scala 57:24]
  reg [2:0] load_type; // @[EXU.scala 58:28]
  wire  es_ready_go = ~ALU_io_alu_busy; // @[EXU.scala 78:20]
  wire  es_allowin = ~es_valid | es_ready_go & io_ms_allowin; // @[EXU.scala 80:29]
  ALU ALU ( // @[EXU.scala 40:21]
    .clock(ALU_clock),
    .reset(ALU_reset),
    .io_src1_value(ALU_io_src1_value),
    .io_src2_value(ALU_io_src2_value),
    .io_ALUop(ALU_io_ALUop),
    .io_src_valid(ALU_io_src_valid),
    .io_alu_busy(ALU_io_alu_busy),
    .io_alu_res(ALU_io_alu_res)
  );
  assign io_es_allowin = ~es_valid | es_ready_go & io_ms_allowin; // @[EXU.scala 80:29]
  assign io_es_to_ms_valid = es_valid & es_ready_go; // @[EXU.scala 79:32]
  assign io_to_ms_pc = es_pc; // @[EXU.scala 111:17]
  assign io_to_ms_alures = ALU_io_alu_res; // @[EXU.scala 56:23 98:13]
  assign io_to_ms_store_data = store_data; // @[EXU.scala 114:25]
  assign io_to_ms_wen = st_we; // @[EXU.scala 115:18]
  assign io_to_ms_wstrb = st_wstrb; // @[EXU.scala 116:20]
  assign io_to_ms_ren = ld_we; // @[EXU.scala 117:18]
  assign io_to_ms_maddr = ALU_io_alu_res; // @[EXU.scala 56:23 98:13]
  assign io_to_ms_rf_dst = es_rd; // @[EXU.scala 119:21]
  assign io_to_ms_rf_we = es_rf_we; // @[EXU.scala 120:20]
  assign io_to_ms_load_type = load_type; // @[EXU.scala 124:24]
  assign io_es_valid = es_valid; // @[EXU.scala 121:17]
  assign io_es_rf_we = es_rf_we; // @[EXU.scala 123:17]
  assign io_es_rf_dst = es_rd; // @[EXU.scala 122:18]
  assign io_es_fwd_ready = es_valid & es_ready_go; // @[EXU.scala 79:32]
  assign io_es_fwd_res = ALU_io_alu_res; // @[EXU.scala 56:23 98:13]
  assign io_es_ld = ld_we & es_valid; // @[EXU.scala 127:23]
  assign ALU_clock = clock;
  assign ALU_reset = reset;
  assign ALU_io_src1_value = ALUop == 32'h6 ? es_pc : src1_value; // @[EXU.scala 94:26]
  assign ALU_io_src2_value = src2_value; // @[EXU.scala 95:20]
  assign ALU_io_ALUop = ALUop; // @[EXU.scala 96:15]
  assign ALU_io_src_valid = es_valid; // @[EXU.scala 97:19]
  always @(posedge clock) begin
    if (reset) begin // @[EXU.scala 42:24]
      es_pc <= 64'h0; // @[EXU.scala 42:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      es_pc <= io_pc; // @[EXU.scala 64:15]
    end
    if (reset) begin // @[EXU.scala 43:27]
      es_valid <= 1'h0; // @[EXU.scala 43:27]
    end else if (es_allowin) begin // @[EXU.scala 60:21]
      es_valid <= io_ds_to_es_valid; // @[EXU.scala 61:18]
    end
    if (reset) begin // @[EXU.scala 47:24]
      es_rd <= 5'h0; // @[EXU.scala 47:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      es_rd <= io_rf_dst; // @[EXU.scala 69:15]
    end
    if (reset) begin // @[EXU.scala 48:27]
      es_rf_we <= 1'h0; // @[EXU.scala 48:27]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      es_rf_we <= io_ctrl_sign_reg_write; // @[EXU.scala 65:18]
    end
    if (reset) begin // @[EXU.scala 50:29]
      src1_value <= 64'h0; // @[EXU.scala 50:29]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      src1_value <= io_src1_value; // @[EXU.scala 67:20]
    end
    if (reset) begin // @[EXU.scala 51:29]
      src2_value <= 64'h0; // @[EXU.scala 51:29]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      src2_value <= io_src2_value; // @[EXU.scala 68:20]
    end
    if (reset) begin // @[EXU.scala 52:29]
      store_data <= 64'h0; // @[EXU.scala 52:29]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      store_data <= io_store_data; // @[EXU.scala 70:20]
    end
    if (reset) begin // @[EXU.scala 53:27]
      st_wstrb <= 8'h0; // @[EXU.scala 53:27]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      st_wstrb <= io_ctrl_sign_Wmask; // @[EXU.scala 71:18]
    end
    if (reset) begin // @[EXU.scala 54:24]
      st_we <= 1'h0; // @[EXU.scala 54:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      st_we <= io_ctrl_sign_Writemem_en; // @[EXU.scala 72:15]
    end
    if (reset) begin // @[EXU.scala 55:24]
      ld_we <= 1'h0; // @[EXU.scala 55:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      ld_we <= io_ctrl_sign_Readmem_en; // @[EXU.scala 73:15]
    end
    if (reset) begin // @[EXU.scala 57:24]
      ALUop <= 32'h0; // @[EXU.scala 57:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      ALUop <= io_ALUop; // @[EXU.scala 74:15]
    end
    if (reset) begin // @[EXU.scala 58:28]
      load_type <= 3'h0; // @[EXU.scala 58:28]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      load_type <= io_load_type; // @[EXU.scala 75:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  es_pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  es_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  es_rd = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  es_rf_we = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  src1_value = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  src2_value = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  store_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  st_wstrb = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  st_we = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ld_we = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ALUop = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  load_type = _RAND_11[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_es_to_ms_valid,
  output        io_ms_allowin,
  input         io_rf_we,
  input  [4:0]  io_rf_dst,
  input  [63:0] io_alu_res,
  input  [63:0] io_store_data,
  input  [2:0]  io_load_type,
  input         io_wen,
  input  [7:0]  io_wstrb,
  input         io_ren,
  input  [63:0] io_maddr,
  output [63:0] io_to_ws_pc,
  output [63:0] io_ms_final_res,
  output        io_ms_to_ws_valid,
  output        io_to_ws_rf_we,
  output [4:0]  io_to_ws_rf_dst,
  output        io_ms_valid,
  output        io_ms_rf_we,
  output [4:0]  io_ms_rf_dst,
  output        io_ms_fwd_ready,
  output [63:0] io_ms_fwd_res,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_wready,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [63:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg  ms_valid; // @[LSU.scala 36:27]
  reg [63:0] ms_pc; // @[LSU.scala 37:24]
  reg  ms_ready_go; // @[LSU.scala 39:30]
  reg  ms_rf_we; // @[LSU.scala 41:27]
  reg [4:0] ms_rf_dst; // @[LSU.scala 42:28]
  reg [63:0] ms_res; // @[LSU.scala 43:25]
  reg [63:0] store_data; // @[LSU.scala 45:29]
  reg  wen; // @[LSU.scala 46:22]
  reg [7:0] wstrb; // @[LSU.scala 47:24]
  reg  ren; // @[LSU.scala 48:22]
  reg [63:0] maddr; // @[LSU.scala 49:24]
  reg [2:0] load_type; // @[LSU.scala 50:28]
  wire  ms_allowin = ~ms_valid | ms_ready_go; // @[LSU.scala 71:29]
  wire  _GEN_8 = io_es_to_ms_valid & ms_allowin ? io_ren : ren; // @[LSU.scala 56:40 64:13 48:22]
  wire  _GEN_11 = io_es_to_ms_valid & ms_allowin ? ~(io_wen | io_ren) : ms_ready_go; // @[LSU.scala 56:40 67:21 39:30]
  reg [63:0] mem_rdata; // @[LSU.scala 75:28]
  wire  _GEN_14 = ms_valid & ren & io_axi_in_rvalid | _GEN_11; // @[LSU.scala 80:52 83:21]
  wire  _GEN_16 = ms_valid & wen & io_axi_in_wready | _GEN_14; // @[LSU.scala 77:46 79:21]
  wire [31:0] _rdata_T_2 = mem_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rdata_T_4 = {_rdata_T_2,mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdata_T_7 = {56'h0,mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdata_T_10 = {32'h0,mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [47:0] _rdata_T_13 = mem_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rdata_T_15 = {_rdata_T_13,mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [55:0] _rdata_T_18 = mem_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rdata_T_20 = {_rdata_T_18,mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdata_T_23 = {48'h0,mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdata_T_25 = 3'h1 == load_type ? _rdata_T_4 : mem_rdata; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_27 = 3'h2 == load_type ? mem_rdata : _rdata_T_25; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_29 = 3'h3 == load_type ? _rdata_T_7 : _rdata_T_27; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_31 = 3'h4 == load_type ? _rdata_T_10 : _rdata_T_29; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_33 = 3'h5 == load_type ? _rdata_T_15 : _rdata_T_31; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_35 = 3'h6 == load_type ? _rdata_T_20 : _rdata_T_33; // @[Mux.scala 81:58]
  wire [63:0] rdata = 3'h7 == load_type ? _rdata_T_23 : _rdata_T_35; // @[Mux.scala 81:58]
  wire  _io_ms_final_res_T = load_type != 3'h0; // @[LSU.scala 114:37]
  assign io_ms_allowin = ~ms_valid | ms_ready_go; // @[LSU.scala 71:29]
  assign io_to_ws_pc = ms_pc; // @[LSU.scala 118:17]
  assign io_ms_final_res = load_type != 3'h0 ? rdata : ms_res; // @[LSU.scala 114:27]
  assign io_ms_to_ws_valid = ms_valid & ms_ready_go; // @[LSU.scala 72:32]
  assign io_to_ws_rf_we = ms_rf_we; // @[LSU.scala 117:20]
  assign io_to_ws_rf_dst = ms_rf_dst; // @[LSU.scala 116:21]
  assign io_ms_valid = ms_valid; // @[LSU.scala 120:17]
  assign io_ms_rf_we = ms_rf_we & ms_valid; // @[LSU.scala 122:28]
  assign io_ms_rf_dst = ms_rf_dst; // @[LSU.scala 121:18]
  assign io_ms_fwd_ready = ms_valid & ms_ready_go; // @[LSU.scala 72:32]
  assign io_ms_fwd_res = _io_ms_final_res_T ? rdata : ms_res; // @[LSU.scala 125:25]
  assign io_axi_out_araddr = maddr[31:0]; // @[LSU.scala 87:23]
  assign io_axi_out_arvalid = ren & ms_valid; // @[LSU.scala 88:31]
  assign io_axi_out_awaddr = maddr[31:0]; // @[LSU.scala 93:23]
  assign io_axi_out_awvalid = wen & ms_valid; // @[LSU.scala 94:31]
  assign io_axi_out_wdata = store_data; // @[LSU.scala 98:22]
  assign io_axi_out_wstrb = wstrb; // @[LSU.scala 99:22]
  assign io_axi_out_wvalid = wen; // @[LSU.scala 101:23]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 36:27]
      ms_valid <= 1'h0; // @[LSU.scala 36:27]
    end else if (ms_allowin) begin // @[LSU.scala 53:21]
      ms_valid <= io_es_to_ms_valid; // @[LSU.scala 54:18]
    end
    if (reset) begin // @[LSU.scala 37:24]
      ms_pc <= 64'h0; // @[LSU.scala 37:24]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      ms_pc <= io_pc; // @[LSU.scala 57:15]
    end
    ms_ready_go <= reset | _GEN_16; // @[LSU.scala 39:{30,30}]
    if (reset) begin // @[LSU.scala 41:27]
      ms_rf_we <= 1'h0; // @[LSU.scala 41:27]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      ms_rf_we <= io_rf_we; // @[LSU.scala 58:18]
    end
    if (reset) begin // @[LSU.scala 42:28]
      ms_rf_dst <= 5'h0; // @[LSU.scala 42:28]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      ms_rf_dst <= io_rf_dst; // @[LSU.scala 59:19]
    end
    if (reset) begin // @[LSU.scala 43:25]
      ms_res <= 64'h0; // @[LSU.scala 43:25]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      ms_res <= io_alu_res; // @[LSU.scala 60:16]
    end
    if (reset) begin // @[LSU.scala 45:29]
      store_data <= 64'h0; // @[LSU.scala 45:29]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      store_data <= io_store_data; // @[LSU.scala 61:20]
    end
    if (reset) begin // @[LSU.scala 46:22]
      wen <= 1'h0; // @[LSU.scala 46:22]
    end else if (ms_valid & wen & io_axi_in_wready) begin // @[LSU.scala 77:46]
      wen <= 1'h0; // @[LSU.scala 78:13]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      wen <= io_wen; // @[LSU.scala 62:13]
    end
    if (reset) begin // @[LSU.scala 47:24]
      wstrb <= 8'h0; // @[LSU.scala 47:24]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      wstrb <= io_wstrb; // @[LSU.scala 63:15]
    end
    if (reset) begin // @[LSU.scala 48:22]
      ren <= 1'h0; // @[LSU.scala 48:22]
    end else if (ms_valid & wen & io_axi_in_wready) begin // @[LSU.scala 77:46]
      ren <= _GEN_8;
    end else if (ms_valid & ren & io_axi_in_rvalid) begin // @[LSU.scala 80:52]
      ren <= 1'h0; // @[LSU.scala 82:13]
    end else begin
      ren <= _GEN_8;
    end
    if (reset) begin // @[LSU.scala 49:24]
      maddr <= 64'h0; // @[LSU.scala 49:24]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      maddr <= io_maddr; // @[LSU.scala 65:15]
    end
    if (reset) begin // @[LSU.scala 50:28]
      load_type <= 3'h0; // @[LSU.scala 50:28]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      load_type <= io_load_type; // @[LSU.scala 66:19]
    end
    if (reset) begin // @[LSU.scala 75:28]
      mem_rdata <= 64'h0; // @[LSU.scala 75:28]
    end else if (!(ms_valid & wen & io_axi_in_wready)) begin // @[LSU.scala 77:46]
      if (ms_valid & ren & io_axi_in_rvalid) begin // @[LSU.scala 80:52]
        mem_rdata <= io_axi_in_rdata; // @[LSU.scala 81:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ms_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  ms_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  ms_ready_go = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ms_rf_we = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ms_rf_dst = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  ms_res = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  store_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  wen = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wstrb = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  ren = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  maddr = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  load_type = _RAND_11[2:0];
  _RAND_12 = {2{`RANDOM}};
  mem_rdata = _RAND_12[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_ms_to_ws_valid,
  input  [63:0] io_ms_final_res,
  input         io_rf_we,
  input  [4:0]  io_rf_dst,
  output        io_we,
  output [4:0]  io_waddr,
  output [63:0] io_wdata,
  output        io_ws_valid,
  output        io_ws_rf_we,
  output [4:0]  io_ws_rf_dst,
  output [63:0] io_ws_fwd_res,
  output [63:0] io_ws_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  ws_valid; // @[WBU.scala 25:27]
  reg [63:0] ws_pc; // @[WBU.scala 26:24]
  reg  ws_rf_we; // @[WBU.scala 30:27]
  reg [4:0] ws_rf_dst; // @[WBU.scala 31:28]
  reg [63:0] ws_res; // @[WBU.scala 32:25]
  assign io_we = ws_rf_we & ws_valid; // @[WBU.scala 61:22]
  assign io_waddr = ws_rf_dst; // @[WBU.scala 62:14]
  assign io_wdata = ws_res; // @[WBU.scala 63:14]
  assign io_ws_valid = ws_valid; // @[WBU.scala 64:17]
  assign io_ws_rf_we = ws_rf_we; // @[WBU.scala 66:17]
  assign io_ws_rf_dst = ws_rf_dst; // @[WBU.scala 65:18]
  assign io_ws_fwd_res = ws_res; // @[WBU.scala 68:19]
  assign io_ws_pc = ws_pc; // @[WBU.scala 69:14]
  always @(posedge clock) begin
    if (reset) begin // @[WBU.scala 25:27]
      ws_valid <= 1'h0; // @[WBU.scala 25:27]
    end else begin
      ws_valid <= io_ms_to_ws_valid;
    end
    if (reset) begin // @[WBU.scala 26:24]
      ws_pc <= 64'h0; // @[WBU.scala 26:24]
    end else if (io_ms_to_ws_valid) begin // @[WBU.scala 43:40]
      ws_pc <= io_pc; // @[WBU.scala 44:15]
    end
    if (reset) begin // @[WBU.scala 30:27]
      ws_rf_we <= 1'h0; // @[WBU.scala 30:27]
    end else if (io_ms_to_ws_valid) begin // @[WBU.scala 43:40]
      ws_rf_we <= io_rf_we; // @[WBU.scala 45:18]
    end
    if (reset) begin // @[WBU.scala 31:28]
      ws_rf_dst <= 5'h0; // @[WBU.scala 31:28]
    end else if (io_ms_to_ws_valid) begin // @[WBU.scala 43:40]
      ws_rf_dst <= io_rf_dst; // @[WBU.scala 46:19]
    end
    if (reset) begin // @[WBU.scala 32:25]
      ws_res <= 64'h0; // @[WBU.scala 32:25]
    end else if (io_ms_to_ws_valid) begin // @[WBU.scala 43:40]
      ws_res <= io_ms_final_res; // @[WBU.scala 47:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ws_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  ws_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  ws_rf_we = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ws_rf_dst = _RAND_3[4:0];
  _RAND_4 = {2{`RANDOM}};
  ws_res = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI_ARBITER(
  input         clock,
  input         reset,
  input  [31:0] io_ifu_axi_in_araddr,
  input  [7:0]  io_ifu_axi_in_arlen,
  input         io_ifu_axi_in_arvalid,
  input         io_ifu_axi_in_rready,
  output [63:0] io_ifu_axi_out_rdata,
  output        io_ifu_axi_out_rlast,
  output        io_ifu_axi_out_rvalid,
  input  [31:0] io_lsu_axi_in_araddr,
  input  [7:0]  io_lsu_axi_in_arlen,
  input         io_lsu_axi_in_arvalid,
  input         io_lsu_axi_in_rready,
  input  [31:0] io_lsu_axi_in_awaddr,
  input  [7:0]  io_lsu_axi_in_awlen,
  input         io_lsu_axi_in_awvalid,
  input  [63:0] io_lsu_axi_in_wdata,
  input  [7:0]  io_lsu_axi_in_wstrb,
  input         io_lsu_axi_in_wvalid,
  input         io_lsu_axi_in_bready,
  output [63:0] io_lsu_axi_out_rdata,
  output        io_lsu_axi_out_rlast,
  output        io_lsu_axi_out_rvalid,
  output        io_lsu_axi_out_wready,
  output        io_lsu_axi_out_bvalid,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rlast,
  input         io_axi_in_rvalid,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output [7:0]  io_axi_out_arlen,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output [7:0]  io_axi_out_awlen,
  output        io_axi_out_awvalid,
  output [63:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[axi_arbiter.scala 18:24]
  wire [1:0] _GEN_0 = io_ifu_axi_in_arvalid ? 2'h1 : state; // @[axi_arbiter.scala 59:46 60:23 18:24]
  wire [31:0] _GEN_1 = io_ifu_axi_in_arvalid ? io_ifu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 59:46 61:28 65:28]
  wire [7:0] _GEN_2 = io_ifu_axi_in_arvalid ? io_ifu_axi_in_arlen : 8'h0; // @[axi_arbiter.scala 59:46 61:28 65:28]
  wire  _GEN_6 = io_ifu_axi_in_arvalid & io_ifu_axi_in_rready; // @[axi_arbiter.scala 59:46 61:28 65:28]
  wire [63:0] _GEN_18 = io_ifu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 59:46 62:32 67:32]
  wire  _GEN_19 = io_ifu_axi_in_arvalid & io_axi_in_rlast; // @[axi_arbiter.scala 59:46 62:32 67:32]
  wire  _GEN_20 = io_ifu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 59:46 62:32 67:32]
  wire [31:0] _GEN_32 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_araddr : _GEN_1; // @[axi_arbiter.scala 54:46 56:28]
  wire [7:0] _GEN_33 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_arlen : _GEN_2; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_36 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_arvalid : io_ifu_axi_in_arvalid; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_37 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_rready : _GEN_6; // @[axi_arbiter.scala 54:46 56:28]
  wire [31:0] _GEN_38 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 54:46 56:28]
  wire [7:0] _GEN_39 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_awlen : 8'h0; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_42 = io_lsu_axi_in_arvalid & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 54:46 56:28]
  wire [63:0] _GEN_43 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wdata : 64'h0; // @[axi_arbiter.scala 54:46 56:28]
  wire [7:0] _GEN_44 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_46 = io_lsu_axi_in_arvalid & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_47 = io_lsu_axi_in_arvalid & io_lsu_axi_in_bready; // @[axi_arbiter.scala 54:46 56:28]
  wire [63:0] _GEN_49 = io_lsu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 54:46 57:32]
  wire  _GEN_50 = io_lsu_axi_in_arvalid & io_axi_in_rlast; // @[axi_arbiter.scala 54:46 57:32]
  wire  _GEN_51 = io_lsu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 54:46 57:32]
  wire  _GEN_53 = io_lsu_axi_in_arvalid & io_axi_in_wready; // @[axi_arbiter.scala 54:46 57:32]
  wire  _GEN_54 = io_lsu_axi_in_arvalid & io_axi_in_bvalid; // @[axi_arbiter.scala 54:46 57:32]
  wire [63:0] _GEN_56 = io_lsu_axi_in_arvalid ? 64'h0 : _GEN_18; // @[axi_arbiter.scala 54:46 58:32]
  wire  _GEN_57 = io_lsu_axi_in_arvalid ? 1'h0 : _GEN_19; // @[axi_arbiter.scala 54:46 58:32]
  wire  _GEN_58 = io_lsu_axi_in_arvalid ? 1'h0 : _GEN_20; // @[axi_arbiter.scala 54:46 58:32]
  wire [31:0] _GEN_63 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_araddr : _GEN_32; // @[axi_arbiter.scala 49:40 51:28]
  wire [7:0] _GEN_64 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_arlen : _GEN_33; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_67 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_arvalid : _GEN_36; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_68 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_rready : _GEN_37; // @[axi_arbiter.scala 49:40 51:28]
  wire [31:0] _GEN_69 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awaddr : _GEN_38; // @[axi_arbiter.scala 49:40 51:28]
  wire [7:0] _GEN_70 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awlen : _GEN_39; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_73 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awvalid : _GEN_42; // @[axi_arbiter.scala 49:40 51:28]
  wire [63:0] _GEN_74 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wdata : _GEN_43; // @[axi_arbiter.scala 49:40 51:28]
  wire [7:0] _GEN_75 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wstrb : _GEN_44; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_77 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wvalid : _GEN_46; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_78 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_bready : _GEN_47; // @[axi_arbiter.scala 49:40 51:28]
  wire [63:0] _GEN_80 = io_lsu_axi_in_awvalid ? io_axi_in_rdata : _GEN_49; // @[axi_arbiter.scala 49:40 52:32]
  wire  _GEN_81 = io_lsu_axi_in_awvalid ? io_axi_in_rlast : _GEN_50; // @[axi_arbiter.scala 49:40 52:32]
  wire  _GEN_82 = io_lsu_axi_in_awvalid ? io_axi_in_rvalid : _GEN_51; // @[axi_arbiter.scala 49:40 52:32]
  wire  _GEN_84 = io_lsu_axi_in_awvalid ? io_axi_in_wready : _GEN_53; // @[axi_arbiter.scala 49:40 52:32]
  wire  _GEN_85 = io_lsu_axi_in_awvalid ? io_axi_in_bvalid : _GEN_54; // @[axi_arbiter.scala 49:40 52:32]
  wire [63:0] _GEN_87 = io_lsu_axi_in_awvalid ? 64'h0 : _GEN_56; // @[axi_arbiter.scala 49:40 53:32]
  wire  _GEN_88 = io_lsu_axi_in_awvalid ? 1'h0 : _GEN_57; // @[axi_arbiter.scala 49:40 53:32]
  wire  _GEN_89 = io_lsu_axi_in_awvalid ? 1'h0 : _GEN_58; // @[axi_arbiter.scala 49:40 53:32]
  wire [1:0] _GEN_94 = io_lsu_axi_out_rvalid & io_lsu_axi_in_rready & io_lsu_axi_out_rlast ? 2'h0 : state; // @[axi_arbiter.scala 82:88 83:23 18:24]
  wire [1:0] _GEN_95 = io_lsu_axi_out_bvalid & io_lsu_axi_in_bready ? 2'h0 : state; // @[axi_arbiter.scala 90:64 91:23 18:24]
  wire [31:0] _GEN_96 = state == 2'h3 ? io_lsu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [7:0] _GEN_97 = state == 2'h3 ? io_lsu_axi_in_arlen : 8'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_100 = state == 2'h3 & io_lsu_axi_in_arvalid; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_101 = state == 2'h3 & io_lsu_axi_in_rready; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [31:0] _GEN_102 = state == 2'h3 ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [7:0] _GEN_103 = state == 2'h3 ? io_lsu_axi_in_awlen : 8'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_106 = state == 2'h3 & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [63:0] _GEN_107 = state == 2'h3 ? io_lsu_axi_in_wdata : 64'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [7:0] _GEN_108 = state == 2'h3 ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_110 = state == 2'h3 & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_111 = state == 2'h3 & io_lsu_axi_in_bready; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [63:0] _GEN_113 = state == 2'h3 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire  _GEN_114 = state == 2'h3 & io_axi_in_rlast; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire  _GEN_115 = state == 2'h3 & io_axi_in_rvalid; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire  _GEN_117 = state == 2'h3 & io_axi_in_wready; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire  _GEN_118 = state == 2'h3 & io_axi_in_bvalid; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire [1:0] _GEN_126 = state == 2'h3 ? _GEN_95 : state; // @[axi_arbiter.scala 18:24 86:39]
  wire [31:0] _GEN_127 = state == 2'h2 ? io_lsu_axi_in_araddr : _GEN_96; // @[axi_arbiter.scala 78:39 79:24]
  wire [7:0] _GEN_128 = state == 2'h2 ? io_lsu_axi_in_arlen : _GEN_97; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_131 = state == 2'h2 ? io_lsu_axi_in_arvalid : _GEN_100; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_132 = state == 2'h2 ? io_lsu_axi_in_rready : _GEN_101; // @[axi_arbiter.scala 78:39 79:24]
  wire [31:0] _GEN_133 = state == 2'h2 ? io_lsu_axi_in_awaddr : _GEN_102; // @[axi_arbiter.scala 78:39 79:24]
  wire [7:0] _GEN_134 = state == 2'h2 ? io_lsu_axi_in_awlen : _GEN_103; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_137 = state == 2'h2 ? io_lsu_axi_in_awvalid : _GEN_106; // @[axi_arbiter.scala 78:39 79:24]
  wire [63:0] _GEN_138 = state == 2'h2 ? io_lsu_axi_in_wdata : _GEN_107; // @[axi_arbiter.scala 78:39 79:24]
  wire [7:0] _GEN_139 = state == 2'h2 ? io_lsu_axi_in_wstrb : _GEN_108; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_141 = state == 2'h2 ? io_lsu_axi_in_wvalid : _GEN_110; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_142 = state == 2'h2 ? io_lsu_axi_in_bready : _GEN_111; // @[axi_arbiter.scala 78:39 79:24]
  wire [63:0] _GEN_144 = state == 2'h2 ? io_axi_in_rdata : _GEN_113; // @[axi_arbiter.scala 78:39 80:28]
  wire  _GEN_145 = state == 2'h2 ? io_axi_in_rlast : _GEN_114; // @[axi_arbiter.scala 78:39 80:28]
  wire  _GEN_146 = state == 2'h2 ? io_axi_in_rvalid : _GEN_115; // @[axi_arbiter.scala 78:39 80:28]
  wire  _GEN_148 = state == 2'h2 ? io_axi_in_wready : _GEN_117; // @[axi_arbiter.scala 78:39 80:28]
  wire  _GEN_149 = state == 2'h2 ? io_axi_in_bvalid : _GEN_118; // @[axi_arbiter.scala 78:39 80:28]
  wire [31:0] _GEN_158 = state == 2'h1 ? io_ifu_axi_in_araddr : _GEN_127; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_159 = state == 2'h1 ? io_ifu_axi_in_arlen : _GEN_128; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_162 = state == 2'h1 ? io_ifu_axi_in_arvalid : _GEN_131; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_163 = state == 2'h1 ? io_ifu_axi_in_rready : _GEN_132; // @[axi_arbiter.scala 70:39 71:24]
  wire [31:0] _GEN_164 = state == 2'h1 ? 32'h0 : _GEN_133; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_165 = state == 2'h1 ? 8'h0 : _GEN_134; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_168 = state == 2'h1 ? 1'h0 : _GEN_137; // @[axi_arbiter.scala 70:39 71:24]
  wire [63:0] _GEN_169 = state == 2'h1 ? 64'h0 : _GEN_138; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_170 = state == 2'h1 ? 8'h0 : _GEN_139; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_172 = state == 2'h1 ? 1'h0 : _GEN_141; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_173 = state == 2'h1 ? 1'h0 : _GEN_142; // @[axi_arbiter.scala 70:39 71:24]
  wire [63:0] _GEN_175 = state == 2'h1 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_176 = state == 2'h1 & io_axi_in_rlast; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_177 = state == 2'h1 & io_axi_in_rvalid; // @[axi_arbiter.scala 70:39 72:28]
  wire [63:0] _GEN_182 = state == 2'h1 ? 64'h0 : _GEN_144; // @[axi_arbiter.scala 70:39 73:28]
  wire  _GEN_183 = state == 2'h1 ? 1'h0 : _GEN_145; // @[axi_arbiter.scala 70:39 73:28]
  wire  _GEN_184 = state == 2'h1 ? 1'h0 : _GEN_146; // @[axi_arbiter.scala 70:39 73:28]
  wire  _GEN_186 = state == 2'h1 ? 1'h0 : _GEN_148; // @[axi_arbiter.scala 70:39 73:28]
  wire  _GEN_187 = state == 2'h1 ? 1'h0 : _GEN_149; // @[axi_arbiter.scala 70:39 73:28]
  assign io_ifu_axi_out_rdata = state == 2'h0 ? _GEN_87 : _GEN_175; // @[axi_arbiter.scala 48:27]
  assign io_ifu_axi_out_rlast = state == 2'h0 ? _GEN_88 : _GEN_176; // @[axi_arbiter.scala 48:27]
  assign io_ifu_axi_out_rvalid = state == 2'h0 ? _GEN_89 : _GEN_177; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_rdata = state == 2'h0 ? _GEN_80 : _GEN_182; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_rlast = state == 2'h0 ? _GEN_81 : _GEN_183; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_rvalid = state == 2'h0 ? _GEN_82 : _GEN_184; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_wready = state == 2'h0 ? _GEN_84 : _GEN_186; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_bvalid = state == 2'h0 ? _GEN_85 : _GEN_187; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_araddr = state == 2'h0 ? _GEN_63 : _GEN_158; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_arlen = state == 2'h0 ? _GEN_64 : _GEN_159; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_arvalid = state == 2'h0 ? _GEN_67 : _GEN_162; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_rready = state == 2'h0 ? _GEN_68 : _GEN_163; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_awaddr = state == 2'h0 ? _GEN_69 : _GEN_164; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_awlen = state == 2'h0 ? _GEN_70 : _GEN_165; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_awvalid = state == 2'h0 ? _GEN_73 : _GEN_168; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_wdata = state == 2'h0 ? _GEN_74 : _GEN_169; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_wstrb = state == 2'h0 ? _GEN_75 : _GEN_170; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_wvalid = state == 2'h0 ? _GEN_77 : _GEN_172; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_bready = state == 2'h0 ? _GEN_78 : _GEN_173; // @[axi_arbiter.scala 48:27]
  always @(posedge clock) begin
    if (reset) begin // @[axi_arbiter.scala 18:24]
      state <= 2'h0; // @[axi_arbiter.scala 18:24]
    end else if (state == 2'h0) begin // @[axi_arbiter.scala 48:27]
      if (io_lsu_axi_in_awvalid) begin // @[axi_arbiter.scala 49:40]
        state <= 2'h3; // @[axi_arbiter.scala 50:23]
      end else if (io_lsu_axi_in_arvalid) begin // @[axi_arbiter.scala 54:46]
        state <= 2'h2; // @[axi_arbiter.scala 55:23]
      end else begin
        state <= _GEN_0;
      end
    end else if (state == 2'h1) begin // @[axi_arbiter.scala 70:39]
      if (io_ifu_axi_out_rvalid & io_ifu_axi_in_rready & io_ifu_axi_out_rlast) begin // @[axi_arbiter.scala 74:88]
        state <= 2'h0; // @[axi_arbiter.scala 75:23]
      end
    end else if (state == 2'h2) begin // @[axi_arbiter.scala 78:39]
      state <= _GEN_94;
    end else begin
      state <= _GEN_126;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module I_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_ifu_araddr,
  input         io_from_ifu_arvalid,
  input         io_from_ifu_rready,
  output [63:0] io_to_ifu_rdata,
  output        io_to_ifu_rlast,
  output        io_to_ifu_rvalid,
  output [31:0] io_to_axi_araddr,
  output [7:0]  io_to_axi_arlen,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rlast,
  input         io_from_axi_rvalid,
  output        io_cache_init,
  input         io_clear_cache
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [511:0] _RAND_2;
  reg [511:0] _RAND_3;
  reg [511:0] _RAND_4;
  reg [511:0] _RAND_5;
  reg [511:0] _RAND_6;
  reg [511:0] _RAND_7;
  reg [511:0] _RAND_8;
  reg [511:0] _RAND_9;
  reg [511:0] _RAND_10;
  reg [511:0] _RAND_11;
  reg [511:0] _RAND_12;
  reg [511:0] _RAND_13;
  reg [511:0] _RAND_14;
  reg [511:0] _RAND_15;
  reg [511:0] _RAND_16;
  reg [511:0] _RAND_17;
  reg [511:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [511:0] _RAND_21;
  reg [511:0] _RAND_22;
  reg [511:0] _RAND_23;
  reg [511:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [511:0] _RAND_26;
  reg [511:0] _RAND_27;
  reg [511:0] _RAND_28;
  reg [511:0] _RAND_29;
  reg [511:0] _RAND_30;
  reg [511:0] _RAND_31;
  reg [511:0] _RAND_32;
  reg [511:0] _RAND_33;
  reg [511:0] _RAND_34;
  reg [511:0] _RAND_35;
  reg [511:0] _RAND_36;
  reg [511:0] _RAND_37;
  reg [511:0] _RAND_38;
  reg [511:0] _RAND_39;
  reg [511:0] _RAND_40;
  reg [511:0] _RAND_41;
  reg [511:0] _RAND_42;
  reg [511:0] _RAND_43;
  reg [511:0] _RAND_44;
  reg [511:0] _RAND_45;
  reg [511:0] _RAND_46;
  reg [511:0] _RAND_47;
  reg [511:0] _RAND_48;
  reg [511:0] _RAND_49;
  reg [511:0] _RAND_50;
  reg [511:0] _RAND_51;
  reg [511:0] _RAND_52;
  reg [511:0] _RAND_53;
  reg [511:0] _RAND_54;
  reg [511:0] _RAND_55;
  reg [511:0] _RAND_56;
  reg [511:0] _RAND_57;
  reg [511:0] _RAND_58;
  reg [511:0] _RAND_59;
  reg [511:0] _RAND_60;
  reg [511:0] _RAND_61;
  reg [511:0] _RAND_62;
  reg [511:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] ram_0_0; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_1; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_2; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_3; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_4; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_5; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_6; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_7; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_8; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_9; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_10; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_11; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_12; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_13; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_14; // @[i_cache.scala 19:24]
  reg [511:0] ram_0_15; // @[i_cache.scala 19:24]
  reg [511:0] ram_1_0; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_1; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_2; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_3; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_4; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_5; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_6; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_7; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_8; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_9; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_10; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_11; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_12; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_13; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_14; // @[i_cache.scala 20:24]
  reg [511:0] ram_1_15; // @[i_cache.scala 20:24]
  reg [511:0] ram_2_0; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_1; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_2; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_3; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_4; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_5; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_6; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_7; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_8; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_9; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_10; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_11; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_12; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_13; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_14; // @[i_cache.scala 21:24]
  reg [511:0] ram_2_15; // @[i_cache.scala 21:24]
  reg [511:0] ram_3_0; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_1; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_2; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_3; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_4; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_5; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_6; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_7; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_8; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_9; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_10; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_11; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_12; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_13; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_14; // @[i_cache.scala 22:24]
  reg [511:0] ram_3_15; // @[i_cache.scala 22:24]
  reg [31:0] tag_0_0; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_1; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_2; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_3; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_4; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_5; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_6; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_7; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_8; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_9; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_10; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_11; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_12; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_13; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_14; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_15; // @[i_cache.scala 23:24]
  reg [31:0] tag_1_0; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_1; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_2; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_3; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_4; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_5; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_6; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_7; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_8; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_9; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_10; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_11; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_12; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_13; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_14; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_15; // @[i_cache.scala 24:24]
  reg [31:0] tag_2_0; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_1; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_2; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_3; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_4; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_5; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_6; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_7; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_8; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_9; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_10; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_11; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_12; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_13; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_14; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_15; // @[i_cache.scala 25:24]
  reg [31:0] tag_3_0; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_1; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_2; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_3; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_4; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_5; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_6; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_7; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_8; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_9; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_10; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_11; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_12; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_13; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_14; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_15; // @[i_cache.scala 26:24]
  reg  valid_0_0; // @[i_cache.scala 27:26]
  reg  valid_0_1; // @[i_cache.scala 27:26]
  reg  valid_0_2; // @[i_cache.scala 27:26]
  reg  valid_0_3; // @[i_cache.scala 27:26]
  reg  valid_0_4; // @[i_cache.scala 27:26]
  reg  valid_0_5; // @[i_cache.scala 27:26]
  reg  valid_0_6; // @[i_cache.scala 27:26]
  reg  valid_0_7; // @[i_cache.scala 27:26]
  reg  valid_0_8; // @[i_cache.scala 27:26]
  reg  valid_0_9; // @[i_cache.scala 27:26]
  reg  valid_0_10; // @[i_cache.scala 27:26]
  reg  valid_0_11; // @[i_cache.scala 27:26]
  reg  valid_0_12; // @[i_cache.scala 27:26]
  reg  valid_0_13; // @[i_cache.scala 27:26]
  reg  valid_0_14; // @[i_cache.scala 27:26]
  reg  valid_0_15; // @[i_cache.scala 27:26]
  reg  valid_1_0; // @[i_cache.scala 28:26]
  reg  valid_1_1; // @[i_cache.scala 28:26]
  reg  valid_1_2; // @[i_cache.scala 28:26]
  reg  valid_1_3; // @[i_cache.scala 28:26]
  reg  valid_1_4; // @[i_cache.scala 28:26]
  reg  valid_1_5; // @[i_cache.scala 28:26]
  reg  valid_1_6; // @[i_cache.scala 28:26]
  reg  valid_1_7; // @[i_cache.scala 28:26]
  reg  valid_1_8; // @[i_cache.scala 28:26]
  reg  valid_1_9; // @[i_cache.scala 28:26]
  reg  valid_1_10; // @[i_cache.scala 28:26]
  reg  valid_1_11; // @[i_cache.scala 28:26]
  reg  valid_1_12; // @[i_cache.scala 28:26]
  reg  valid_1_13; // @[i_cache.scala 28:26]
  reg  valid_1_14; // @[i_cache.scala 28:26]
  reg  valid_1_15; // @[i_cache.scala 28:26]
  reg  valid_2_0; // @[i_cache.scala 29:26]
  reg  valid_2_1; // @[i_cache.scala 29:26]
  reg  valid_2_2; // @[i_cache.scala 29:26]
  reg  valid_2_3; // @[i_cache.scala 29:26]
  reg  valid_2_4; // @[i_cache.scala 29:26]
  reg  valid_2_5; // @[i_cache.scala 29:26]
  reg  valid_2_6; // @[i_cache.scala 29:26]
  reg  valid_2_7; // @[i_cache.scala 29:26]
  reg  valid_2_8; // @[i_cache.scala 29:26]
  reg  valid_2_9; // @[i_cache.scala 29:26]
  reg  valid_2_10; // @[i_cache.scala 29:26]
  reg  valid_2_11; // @[i_cache.scala 29:26]
  reg  valid_2_12; // @[i_cache.scala 29:26]
  reg  valid_2_13; // @[i_cache.scala 29:26]
  reg  valid_2_14; // @[i_cache.scala 29:26]
  reg  valid_2_15; // @[i_cache.scala 29:26]
  reg  valid_3_0; // @[i_cache.scala 30:26]
  reg  valid_3_1; // @[i_cache.scala 30:26]
  reg  valid_3_2; // @[i_cache.scala 30:26]
  reg  valid_3_3; // @[i_cache.scala 30:26]
  reg  valid_3_4; // @[i_cache.scala 30:26]
  reg  valid_3_5; // @[i_cache.scala 30:26]
  reg  valid_3_6; // @[i_cache.scala 30:26]
  reg  valid_3_7; // @[i_cache.scala 30:26]
  reg  valid_3_8; // @[i_cache.scala 30:26]
  reg  valid_3_9; // @[i_cache.scala 30:26]
  reg  valid_3_10; // @[i_cache.scala 30:26]
  reg  valid_3_11; // @[i_cache.scala 30:26]
  reg  valid_3_12; // @[i_cache.scala 30:26]
  reg  valid_3_13; // @[i_cache.scala 30:26]
  reg  valid_3_14; // @[i_cache.scala 30:26]
  reg  valid_3_15; // @[i_cache.scala 30:26]
  reg [63:0] receive_data_0; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_1; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_2; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_3; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_4; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_5; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_6; // @[i_cache.scala 38:31]
  reg [63:0] receive_data_7; // @[i_cache.scala 38:31]
  reg [2:0] receive_num; // @[i_cache.scala 39:30]
  reg [7:0] quene_0; // @[i_cache.scala 40:24]
  reg [7:0] quene_1; // @[i_cache.scala 40:24]
  reg [7:0] quene_2; // @[i_cache.scala 40:24]
  reg [7:0] quene_3; // @[i_cache.scala 40:24]
  reg [7:0] quene_4; // @[i_cache.scala 40:24]
  reg [7:0] quene_5; // @[i_cache.scala 40:24]
  reg [7:0] quene_6; // @[i_cache.scala 40:24]
  reg [7:0] quene_7; // @[i_cache.scala 40:24]
  reg [7:0] quene_8; // @[i_cache.scala 40:24]
  reg [7:0] quene_9; // @[i_cache.scala 40:24]
  reg [7:0] quene_10; // @[i_cache.scala 40:24]
  reg [7:0] quene_11; // @[i_cache.scala 40:24]
  reg [7:0] quene_12; // @[i_cache.scala 40:24]
  reg [7:0] quene_13; // @[i_cache.scala 40:24]
  reg [7:0] quene_14; // @[i_cache.scala 40:24]
  reg [7:0] quene_15; // @[i_cache.scala 40:24]
  wire [5:0] offset = io_from_ifu_araddr[5:0]; // @[i_cache.scala 42:36]
  wire [3:0] index = io_from_ifu_araddr[9:6]; // @[i_cache.scala 43:35]
  wire [21:0] tag = io_from_ifu_araddr[31:10]; // @[i_cache.scala 44:33]
  wire [8:0] shift_bit = {offset, 3'h0}; // @[i_cache.scala 45:28]
  wire [31:0] _GEN_1 = 4'h1 == index ? tag_0_1 : tag_0_0; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_2 = 4'h2 == index ? tag_0_2 : _GEN_1; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_3 = 4'h3 == index ? tag_0_3 : _GEN_2; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_4 = 4'h4 == index ? tag_0_4 : _GEN_3; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_5 = 4'h5 == index ? tag_0_5 : _GEN_4; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_6 = 4'h6 == index ? tag_0_6 : _GEN_5; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_7 = 4'h7 == index ? tag_0_7 : _GEN_6; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_8 = 4'h8 == index ? tag_0_8 : _GEN_7; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_9 = 4'h9 == index ? tag_0_9 : _GEN_8; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_10 = 4'ha == index ? tag_0_10 : _GEN_9; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_11 = 4'hb == index ? tag_0_11 : _GEN_10; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_12 = 4'hc == index ? tag_0_12 : _GEN_11; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_13 = 4'hd == index ? tag_0_13 : _GEN_12; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_14 = 4'he == index ? tag_0_14 : _GEN_13; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_15 = 4'hf == index ? tag_0_15 : _GEN_14; // @[i_cache.scala 47:{31,31}]
  wire [31:0] _GEN_2956 = {{10'd0}, tag}; // @[i_cache.scala 47:31]
  wire  _GEN_17 = 4'h1 == index ? valid_0_1 : valid_0_0; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_18 = 4'h2 == index ? valid_0_2 : _GEN_17; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_19 = 4'h3 == index ? valid_0_3 : _GEN_18; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_20 = 4'h4 == index ? valid_0_4 : _GEN_19; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_21 = 4'h5 == index ? valid_0_5 : _GEN_20; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_22 = 4'h6 == index ? valid_0_6 : _GEN_21; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_23 = 4'h7 == index ? valid_0_7 : _GEN_22; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_24 = 4'h8 == index ? valid_0_8 : _GEN_23; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_25 = 4'h9 == index ? valid_0_9 : _GEN_24; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_26 = 4'ha == index ? valid_0_10 : _GEN_25; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_27 = 4'hb == index ? valid_0_11 : _GEN_26; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_28 = 4'hc == index ? valid_0_12 : _GEN_27; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_29 = 4'hd == index ? valid_0_13 : _GEN_28; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_30 = 4'he == index ? valid_0_14 : _GEN_29; // @[i_cache.scala 47:{57,57}]
  wire  _GEN_31 = 4'hf == index ? valid_0_15 : _GEN_30; // @[i_cache.scala 47:{57,57}]
  wire  way0_hit = _GEN_15 == _GEN_2956 & _GEN_31; // @[i_cache.scala 47:40]
  wire [31:0] _GEN_33 = 4'h1 == index ? tag_1_1 : tag_1_0; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_34 = 4'h2 == index ? tag_1_2 : _GEN_33; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_35 = 4'h3 == index ? tag_1_3 : _GEN_34; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_36 = 4'h4 == index ? tag_1_4 : _GEN_35; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_37 = 4'h5 == index ? tag_1_5 : _GEN_36; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_38 = 4'h6 == index ? tag_1_6 : _GEN_37; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_39 = 4'h7 == index ? tag_1_7 : _GEN_38; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_40 = 4'h8 == index ? tag_1_8 : _GEN_39; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_41 = 4'h9 == index ? tag_1_9 : _GEN_40; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_42 = 4'ha == index ? tag_1_10 : _GEN_41; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_43 = 4'hb == index ? tag_1_11 : _GEN_42; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_44 = 4'hc == index ? tag_1_12 : _GEN_43; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_45 = 4'hd == index ? tag_1_13 : _GEN_44; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_46 = 4'he == index ? tag_1_14 : _GEN_45; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_47 = 4'hf == index ? tag_1_15 : _GEN_46; // @[i_cache.scala 49:{31,31}]
  wire  _GEN_49 = 4'h1 == index ? valid_1_1 : valid_1_0; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_50 = 4'h2 == index ? valid_1_2 : _GEN_49; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_51 = 4'h3 == index ? valid_1_3 : _GEN_50; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_52 = 4'h4 == index ? valid_1_4 : _GEN_51; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_53 = 4'h5 == index ? valid_1_5 : _GEN_52; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_54 = 4'h6 == index ? valid_1_6 : _GEN_53; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_55 = 4'h7 == index ? valid_1_7 : _GEN_54; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_56 = 4'h8 == index ? valid_1_8 : _GEN_55; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_57 = 4'h9 == index ? valid_1_9 : _GEN_56; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_58 = 4'ha == index ? valid_1_10 : _GEN_57; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_59 = 4'hb == index ? valid_1_11 : _GEN_58; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_60 = 4'hc == index ? valid_1_12 : _GEN_59; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_61 = 4'hd == index ? valid_1_13 : _GEN_60; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_62 = 4'he == index ? valid_1_14 : _GEN_61; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_63 = 4'hf == index ? valid_1_15 : _GEN_62; // @[i_cache.scala 49:{57,57}]
  wire  way1_hit = _GEN_47 == _GEN_2956 & _GEN_63; // @[i_cache.scala 49:40]
  wire [31:0] _GEN_65 = 4'h1 == index ? tag_2_1 : tag_2_0; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_66 = 4'h2 == index ? tag_2_2 : _GEN_65; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_67 = 4'h3 == index ? tag_2_3 : _GEN_66; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_68 = 4'h4 == index ? tag_2_4 : _GEN_67; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_69 = 4'h5 == index ? tag_2_5 : _GEN_68; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_70 = 4'h6 == index ? tag_2_6 : _GEN_69; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_71 = 4'h7 == index ? tag_2_7 : _GEN_70; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_72 = 4'h8 == index ? tag_2_8 : _GEN_71; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_73 = 4'h9 == index ? tag_2_9 : _GEN_72; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_74 = 4'ha == index ? tag_2_10 : _GEN_73; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_75 = 4'hb == index ? tag_2_11 : _GEN_74; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_76 = 4'hc == index ? tag_2_12 : _GEN_75; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_77 = 4'hd == index ? tag_2_13 : _GEN_76; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_78 = 4'he == index ? tag_2_14 : _GEN_77; // @[i_cache.scala 50:{31,31}]
  wire [31:0] _GEN_79 = 4'hf == index ? tag_2_15 : _GEN_78; // @[i_cache.scala 50:{31,31}]
  wire  _GEN_81 = 4'h1 == index ? valid_2_1 : valid_2_0; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_82 = 4'h2 == index ? valid_2_2 : _GEN_81; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_83 = 4'h3 == index ? valid_2_3 : _GEN_82; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_84 = 4'h4 == index ? valid_2_4 : _GEN_83; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_85 = 4'h5 == index ? valid_2_5 : _GEN_84; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_86 = 4'h6 == index ? valid_2_6 : _GEN_85; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_87 = 4'h7 == index ? valid_2_7 : _GEN_86; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_88 = 4'h8 == index ? valid_2_8 : _GEN_87; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_89 = 4'h9 == index ? valid_2_9 : _GEN_88; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_90 = 4'ha == index ? valid_2_10 : _GEN_89; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_91 = 4'hb == index ? valid_2_11 : _GEN_90; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_92 = 4'hc == index ? valid_2_12 : _GEN_91; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_93 = 4'hd == index ? valid_2_13 : _GEN_92; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_94 = 4'he == index ? valid_2_14 : _GEN_93; // @[i_cache.scala 50:{57,57}]
  wire  _GEN_95 = 4'hf == index ? valid_2_15 : _GEN_94; // @[i_cache.scala 50:{57,57}]
  wire  way2_hit = _GEN_79 == _GEN_2956 & _GEN_95; // @[i_cache.scala 50:40]
  wire [31:0] _GEN_97 = 4'h1 == index ? tag_3_1 : tag_3_0; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_98 = 4'h2 == index ? tag_3_2 : _GEN_97; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_99 = 4'h3 == index ? tag_3_3 : _GEN_98; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_100 = 4'h4 == index ? tag_3_4 : _GEN_99; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_101 = 4'h5 == index ? tag_3_5 : _GEN_100; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_102 = 4'h6 == index ? tag_3_6 : _GEN_101; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_103 = 4'h7 == index ? tag_3_7 : _GEN_102; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_104 = 4'h8 == index ? tag_3_8 : _GEN_103; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_105 = 4'h9 == index ? tag_3_9 : _GEN_104; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_106 = 4'ha == index ? tag_3_10 : _GEN_105; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_107 = 4'hb == index ? tag_3_11 : _GEN_106; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_108 = 4'hc == index ? tag_3_12 : _GEN_107; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_109 = 4'hd == index ? tag_3_13 : _GEN_108; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_110 = 4'he == index ? tag_3_14 : _GEN_109; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_111 = 4'hf == index ? tag_3_15 : _GEN_110; // @[i_cache.scala 51:{31,31}]
  wire  _GEN_113 = 4'h1 == index ? valid_3_1 : valid_3_0; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_114 = 4'h2 == index ? valid_3_2 : _GEN_113; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_115 = 4'h3 == index ? valid_3_3 : _GEN_114; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_116 = 4'h4 == index ? valid_3_4 : _GEN_115; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_117 = 4'h5 == index ? valid_3_5 : _GEN_116; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_118 = 4'h6 == index ? valid_3_6 : _GEN_117; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_119 = 4'h7 == index ? valid_3_7 : _GEN_118; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_120 = 4'h8 == index ? valid_3_8 : _GEN_119; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_121 = 4'h9 == index ? valid_3_9 : _GEN_120; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_122 = 4'ha == index ? valid_3_10 : _GEN_121; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_123 = 4'hb == index ? valid_3_11 : _GEN_122; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_124 = 4'hc == index ? valid_3_12 : _GEN_123; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_125 = 4'hd == index ? valid_3_13 : _GEN_124; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_126 = 4'he == index ? valid_3_14 : _GEN_125; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_127 = 4'hf == index ? valid_3_15 : _GEN_126; // @[i_cache.scala 51:{57,57}]
  wire  way3_hit = _GEN_111 == _GEN_2956 & _GEN_127; // @[i_cache.scala 51:40]
  wire [2:0] _unuse_way_T_4 = ~_GEN_127 ? 3'h4 : 3'h0; // @[i_cache.scala 52:108]
  wire [2:0] _unuse_way_T_5 = ~_GEN_95 ? 3'h3 : _unuse_way_T_4; // @[i_cache.scala 52:79]
  wire [2:0] _unuse_way_T_6 = ~_GEN_63 ? 3'h2 : _unuse_way_T_5; // @[i_cache.scala 52:50]
  wire [2:0] unuse_way = ~_GEN_31 ? 3'h1 : _unuse_way_T_6; // @[i_cache.scala 52:21]
  reg [2:0] state; // @[i_cache.scala 54:24]
  wire  _T_4 = way0_hit | way1_hit | way2_hit | way3_hit; // @[i_cache.scala 65:46]
  wire [2:0] _GEN_130 = io_from_ifu_rready ? 3'h0 : state; // @[i_cache.scala 54:24 66:41 67:27]
  wire [63:0] _GEN_133 = 3'h0 == receive_num ? io_from_axi_rdata : receive_data_0; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_134 = 3'h1 == receive_num ? io_from_axi_rdata : receive_data_1; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_135 = 3'h2 == receive_num ? io_from_axi_rdata : receive_data_2; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_136 = 3'h3 == receive_num ? io_from_axi_rdata : receive_data_3; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_137 = 3'h4 == receive_num ? io_from_axi_rdata : receive_data_4; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_138 = 3'h5 == receive_num ? io_from_axi_rdata : receive_data_5; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_139 = 3'h6 == receive_num ? io_from_axi_rdata : receive_data_6; // @[i_cache.scala 38:31 76:{43,43}]
  wire [63:0] _GEN_140 = 3'h7 == receive_num ? io_from_axi_rdata : receive_data_7; // @[i_cache.scala 38:31 76:{43,43}]
  wire [2:0] _receive_num_T_1 = receive_num + 3'h1; // @[i_cache.scala 77:44]
  wire [2:0] _GEN_141 = io_from_axi_rlast ? 3'h3 : state; // @[i_cache.scala 54:24 78:40 79:27]
  wire [63:0] _GEN_142 = io_from_axi_rvalid ? _GEN_133 : receive_data_0; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_143 = io_from_axi_rvalid ? _GEN_134 : receive_data_1; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_144 = io_from_axi_rvalid ? _GEN_135 : receive_data_2; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_145 = io_from_axi_rvalid ? _GEN_136 : receive_data_3; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_146 = io_from_axi_rvalid ? _GEN_137 : receive_data_4; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_147 = io_from_axi_rvalid ? _GEN_138 : receive_data_5; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_148 = io_from_axi_rvalid ? _GEN_139 : receive_data_6; // @[i_cache.scala 38:31 75:37]
  wire [63:0] _GEN_149 = io_from_axi_rvalid ? _GEN_140 : receive_data_7; // @[i_cache.scala 38:31 75:37]
  wire [2:0] _GEN_150 = io_from_axi_rvalid ? _receive_num_T_1 : receive_num; // @[i_cache.scala 75:37 77:29 39:30]
  wire [2:0] _GEN_151 = io_from_axi_rvalid ? _GEN_141 : state; // @[i_cache.scala 54:24 75:37]
  wire [511:0] _ram_0_T = {receive_data_7,receive_data_6,receive_data_5,receive_data_4,receive_data_3,receive_data_2,
    receive_data_1,receive_data_0}; // @[Cat.scala 31:58]
  wire [511:0] _GEN_152 = 4'h0 == index ? _ram_0_T : ram_0_0; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_153 = 4'h1 == index ? _ram_0_T : ram_0_1; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_154 = 4'h2 == index ? _ram_0_T : ram_0_2; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_155 = 4'h3 == index ? _ram_0_T : ram_0_3; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_156 = 4'h4 == index ? _ram_0_T : ram_0_4; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_157 = 4'h5 == index ? _ram_0_T : ram_0_5; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_158 = 4'h6 == index ? _ram_0_T : ram_0_6; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_159 = 4'h7 == index ? _ram_0_T : ram_0_7; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_160 = 4'h8 == index ? _ram_0_T : ram_0_8; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_161 = 4'h9 == index ? _ram_0_T : ram_0_9; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_162 = 4'ha == index ? _ram_0_T : ram_0_10; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_163 = 4'hb == index ? _ram_0_T : ram_0_11; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_164 = 4'hc == index ? _ram_0_T : ram_0_12; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_165 = 4'hd == index ? _ram_0_T : ram_0_13; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_166 = 4'he == index ? _ram_0_T : ram_0_14; // @[i_cache.scala 19:24 86:{30,30}]
  wire [511:0] _GEN_167 = 4'hf == index ? _ram_0_T : ram_0_15; // @[i_cache.scala 19:24 86:{30,30}]
  wire [31:0] _GEN_168 = 4'h0 == index ? _GEN_2956 : tag_0_0; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_169 = 4'h1 == index ? _GEN_2956 : tag_0_1; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_170 = 4'h2 == index ? _GEN_2956 : tag_0_2; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_171 = 4'h3 == index ? _GEN_2956 : tag_0_3; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_172 = 4'h4 == index ? _GEN_2956 : tag_0_4; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_173 = 4'h5 == index ? _GEN_2956 : tag_0_5; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_174 = 4'h6 == index ? _GEN_2956 : tag_0_6; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_175 = 4'h7 == index ? _GEN_2956 : tag_0_7; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_176 = 4'h8 == index ? _GEN_2956 : tag_0_8; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_177 = 4'h9 == index ? _GEN_2956 : tag_0_9; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_178 = 4'ha == index ? _GEN_2956 : tag_0_10; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_179 = 4'hb == index ? _GEN_2956 : tag_0_11; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_180 = 4'hc == index ? _GEN_2956 : tag_0_12; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_181 = 4'hd == index ? _GEN_2956 : tag_0_13; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_182 = 4'he == index ? _GEN_2956 : tag_0_14; // @[i_cache.scala 23:24 87:{30,30}]
  wire [31:0] _GEN_183 = 4'hf == index ? _GEN_2956 : tag_0_15; // @[i_cache.scala 23:24 87:{30,30}]
  wire  _GEN_2969 = 4'h0 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_184 = 4'h0 == index | valid_0_0; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2970 = 4'h1 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_185 = 4'h1 == index | valid_0_1; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2971 = 4'h2 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_186 = 4'h2 == index | valid_0_2; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2972 = 4'h3 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_187 = 4'h3 == index | valid_0_3; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2973 = 4'h4 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_188 = 4'h4 == index | valid_0_4; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2974 = 4'h5 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_189 = 4'h5 == index | valid_0_5; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2975 = 4'h6 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_190 = 4'h6 == index | valid_0_6; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2976 = 4'h7 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_191 = 4'h7 == index | valid_0_7; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2977 = 4'h8 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_192 = 4'h8 == index | valid_0_8; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2978 = 4'h9 == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_193 = 4'h9 == index | valid_0_9; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2979 = 4'ha == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_194 = 4'ha == index | valid_0_10; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2980 = 4'hb == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_195 = 4'hb == index | valid_0_11; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2981 = 4'hc == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_196 = 4'hc == index | valid_0_12; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2982 = 4'hd == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_197 = 4'hd == index | valid_0_13; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2983 = 4'he == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_198 = 4'he == index | valid_0_14; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_2984 = 4'hf == index; // @[i_cache.scala 27:26 88:{32,32}]
  wire  _GEN_199 = 4'hf == index | valid_0_15; // @[i_cache.scala 27:26 88:{32,32}]
  wire [7:0] _GEN_201 = 4'h1 == index ? quene_1 : quene_0; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_202 = 4'h2 == index ? quene_2 : _GEN_201; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_203 = 4'h3 == index ? quene_3 : _GEN_202; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_204 = 4'h4 == index ? quene_4 : _GEN_203; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_205 = 4'h5 == index ? quene_5 : _GEN_204; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_206 = 4'h6 == index ? quene_6 : _GEN_205; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_207 = 4'h7 == index ? quene_7 : _GEN_206; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_208 = 4'h8 == index ? quene_8 : _GEN_207; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_209 = 4'h9 == index ? quene_9 : _GEN_208; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_210 = 4'ha == index ? quene_10 : _GEN_209; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_211 = 4'hb == index ? quene_11 : _GEN_210; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_212 = 4'hc == index ? quene_12 : _GEN_211; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_213 = 4'hd == index ? quene_13 : _GEN_212; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_214 = 4'he == index ? quene_14 : _GEN_213; // @[i_cache.scala 89:{46,46}]
  wire [7:0] _GEN_215 = 4'hf == index ? quene_15 : _GEN_214; // @[i_cache.scala 89:{46,46}]
  wire [9:0] _GEN_2985 = {_GEN_215, 2'h0}; // @[i_cache.scala 89:46]
  wire [10:0] _quene_T = {{1'd0}, _GEN_2985}; // @[i_cache.scala 89:46]
  wire [7:0] _GEN_216 = 4'h0 == index ? _quene_T[7:0] : quene_0; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_217 = 4'h1 == index ? _quene_T[7:0] : quene_1; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_218 = 4'h2 == index ? _quene_T[7:0] : quene_2; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_219 = 4'h3 == index ? _quene_T[7:0] : quene_3; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_220 = 4'h4 == index ? _quene_T[7:0] : quene_4; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_221 = 4'h5 == index ? _quene_T[7:0] : quene_5; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_222 = 4'h6 == index ? _quene_T[7:0] : quene_6; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_223 = 4'h7 == index ? _quene_T[7:0] : quene_7; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_224 = 4'h8 == index ? _quene_T[7:0] : quene_8; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_225 = 4'h9 == index ? _quene_T[7:0] : quene_9; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_226 = 4'ha == index ? _quene_T[7:0] : quene_10; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_227 = 4'hb == index ? _quene_T[7:0] : quene_11; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_228 = 4'hc == index ? _quene_T[7:0] : quene_12; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_229 = 4'hd == index ? _quene_T[7:0] : quene_13; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_230 = 4'he == index ? _quene_T[7:0] : quene_14; // @[i_cache.scala 40:24 89:{30,30}]
  wire [7:0] _GEN_231 = 4'hf == index ? _quene_T[7:0] : quene_15; // @[i_cache.scala 40:24 89:{30,30}]
  wire [511:0] _GEN_232 = 4'h0 == index ? _ram_0_T : ram_1_0; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_233 = 4'h1 == index ? _ram_0_T : ram_1_1; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_234 = 4'h2 == index ? _ram_0_T : ram_1_2; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_235 = 4'h3 == index ? _ram_0_T : ram_1_3; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_236 = 4'h4 == index ? _ram_0_T : ram_1_4; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_237 = 4'h5 == index ? _ram_0_T : ram_1_5; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_238 = 4'h6 == index ? _ram_0_T : ram_1_6; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_239 = 4'h7 == index ? _ram_0_T : ram_1_7; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_240 = 4'h8 == index ? _ram_0_T : ram_1_8; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_241 = 4'h9 == index ? _ram_0_T : ram_1_9; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_242 = 4'ha == index ? _ram_0_T : ram_1_10; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_243 = 4'hb == index ? _ram_0_T : ram_1_11; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_244 = 4'hc == index ? _ram_0_T : ram_1_12; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_245 = 4'hd == index ? _ram_0_T : ram_1_13; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_246 = 4'he == index ? _ram_0_T : ram_1_14; // @[i_cache.scala 20:24 91:{30,30}]
  wire [511:0] _GEN_247 = 4'hf == index ? _ram_0_T : ram_1_15; // @[i_cache.scala 20:24 91:{30,30}]
  wire [31:0] _GEN_248 = 4'h0 == index ? _GEN_2956 : tag_1_0; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_249 = 4'h1 == index ? _GEN_2956 : tag_1_1; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_250 = 4'h2 == index ? _GEN_2956 : tag_1_2; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_251 = 4'h3 == index ? _GEN_2956 : tag_1_3; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_252 = 4'h4 == index ? _GEN_2956 : tag_1_4; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_253 = 4'h5 == index ? _GEN_2956 : tag_1_5; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_254 = 4'h6 == index ? _GEN_2956 : tag_1_6; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_255 = 4'h7 == index ? _GEN_2956 : tag_1_7; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_256 = 4'h8 == index ? _GEN_2956 : tag_1_8; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_257 = 4'h9 == index ? _GEN_2956 : tag_1_9; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_258 = 4'ha == index ? _GEN_2956 : tag_1_10; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_259 = 4'hb == index ? _GEN_2956 : tag_1_11; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_260 = 4'hc == index ? _GEN_2956 : tag_1_12; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_261 = 4'hd == index ? _GEN_2956 : tag_1_13; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_262 = 4'he == index ? _GEN_2956 : tag_1_14; // @[i_cache.scala 24:24 92:{30,30}]
  wire [31:0] _GEN_263 = 4'hf == index ? _GEN_2956 : tag_1_15; // @[i_cache.scala 24:24 92:{30,30}]
  wire  _GEN_264 = _GEN_2969 | valid_1_0; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_265 = _GEN_2970 | valid_1_1; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_266 = _GEN_2971 | valid_1_2; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_267 = _GEN_2972 | valid_1_3; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_268 = _GEN_2973 | valid_1_4; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_269 = _GEN_2974 | valid_1_5; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_270 = _GEN_2975 | valid_1_6; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_271 = _GEN_2976 | valid_1_7; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_272 = _GEN_2977 | valid_1_8; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_273 = _GEN_2978 | valid_1_9; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_274 = _GEN_2979 | valid_1_10; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_275 = _GEN_2980 | valid_1_11; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_276 = _GEN_2981 | valid_1_12; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_277 = _GEN_2982 | valid_1_13; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_278 = _GEN_2983 | valid_1_14; // @[i_cache.scala 28:26 93:{32,32}]
  wire  _GEN_279 = _GEN_2984 | valid_1_15; // @[i_cache.scala 28:26 93:{32,32}]
  wire [10:0] _quene_T_2 = _quene_T | 11'h1; // @[i_cache.scala 94:55]
  wire [7:0] _GEN_280 = 4'h0 == index ? _quene_T_2[7:0] : quene_0; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_281 = 4'h1 == index ? _quene_T_2[7:0] : quene_1; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_282 = 4'h2 == index ? _quene_T_2[7:0] : quene_2; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_283 = 4'h3 == index ? _quene_T_2[7:0] : quene_3; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_284 = 4'h4 == index ? _quene_T_2[7:0] : quene_4; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_285 = 4'h5 == index ? _quene_T_2[7:0] : quene_5; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_286 = 4'h6 == index ? _quene_T_2[7:0] : quene_6; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_287 = 4'h7 == index ? _quene_T_2[7:0] : quene_7; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_288 = 4'h8 == index ? _quene_T_2[7:0] : quene_8; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_289 = 4'h9 == index ? _quene_T_2[7:0] : quene_9; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_290 = 4'ha == index ? _quene_T_2[7:0] : quene_10; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_291 = 4'hb == index ? _quene_T_2[7:0] : quene_11; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_292 = 4'hc == index ? _quene_T_2[7:0] : quene_12; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_293 = 4'hd == index ? _quene_T_2[7:0] : quene_13; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_294 = 4'he == index ? _quene_T_2[7:0] : quene_14; // @[i_cache.scala 40:24 94:{30,30}]
  wire [7:0] _GEN_295 = 4'hf == index ? _quene_T_2[7:0] : quene_15; // @[i_cache.scala 40:24 94:{30,30}]
  wire [511:0] _GEN_296 = 4'h0 == index ? _ram_0_T : ram_2_0; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_297 = 4'h1 == index ? _ram_0_T : ram_2_1; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_298 = 4'h2 == index ? _ram_0_T : ram_2_2; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_299 = 4'h3 == index ? _ram_0_T : ram_2_3; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_300 = 4'h4 == index ? _ram_0_T : ram_2_4; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_301 = 4'h5 == index ? _ram_0_T : ram_2_5; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_302 = 4'h6 == index ? _ram_0_T : ram_2_6; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_303 = 4'h7 == index ? _ram_0_T : ram_2_7; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_304 = 4'h8 == index ? _ram_0_T : ram_2_8; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_305 = 4'h9 == index ? _ram_0_T : ram_2_9; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_306 = 4'ha == index ? _ram_0_T : ram_2_10; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_307 = 4'hb == index ? _ram_0_T : ram_2_11; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_308 = 4'hc == index ? _ram_0_T : ram_2_12; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_309 = 4'hd == index ? _ram_0_T : ram_2_13; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_310 = 4'he == index ? _ram_0_T : ram_2_14; // @[i_cache.scala 21:24 96:{30,30}]
  wire [511:0] _GEN_311 = 4'hf == index ? _ram_0_T : ram_2_15; // @[i_cache.scala 21:24 96:{30,30}]
  wire [31:0] _GEN_312 = 4'h0 == index ? _GEN_2956 : tag_2_0; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_313 = 4'h1 == index ? _GEN_2956 : tag_2_1; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_314 = 4'h2 == index ? _GEN_2956 : tag_2_2; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_315 = 4'h3 == index ? _GEN_2956 : tag_2_3; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_316 = 4'h4 == index ? _GEN_2956 : tag_2_4; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_317 = 4'h5 == index ? _GEN_2956 : tag_2_5; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_318 = 4'h6 == index ? _GEN_2956 : tag_2_6; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_319 = 4'h7 == index ? _GEN_2956 : tag_2_7; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_320 = 4'h8 == index ? _GEN_2956 : tag_2_8; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_321 = 4'h9 == index ? _GEN_2956 : tag_2_9; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_322 = 4'ha == index ? _GEN_2956 : tag_2_10; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_323 = 4'hb == index ? _GEN_2956 : tag_2_11; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_324 = 4'hc == index ? _GEN_2956 : tag_2_12; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_325 = 4'hd == index ? _GEN_2956 : tag_2_13; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_326 = 4'he == index ? _GEN_2956 : tag_2_14; // @[i_cache.scala 25:24 97:{30,30}]
  wire [31:0] _GEN_327 = 4'hf == index ? _GEN_2956 : tag_2_15; // @[i_cache.scala 25:24 97:{30,30}]
  wire  _GEN_328 = _GEN_2969 | valid_2_0; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_329 = _GEN_2970 | valid_2_1; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_330 = _GEN_2971 | valid_2_2; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_331 = _GEN_2972 | valid_2_3; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_332 = _GEN_2973 | valid_2_4; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_333 = _GEN_2974 | valid_2_5; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_334 = _GEN_2975 | valid_2_6; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_335 = _GEN_2976 | valid_2_7; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_336 = _GEN_2977 | valid_2_8; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_337 = _GEN_2978 | valid_2_9; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_338 = _GEN_2979 | valid_2_10; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_339 = _GEN_2980 | valid_2_11; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_340 = _GEN_2981 | valid_2_12; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_341 = _GEN_2982 | valid_2_13; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_342 = _GEN_2983 | valid_2_14; // @[i_cache.scala 29:26 98:{32,32}]
  wire  _GEN_343 = _GEN_2984 | valid_2_15; // @[i_cache.scala 29:26 98:{32,32}]
  wire [10:0] _quene_T_4 = _quene_T | 11'h2; // @[i_cache.scala 99:55]
  wire [7:0] _GEN_344 = 4'h0 == index ? _quene_T_4[7:0] : quene_0; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_345 = 4'h1 == index ? _quene_T_4[7:0] : quene_1; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_346 = 4'h2 == index ? _quene_T_4[7:0] : quene_2; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_347 = 4'h3 == index ? _quene_T_4[7:0] : quene_3; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_348 = 4'h4 == index ? _quene_T_4[7:0] : quene_4; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_349 = 4'h5 == index ? _quene_T_4[7:0] : quene_5; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_350 = 4'h6 == index ? _quene_T_4[7:0] : quene_6; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_351 = 4'h7 == index ? _quene_T_4[7:0] : quene_7; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_352 = 4'h8 == index ? _quene_T_4[7:0] : quene_8; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_353 = 4'h9 == index ? _quene_T_4[7:0] : quene_9; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_354 = 4'ha == index ? _quene_T_4[7:0] : quene_10; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_355 = 4'hb == index ? _quene_T_4[7:0] : quene_11; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_356 = 4'hc == index ? _quene_T_4[7:0] : quene_12; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_357 = 4'hd == index ? _quene_T_4[7:0] : quene_13; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_358 = 4'he == index ? _quene_T_4[7:0] : quene_14; // @[i_cache.scala 40:24 99:{30,30}]
  wire [7:0] _GEN_359 = 4'hf == index ? _quene_T_4[7:0] : quene_15; // @[i_cache.scala 40:24 99:{30,30}]
  wire [511:0] _GEN_360 = 4'h0 == index ? _ram_0_T : ram_3_0; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_361 = 4'h1 == index ? _ram_0_T : ram_3_1; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_362 = 4'h2 == index ? _ram_0_T : ram_3_2; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_363 = 4'h3 == index ? _ram_0_T : ram_3_3; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_364 = 4'h4 == index ? _ram_0_T : ram_3_4; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_365 = 4'h5 == index ? _ram_0_T : ram_3_5; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_366 = 4'h6 == index ? _ram_0_T : ram_3_6; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_367 = 4'h7 == index ? _ram_0_T : ram_3_7; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_368 = 4'h8 == index ? _ram_0_T : ram_3_8; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_369 = 4'h9 == index ? _ram_0_T : ram_3_9; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_370 = 4'ha == index ? _ram_0_T : ram_3_10; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_371 = 4'hb == index ? _ram_0_T : ram_3_11; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_372 = 4'hc == index ? _ram_0_T : ram_3_12; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_373 = 4'hd == index ? _ram_0_T : ram_3_13; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_374 = 4'he == index ? _ram_0_T : ram_3_14; // @[i_cache.scala 101:{30,30} 22:24]
  wire [511:0] _GEN_375 = 4'hf == index ? _ram_0_T : ram_3_15; // @[i_cache.scala 101:{30,30} 22:24]
  wire [31:0] _GEN_376 = 4'h0 == index ? _GEN_2956 : tag_3_0; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_377 = 4'h1 == index ? _GEN_2956 : tag_3_1; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_378 = 4'h2 == index ? _GEN_2956 : tag_3_2; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_379 = 4'h3 == index ? _GEN_2956 : tag_3_3; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_380 = 4'h4 == index ? _GEN_2956 : tag_3_4; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_381 = 4'h5 == index ? _GEN_2956 : tag_3_5; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_382 = 4'h6 == index ? _GEN_2956 : tag_3_6; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_383 = 4'h7 == index ? _GEN_2956 : tag_3_7; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_384 = 4'h8 == index ? _GEN_2956 : tag_3_8; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_385 = 4'h9 == index ? _GEN_2956 : tag_3_9; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_386 = 4'ha == index ? _GEN_2956 : tag_3_10; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_387 = 4'hb == index ? _GEN_2956 : tag_3_11; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_388 = 4'hc == index ? _GEN_2956 : tag_3_12; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_389 = 4'hd == index ? _GEN_2956 : tag_3_13; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_390 = 4'he == index ? _GEN_2956 : tag_3_14; // @[i_cache.scala 102:{30,30} 26:24]
  wire [31:0] _GEN_391 = 4'hf == index ? _GEN_2956 : tag_3_15; // @[i_cache.scala 102:{30,30} 26:24]
  wire  _GEN_392 = _GEN_2969 | valid_3_0; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_393 = _GEN_2970 | valid_3_1; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_394 = _GEN_2971 | valid_3_2; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_395 = _GEN_2972 | valid_3_3; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_396 = _GEN_2973 | valid_3_4; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_397 = _GEN_2974 | valid_3_5; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_398 = _GEN_2975 | valid_3_6; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_399 = _GEN_2976 | valid_3_7; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_400 = _GEN_2977 | valid_3_8; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_401 = _GEN_2978 | valid_3_9; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_402 = _GEN_2979 | valid_3_10; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_403 = _GEN_2980 | valid_3_11; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_404 = _GEN_2981 | valid_3_12; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_405 = _GEN_2982 | valid_3_13; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_406 = _GEN_2983 | valid_3_14; // @[i_cache.scala 103:{32,32} 30:26]
  wire  _GEN_407 = _GEN_2984 | valid_3_15; // @[i_cache.scala 103:{32,32} 30:26]
  wire [10:0] _quene_T_6 = _quene_T | 11'h3; // @[i_cache.scala 104:55]
  wire [7:0] _GEN_408 = 4'h0 == index ? _quene_T_6[7:0] : quene_0; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_409 = 4'h1 == index ? _quene_T_6[7:0] : quene_1; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_410 = 4'h2 == index ? _quene_T_6[7:0] : quene_2; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_411 = 4'h3 == index ? _quene_T_6[7:0] : quene_3; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_412 = 4'h4 == index ? _quene_T_6[7:0] : quene_4; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_413 = 4'h5 == index ? _quene_T_6[7:0] : quene_5; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_414 = 4'h6 == index ? _quene_T_6[7:0] : quene_6; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_415 = 4'h7 == index ? _quene_T_6[7:0] : quene_7; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_416 = 4'h8 == index ? _quene_T_6[7:0] : quene_8; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_417 = 4'h9 == index ? _quene_T_6[7:0] : quene_9; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_418 = 4'ha == index ? _quene_T_6[7:0] : quene_10; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_419 = 4'hb == index ? _quene_T_6[7:0] : quene_11; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_420 = 4'hc == index ? _quene_T_6[7:0] : quene_12; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_421 = 4'hd == index ? _quene_T_6[7:0] : quene_13; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_422 = 4'he == index ? _quene_T_6[7:0] : quene_14; // @[i_cache.scala 104:{30,30} 40:24]
  wire [7:0] _GEN_423 = 4'hf == index ? _quene_T_6[7:0] : quene_15; // @[i_cache.scala 104:{30,30} 40:24]
  wire [511:0] _GEN_680 = _GEN_215[7:6] == 2'h2 ? _GEN_296 : ram_2_0; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_681 = _GEN_215[7:6] == 2'h2 ? _GEN_297 : ram_2_1; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_682 = _GEN_215[7:6] == 2'h2 ? _GEN_298 : ram_2_2; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_683 = _GEN_215[7:6] == 2'h2 ? _GEN_299 : ram_2_3; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_684 = _GEN_215[7:6] == 2'h2 ? _GEN_300 : ram_2_4; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_685 = _GEN_215[7:6] == 2'h2 ? _GEN_301 : ram_2_5; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_686 = _GEN_215[7:6] == 2'h2 ? _GEN_302 : ram_2_6; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_687 = _GEN_215[7:6] == 2'h2 ? _GEN_303 : ram_2_7; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_688 = _GEN_215[7:6] == 2'h2 ? _GEN_304 : ram_2_8; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_689 = _GEN_215[7:6] == 2'h2 ? _GEN_305 : ram_2_9; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_690 = _GEN_215[7:6] == 2'h2 ? _GEN_306 : ram_2_10; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_691 = _GEN_215[7:6] == 2'h2 ? _GEN_307 : ram_2_11; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_692 = _GEN_215[7:6] == 2'h2 ? _GEN_308 : ram_2_12; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_693 = _GEN_215[7:6] == 2'h2 ? _GEN_309 : ram_2_13; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_694 = _GEN_215[7:6] == 2'h2 ? _GEN_310 : ram_2_14; // @[i_cache.scala 116:52 21:24]
  wire [511:0] _GEN_695 = _GEN_215[7:6] == 2'h2 ? _GEN_311 : ram_2_15; // @[i_cache.scala 116:52 21:24]
  wire [31:0] _GEN_696 = _GEN_215[7:6] == 2'h2 ? _GEN_312 : tag_2_0; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_697 = _GEN_215[7:6] == 2'h2 ? _GEN_313 : tag_2_1; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_698 = _GEN_215[7:6] == 2'h2 ? _GEN_314 : tag_2_2; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_699 = _GEN_215[7:6] == 2'h2 ? _GEN_315 : tag_2_3; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_700 = _GEN_215[7:6] == 2'h2 ? _GEN_316 : tag_2_4; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_701 = _GEN_215[7:6] == 2'h2 ? _GEN_317 : tag_2_5; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_702 = _GEN_215[7:6] == 2'h2 ? _GEN_318 : tag_2_6; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_703 = _GEN_215[7:6] == 2'h2 ? _GEN_319 : tag_2_7; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_704 = _GEN_215[7:6] == 2'h2 ? _GEN_320 : tag_2_8; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_705 = _GEN_215[7:6] == 2'h2 ? _GEN_321 : tag_2_9; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_706 = _GEN_215[7:6] == 2'h2 ? _GEN_322 : tag_2_10; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_707 = _GEN_215[7:6] == 2'h2 ? _GEN_323 : tag_2_11; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_708 = _GEN_215[7:6] == 2'h2 ? _GEN_324 : tag_2_12; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_709 = _GEN_215[7:6] == 2'h2 ? _GEN_325 : tag_2_13; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_710 = _GEN_215[7:6] == 2'h2 ? _GEN_326 : tag_2_14; // @[i_cache.scala 116:52 25:24]
  wire [31:0] _GEN_711 = _GEN_215[7:6] == 2'h2 ? _GEN_327 : tag_2_15; // @[i_cache.scala 116:52 25:24]
  wire  _GEN_712 = _GEN_215[7:6] == 2'h2 ? _GEN_328 : valid_2_0; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_713 = _GEN_215[7:6] == 2'h2 ? _GEN_329 : valid_2_1; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_714 = _GEN_215[7:6] == 2'h2 ? _GEN_330 : valid_2_2; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_715 = _GEN_215[7:6] == 2'h2 ? _GEN_331 : valid_2_3; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_716 = _GEN_215[7:6] == 2'h2 ? _GEN_332 : valid_2_4; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_717 = _GEN_215[7:6] == 2'h2 ? _GEN_333 : valid_2_5; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_718 = _GEN_215[7:6] == 2'h2 ? _GEN_334 : valid_2_6; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_719 = _GEN_215[7:6] == 2'h2 ? _GEN_335 : valid_2_7; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_720 = _GEN_215[7:6] == 2'h2 ? _GEN_336 : valid_2_8; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_721 = _GEN_215[7:6] == 2'h2 ? _GEN_337 : valid_2_9; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_722 = _GEN_215[7:6] == 2'h2 ? _GEN_338 : valid_2_10; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_723 = _GEN_215[7:6] == 2'h2 ? _GEN_339 : valid_2_11; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_724 = _GEN_215[7:6] == 2'h2 ? _GEN_340 : valid_2_12; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_725 = _GEN_215[7:6] == 2'h2 ? _GEN_341 : valid_2_13; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_726 = _GEN_215[7:6] == 2'h2 ? _GEN_342 : valid_2_14; // @[i_cache.scala 116:52 29:26]
  wire  _GEN_727 = _GEN_215[7:6] == 2'h2 ? _GEN_343 : valid_2_15; // @[i_cache.scala 116:52 29:26]
  wire [7:0] _GEN_728 = _GEN_215[7:6] == 2'h2 ? _GEN_344 : _GEN_408; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_729 = _GEN_215[7:6] == 2'h2 ? _GEN_345 : _GEN_409; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_730 = _GEN_215[7:6] == 2'h2 ? _GEN_346 : _GEN_410; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_731 = _GEN_215[7:6] == 2'h2 ? _GEN_347 : _GEN_411; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_732 = _GEN_215[7:6] == 2'h2 ? _GEN_348 : _GEN_412; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_733 = _GEN_215[7:6] == 2'h2 ? _GEN_349 : _GEN_413; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_734 = _GEN_215[7:6] == 2'h2 ? _GEN_350 : _GEN_414; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_735 = _GEN_215[7:6] == 2'h2 ? _GEN_351 : _GEN_415; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_736 = _GEN_215[7:6] == 2'h2 ? _GEN_352 : _GEN_416; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_737 = _GEN_215[7:6] == 2'h2 ? _GEN_353 : _GEN_417; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_738 = _GEN_215[7:6] == 2'h2 ? _GEN_354 : _GEN_418; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_739 = _GEN_215[7:6] == 2'h2 ? _GEN_355 : _GEN_419; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_740 = _GEN_215[7:6] == 2'h2 ? _GEN_356 : _GEN_420; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_741 = _GEN_215[7:6] == 2'h2 ? _GEN_357 : _GEN_421; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_742 = _GEN_215[7:6] == 2'h2 ? _GEN_358 : _GEN_422; // @[i_cache.scala 116:52]
  wire [7:0] _GEN_743 = _GEN_215[7:6] == 2'h2 ? _GEN_359 : _GEN_423; // @[i_cache.scala 116:52]
  wire [511:0] _GEN_744 = _GEN_215[7:6] == 2'h2 ? ram_3_0 : _GEN_360; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_745 = _GEN_215[7:6] == 2'h2 ? ram_3_1 : _GEN_361; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_746 = _GEN_215[7:6] == 2'h2 ? ram_3_2 : _GEN_362; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_747 = _GEN_215[7:6] == 2'h2 ? ram_3_3 : _GEN_363; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_748 = _GEN_215[7:6] == 2'h2 ? ram_3_4 : _GEN_364; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_749 = _GEN_215[7:6] == 2'h2 ? ram_3_5 : _GEN_365; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_750 = _GEN_215[7:6] == 2'h2 ? ram_3_6 : _GEN_366; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_751 = _GEN_215[7:6] == 2'h2 ? ram_3_7 : _GEN_367; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_752 = _GEN_215[7:6] == 2'h2 ? ram_3_8 : _GEN_368; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_753 = _GEN_215[7:6] == 2'h2 ? ram_3_9 : _GEN_369; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_754 = _GEN_215[7:6] == 2'h2 ? ram_3_10 : _GEN_370; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_755 = _GEN_215[7:6] == 2'h2 ? ram_3_11 : _GEN_371; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_756 = _GEN_215[7:6] == 2'h2 ? ram_3_12 : _GEN_372; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_757 = _GEN_215[7:6] == 2'h2 ? ram_3_13 : _GEN_373; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_758 = _GEN_215[7:6] == 2'h2 ? ram_3_14 : _GEN_374; // @[i_cache.scala 116:52 22:24]
  wire [511:0] _GEN_759 = _GEN_215[7:6] == 2'h2 ? ram_3_15 : _GEN_375; // @[i_cache.scala 116:52 22:24]
  wire [31:0] _GEN_760 = _GEN_215[7:6] == 2'h2 ? tag_3_0 : _GEN_376; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_761 = _GEN_215[7:6] == 2'h2 ? tag_3_1 : _GEN_377; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_762 = _GEN_215[7:6] == 2'h2 ? tag_3_2 : _GEN_378; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_763 = _GEN_215[7:6] == 2'h2 ? tag_3_3 : _GEN_379; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_764 = _GEN_215[7:6] == 2'h2 ? tag_3_4 : _GEN_380; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_765 = _GEN_215[7:6] == 2'h2 ? tag_3_5 : _GEN_381; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_766 = _GEN_215[7:6] == 2'h2 ? tag_3_6 : _GEN_382; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_767 = _GEN_215[7:6] == 2'h2 ? tag_3_7 : _GEN_383; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_768 = _GEN_215[7:6] == 2'h2 ? tag_3_8 : _GEN_384; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_769 = _GEN_215[7:6] == 2'h2 ? tag_3_9 : _GEN_385; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_770 = _GEN_215[7:6] == 2'h2 ? tag_3_10 : _GEN_386; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_771 = _GEN_215[7:6] == 2'h2 ? tag_3_11 : _GEN_387; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_772 = _GEN_215[7:6] == 2'h2 ? tag_3_12 : _GEN_388; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_773 = _GEN_215[7:6] == 2'h2 ? tag_3_13 : _GEN_389; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_774 = _GEN_215[7:6] == 2'h2 ? tag_3_14 : _GEN_390; // @[i_cache.scala 116:52 26:24]
  wire [31:0] _GEN_775 = _GEN_215[7:6] == 2'h2 ? tag_3_15 : _GEN_391; // @[i_cache.scala 116:52 26:24]
  wire  _GEN_776 = _GEN_215[7:6] == 2'h2 ? valid_3_0 : _GEN_392; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_777 = _GEN_215[7:6] == 2'h2 ? valid_3_1 : _GEN_393; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_778 = _GEN_215[7:6] == 2'h2 ? valid_3_2 : _GEN_394; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_779 = _GEN_215[7:6] == 2'h2 ? valid_3_3 : _GEN_395; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_780 = _GEN_215[7:6] == 2'h2 ? valid_3_4 : _GEN_396; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_781 = _GEN_215[7:6] == 2'h2 ? valid_3_5 : _GEN_397; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_782 = _GEN_215[7:6] == 2'h2 ? valid_3_6 : _GEN_398; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_783 = _GEN_215[7:6] == 2'h2 ? valid_3_7 : _GEN_399; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_784 = _GEN_215[7:6] == 2'h2 ? valid_3_8 : _GEN_400; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_785 = _GEN_215[7:6] == 2'h2 ? valid_3_9 : _GEN_401; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_786 = _GEN_215[7:6] == 2'h2 ? valid_3_10 : _GEN_402; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_787 = _GEN_215[7:6] == 2'h2 ? valid_3_11 : _GEN_403; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_788 = _GEN_215[7:6] == 2'h2 ? valid_3_12 : _GEN_404; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_789 = _GEN_215[7:6] == 2'h2 ? valid_3_13 : _GEN_405; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_790 = _GEN_215[7:6] == 2'h2 ? valid_3_14 : _GEN_406; // @[i_cache.scala 116:52 30:26]
  wire  _GEN_791 = _GEN_215[7:6] == 2'h2 ? valid_3_15 : _GEN_407; // @[i_cache.scala 116:52 30:26]
  wire [511:0] _GEN_792 = _GEN_215[7:6] == 2'h1 ? _GEN_232 : ram_1_0; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_793 = _GEN_215[7:6] == 2'h1 ? _GEN_233 : ram_1_1; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_794 = _GEN_215[7:6] == 2'h1 ? _GEN_234 : ram_1_2; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_795 = _GEN_215[7:6] == 2'h1 ? _GEN_235 : ram_1_3; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_796 = _GEN_215[7:6] == 2'h1 ? _GEN_236 : ram_1_4; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_797 = _GEN_215[7:6] == 2'h1 ? _GEN_237 : ram_1_5; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_798 = _GEN_215[7:6] == 2'h1 ? _GEN_238 : ram_1_6; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_799 = _GEN_215[7:6] == 2'h1 ? _GEN_239 : ram_1_7; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_800 = _GEN_215[7:6] == 2'h1 ? _GEN_240 : ram_1_8; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_801 = _GEN_215[7:6] == 2'h1 ? _GEN_241 : ram_1_9; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_802 = _GEN_215[7:6] == 2'h1 ? _GEN_242 : ram_1_10; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_803 = _GEN_215[7:6] == 2'h1 ? _GEN_243 : ram_1_11; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_804 = _GEN_215[7:6] == 2'h1 ? _GEN_244 : ram_1_12; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_805 = _GEN_215[7:6] == 2'h1 ? _GEN_245 : ram_1_13; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_806 = _GEN_215[7:6] == 2'h1 ? _GEN_246 : ram_1_14; // @[i_cache.scala 111:52 20:24]
  wire [511:0] _GEN_807 = _GEN_215[7:6] == 2'h1 ? _GEN_247 : ram_1_15; // @[i_cache.scala 111:52 20:24]
  wire [31:0] _GEN_808 = _GEN_215[7:6] == 2'h1 ? _GEN_248 : tag_1_0; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_809 = _GEN_215[7:6] == 2'h1 ? _GEN_249 : tag_1_1; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_810 = _GEN_215[7:6] == 2'h1 ? _GEN_250 : tag_1_2; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_811 = _GEN_215[7:6] == 2'h1 ? _GEN_251 : tag_1_3; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_812 = _GEN_215[7:6] == 2'h1 ? _GEN_252 : tag_1_4; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_813 = _GEN_215[7:6] == 2'h1 ? _GEN_253 : tag_1_5; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_814 = _GEN_215[7:6] == 2'h1 ? _GEN_254 : tag_1_6; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_815 = _GEN_215[7:6] == 2'h1 ? _GEN_255 : tag_1_7; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_816 = _GEN_215[7:6] == 2'h1 ? _GEN_256 : tag_1_8; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_817 = _GEN_215[7:6] == 2'h1 ? _GEN_257 : tag_1_9; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_818 = _GEN_215[7:6] == 2'h1 ? _GEN_258 : tag_1_10; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_819 = _GEN_215[7:6] == 2'h1 ? _GEN_259 : tag_1_11; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_820 = _GEN_215[7:6] == 2'h1 ? _GEN_260 : tag_1_12; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_821 = _GEN_215[7:6] == 2'h1 ? _GEN_261 : tag_1_13; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_822 = _GEN_215[7:6] == 2'h1 ? _GEN_262 : tag_1_14; // @[i_cache.scala 111:52 24:24]
  wire [31:0] _GEN_823 = _GEN_215[7:6] == 2'h1 ? _GEN_263 : tag_1_15; // @[i_cache.scala 111:52 24:24]
  wire  _GEN_824 = _GEN_215[7:6] == 2'h1 ? _GEN_264 : valid_1_0; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_825 = _GEN_215[7:6] == 2'h1 ? _GEN_265 : valid_1_1; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_826 = _GEN_215[7:6] == 2'h1 ? _GEN_266 : valid_1_2; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_827 = _GEN_215[7:6] == 2'h1 ? _GEN_267 : valid_1_3; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_828 = _GEN_215[7:6] == 2'h1 ? _GEN_268 : valid_1_4; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_829 = _GEN_215[7:6] == 2'h1 ? _GEN_269 : valid_1_5; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_830 = _GEN_215[7:6] == 2'h1 ? _GEN_270 : valid_1_6; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_831 = _GEN_215[7:6] == 2'h1 ? _GEN_271 : valid_1_7; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_832 = _GEN_215[7:6] == 2'h1 ? _GEN_272 : valid_1_8; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_833 = _GEN_215[7:6] == 2'h1 ? _GEN_273 : valid_1_9; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_834 = _GEN_215[7:6] == 2'h1 ? _GEN_274 : valid_1_10; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_835 = _GEN_215[7:6] == 2'h1 ? _GEN_275 : valid_1_11; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_836 = _GEN_215[7:6] == 2'h1 ? _GEN_276 : valid_1_12; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_837 = _GEN_215[7:6] == 2'h1 ? _GEN_277 : valid_1_13; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_838 = _GEN_215[7:6] == 2'h1 ? _GEN_278 : valid_1_14; // @[i_cache.scala 111:52 28:26]
  wire  _GEN_839 = _GEN_215[7:6] == 2'h1 ? _GEN_279 : valid_1_15; // @[i_cache.scala 111:52 28:26]
  wire [7:0] _GEN_840 = _GEN_215[7:6] == 2'h1 ? _GEN_280 : _GEN_728; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_841 = _GEN_215[7:6] == 2'h1 ? _GEN_281 : _GEN_729; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_842 = _GEN_215[7:6] == 2'h1 ? _GEN_282 : _GEN_730; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_843 = _GEN_215[7:6] == 2'h1 ? _GEN_283 : _GEN_731; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_844 = _GEN_215[7:6] == 2'h1 ? _GEN_284 : _GEN_732; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_845 = _GEN_215[7:6] == 2'h1 ? _GEN_285 : _GEN_733; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_846 = _GEN_215[7:6] == 2'h1 ? _GEN_286 : _GEN_734; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_847 = _GEN_215[7:6] == 2'h1 ? _GEN_287 : _GEN_735; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_848 = _GEN_215[7:6] == 2'h1 ? _GEN_288 : _GEN_736; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_849 = _GEN_215[7:6] == 2'h1 ? _GEN_289 : _GEN_737; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_850 = _GEN_215[7:6] == 2'h1 ? _GEN_290 : _GEN_738; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_851 = _GEN_215[7:6] == 2'h1 ? _GEN_291 : _GEN_739; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_852 = _GEN_215[7:6] == 2'h1 ? _GEN_292 : _GEN_740; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_853 = _GEN_215[7:6] == 2'h1 ? _GEN_293 : _GEN_741; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_854 = _GEN_215[7:6] == 2'h1 ? _GEN_294 : _GEN_742; // @[i_cache.scala 111:52]
  wire [7:0] _GEN_855 = _GEN_215[7:6] == 2'h1 ? _GEN_295 : _GEN_743; // @[i_cache.scala 111:52]
  wire [511:0] _GEN_856 = _GEN_215[7:6] == 2'h1 ? ram_2_0 : _GEN_680; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_857 = _GEN_215[7:6] == 2'h1 ? ram_2_1 : _GEN_681; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_858 = _GEN_215[7:6] == 2'h1 ? ram_2_2 : _GEN_682; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_859 = _GEN_215[7:6] == 2'h1 ? ram_2_3 : _GEN_683; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_860 = _GEN_215[7:6] == 2'h1 ? ram_2_4 : _GEN_684; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_861 = _GEN_215[7:6] == 2'h1 ? ram_2_5 : _GEN_685; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_862 = _GEN_215[7:6] == 2'h1 ? ram_2_6 : _GEN_686; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_863 = _GEN_215[7:6] == 2'h1 ? ram_2_7 : _GEN_687; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_864 = _GEN_215[7:6] == 2'h1 ? ram_2_8 : _GEN_688; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_865 = _GEN_215[7:6] == 2'h1 ? ram_2_9 : _GEN_689; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_866 = _GEN_215[7:6] == 2'h1 ? ram_2_10 : _GEN_690; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_867 = _GEN_215[7:6] == 2'h1 ? ram_2_11 : _GEN_691; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_868 = _GEN_215[7:6] == 2'h1 ? ram_2_12 : _GEN_692; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_869 = _GEN_215[7:6] == 2'h1 ? ram_2_13 : _GEN_693; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_870 = _GEN_215[7:6] == 2'h1 ? ram_2_14 : _GEN_694; // @[i_cache.scala 111:52 21:24]
  wire [511:0] _GEN_871 = _GEN_215[7:6] == 2'h1 ? ram_2_15 : _GEN_695; // @[i_cache.scala 111:52 21:24]
  wire [31:0] _GEN_872 = _GEN_215[7:6] == 2'h1 ? tag_2_0 : _GEN_696; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_873 = _GEN_215[7:6] == 2'h1 ? tag_2_1 : _GEN_697; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_874 = _GEN_215[7:6] == 2'h1 ? tag_2_2 : _GEN_698; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_875 = _GEN_215[7:6] == 2'h1 ? tag_2_3 : _GEN_699; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_876 = _GEN_215[7:6] == 2'h1 ? tag_2_4 : _GEN_700; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_877 = _GEN_215[7:6] == 2'h1 ? tag_2_5 : _GEN_701; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_878 = _GEN_215[7:6] == 2'h1 ? tag_2_6 : _GEN_702; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_879 = _GEN_215[7:6] == 2'h1 ? tag_2_7 : _GEN_703; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_880 = _GEN_215[7:6] == 2'h1 ? tag_2_8 : _GEN_704; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_881 = _GEN_215[7:6] == 2'h1 ? tag_2_9 : _GEN_705; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_882 = _GEN_215[7:6] == 2'h1 ? tag_2_10 : _GEN_706; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_883 = _GEN_215[7:6] == 2'h1 ? tag_2_11 : _GEN_707; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_884 = _GEN_215[7:6] == 2'h1 ? tag_2_12 : _GEN_708; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_885 = _GEN_215[7:6] == 2'h1 ? tag_2_13 : _GEN_709; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_886 = _GEN_215[7:6] == 2'h1 ? tag_2_14 : _GEN_710; // @[i_cache.scala 111:52 25:24]
  wire [31:0] _GEN_887 = _GEN_215[7:6] == 2'h1 ? tag_2_15 : _GEN_711; // @[i_cache.scala 111:52 25:24]
  wire  _GEN_888 = _GEN_215[7:6] == 2'h1 ? valid_2_0 : _GEN_712; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_889 = _GEN_215[7:6] == 2'h1 ? valid_2_1 : _GEN_713; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_890 = _GEN_215[7:6] == 2'h1 ? valid_2_2 : _GEN_714; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_891 = _GEN_215[7:6] == 2'h1 ? valid_2_3 : _GEN_715; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_892 = _GEN_215[7:6] == 2'h1 ? valid_2_4 : _GEN_716; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_893 = _GEN_215[7:6] == 2'h1 ? valid_2_5 : _GEN_717; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_894 = _GEN_215[7:6] == 2'h1 ? valid_2_6 : _GEN_718; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_895 = _GEN_215[7:6] == 2'h1 ? valid_2_7 : _GEN_719; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_896 = _GEN_215[7:6] == 2'h1 ? valid_2_8 : _GEN_720; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_897 = _GEN_215[7:6] == 2'h1 ? valid_2_9 : _GEN_721; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_898 = _GEN_215[7:6] == 2'h1 ? valid_2_10 : _GEN_722; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_899 = _GEN_215[7:6] == 2'h1 ? valid_2_11 : _GEN_723; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_900 = _GEN_215[7:6] == 2'h1 ? valid_2_12 : _GEN_724; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_901 = _GEN_215[7:6] == 2'h1 ? valid_2_13 : _GEN_725; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_902 = _GEN_215[7:6] == 2'h1 ? valid_2_14 : _GEN_726; // @[i_cache.scala 111:52 29:26]
  wire  _GEN_903 = _GEN_215[7:6] == 2'h1 ? valid_2_15 : _GEN_727; // @[i_cache.scala 111:52 29:26]
  wire [511:0] _GEN_904 = _GEN_215[7:6] == 2'h1 ? ram_3_0 : _GEN_744; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_905 = _GEN_215[7:6] == 2'h1 ? ram_3_1 : _GEN_745; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_906 = _GEN_215[7:6] == 2'h1 ? ram_3_2 : _GEN_746; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_907 = _GEN_215[7:6] == 2'h1 ? ram_3_3 : _GEN_747; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_908 = _GEN_215[7:6] == 2'h1 ? ram_3_4 : _GEN_748; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_909 = _GEN_215[7:6] == 2'h1 ? ram_3_5 : _GEN_749; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_910 = _GEN_215[7:6] == 2'h1 ? ram_3_6 : _GEN_750; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_911 = _GEN_215[7:6] == 2'h1 ? ram_3_7 : _GEN_751; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_912 = _GEN_215[7:6] == 2'h1 ? ram_3_8 : _GEN_752; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_913 = _GEN_215[7:6] == 2'h1 ? ram_3_9 : _GEN_753; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_914 = _GEN_215[7:6] == 2'h1 ? ram_3_10 : _GEN_754; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_915 = _GEN_215[7:6] == 2'h1 ? ram_3_11 : _GEN_755; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_916 = _GEN_215[7:6] == 2'h1 ? ram_3_12 : _GEN_756; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_917 = _GEN_215[7:6] == 2'h1 ? ram_3_13 : _GEN_757; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_918 = _GEN_215[7:6] == 2'h1 ? ram_3_14 : _GEN_758; // @[i_cache.scala 111:52 22:24]
  wire [511:0] _GEN_919 = _GEN_215[7:6] == 2'h1 ? ram_3_15 : _GEN_759; // @[i_cache.scala 111:52 22:24]
  wire [31:0] _GEN_920 = _GEN_215[7:6] == 2'h1 ? tag_3_0 : _GEN_760; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_921 = _GEN_215[7:6] == 2'h1 ? tag_3_1 : _GEN_761; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_922 = _GEN_215[7:6] == 2'h1 ? tag_3_2 : _GEN_762; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_923 = _GEN_215[7:6] == 2'h1 ? tag_3_3 : _GEN_763; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_924 = _GEN_215[7:6] == 2'h1 ? tag_3_4 : _GEN_764; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_925 = _GEN_215[7:6] == 2'h1 ? tag_3_5 : _GEN_765; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_926 = _GEN_215[7:6] == 2'h1 ? tag_3_6 : _GEN_766; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_927 = _GEN_215[7:6] == 2'h1 ? tag_3_7 : _GEN_767; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_928 = _GEN_215[7:6] == 2'h1 ? tag_3_8 : _GEN_768; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_929 = _GEN_215[7:6] == 2'h1 ? tag_3_9 : _GEN_769; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_930 = _GEN_215[7:6] == 2'h1 ? tag_3_10 : _GEN_770; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_931 = _GEN_215[7:6] == 2'h1 ? tag_3_11 : _GEN_771; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_932 = _GEN_215[7:6] == 2'h1 ? tag_3_12 : _GEN_772; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_933 = _GEN_215[7:6] == 2'h1 ? tag_3_13 : _GEN_773; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_934 = _GEN_215[7:6] == 2'h1 ? tag_3_14 : _GEN_774; // @[i_cache.scala 111:52 26:24]
  wire [31:0] _GEN_935 = _GEN_215[7:6] == 2'h1 ? tag_3_15 : _GEN_775; // @[i_cache.scala 111:52 26:24]
  wire  _GEN_936 = _GEN_215[7:6] == 2'h1 ? valid_3_0 : _GEN_776; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_937 = _GEN_215[7:6] == 2'h1 ? valid_3_1 : _GEN_777; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_938 = _GEN_215[7:6] == 2'h1 ? valid_3_2 : _GEN_778; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_939 = _GEN_215[7:6] == 2'h1 ? valid_3_3 : _GEN_779; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_940 = _GEN_215[7:6] == 2'h1 ? valid_3_4 : _GEN_780; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_941 = _GEN_215[7:6] == 2'h1 ? valid_3_5 : _GEN_781; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_942 = _GEN_215[7:6] == 2'h1 ? valid_3_6 : _GEN_782; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_943 = _GEN_215[7:6] == 2'h1 ? valid_3_7 : _GEN_783; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_944 = _GEN_215[7:6] == 2'h1 ? valid_3_8 : _GEN_784; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_945 = _GEN_215[7:6] == 2'h1 ? valid_3_9 : _GEN_785; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_946 = _GEN_215[7:6] == 2'h1 ? valid_3_10 : _GEN_786; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_947 = _GEN_215[7:6] == 2'h1 ? valid_3_11 : _GEN_787; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_948 = _GEN_215[7:6] == 2'h1 ? valid_3_12 : _GEN_788; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_949 = _GEN_215[7:6] == 2'h1 ? valid_3_13 : _GEN_789; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_950 = _GEN_215[7:6] == 2'h1 ? valid_3_14 : _GEN_790; // @[i_cache.scala 111:52 30:26]
  wire  _GEN_951 = _GEN_215[7:6] == 2'h1 ? valid_3_15 : _GEN_791; // @[i_cache.scala 111:52 30:26]
  wire [511:0] _GEN_952 = _GEN_215[7:6] == 2'h0 ? _GEN_152 : ram_0_0; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_953 = _GEN_215[7:6] == 2'h0 ? _GEN_153 : ram_0_1; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_954 = _GEN_215[7:6] == 2'h0 ? _GEN_154 : ram_0_2; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_955 = _GEN_215[7:6] == 2'h0 ? _GEN_155 : ram_0_3; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_956 = _GEN_215[7:6] == 2'h0 ? _GEN_156 : ram_0_4; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_957 = _GEN_215[7:6] == 2'h0 ? _GEN_157 : ram_0_5; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_958 = _GEN_215[7:6] == 2'h0 ? _GEN_158 : ram_0_6; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_959 = _GEN_215[7:6] == 2'h0 ? _GEN_159 : ram_0_7; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_960 = _GEN_215[7:6] == 2'h0 ? _GEN_160 : ram_0_8; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_961 = _GEN_215[7:6] == 2'h0 ? _GEN_161 : ram_0_9; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_962 = _GEN_215[7:6] == 2'h0 ? _GEN_162 : ram_0_10; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_963 = _GEN_215[7:6] == 2'h0 ? _GEN_163 : ram_0_11; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_964 = _GEN_215[7:6] == 2'h0 ? _GEN_164 : ram_0_12; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_965 = _GEN_215[7:6] == 2'h0 ? _GEN_165 : ram_0_13; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_966 = _GEN_215[7:6] == 2'h0 ? _GEN_166 : ram_0_14; // @[i_cache.scala 106:46 19:24]
  wire [511:0] _GEN_967 = _GEN_215[7:6] == 2'h0 ? _GEN_167 : ram_0_15; // @[i_cache.scala 106:46 19:24]
  wire [31:0] _GEN_968 = _GEN_215[7:6] == 2'h0 ? _GEN_168 : tag_0_0; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_969 = _GEN_215[7:6] == 2'h0 ? _GEN_169 : tag_0_1; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_970 = _GEN_215[7:6] == 2'h0 ? _GEN_170 : tag_0_2; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_971 = _GEN_215[7:6] == 2'h0 ? _GEN_171 : tag_0_3; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_972 = _GEN_215[7:6] == 2'h0 ? _GEN_172 : tag_0_4; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_973 = _GEN_215[7:6] == 2'h0 ? _GEN_173 : tag_0_5; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_974 = _GEN_215[7:6] == 2'h0 ? _GEN_174 : tag_0_6; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_975 = _GEN_215[7:6] == 2'h0 ? _GEN_175 : tag_0_7; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_976 = _GEN_215[7:6] == 2'h0 ? _GEN_176 : tag_0_8; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_977 = _GEN_215[7:6] == 2'h0 ? _GEN_177 : tag_0_9; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_978 = _GEN_215[7:6] == 2'h0 ? _GEN_178 : tag_0_10; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_979 = _GEN_215[7:6] == 2'h0 ? _GEN_179 : tag_0_11; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_980 = _GEN_215[7:6] == 2'h0 ? _GEN_180 : tag_0_12; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_981 = _GEN_215[7:6] == 2'h0 ? _GEN_181 : tag_0_13; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_982 = _GEN_215[7:6] == 2'h0 ? _GEN_182 : tag_0_14; // @[i_cache.scala 106:46 23:24]
  wire [31:0] _GEN_983 = _GEN_215[7:6] == 2'h0 ? _GEN_183 : tag_0_15; // @[i_cache.scala 106:46 23:24]
  wire  _GEN_984 = _GEN_215[7:6] == 2'h0 ? _GEN_184 : valid_0_0; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_985 = _GEN_215[7:6] == 2'h0 ? _GEN_185 : valid_0_1; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_986 = _GEN_215[7:6] == 2'h0 ? _GEN_186 : valid_0_2; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_987 = _GEN_215[7:6] == 2'h0 ? _GEN_187 : valid_0_3; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_988 = _GEN_215[7:6] == 2'h0 ? _GEN_188 : valid_0_4; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_989 = _GEN_215[7:6] == 2'h0 ? _GEN_189 : valid_0_5; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_990 = _GEN_215[7:6] == 2'h0 ? _GEN_190 : valid_0_6; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_991 = _GEN_215[7:6] == 2'h0 ? _GEN_191 : valid_0_7; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_992 = _GEN_215[7:6] == 2'h0 ? _GEN_192 : valid_0_8; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_993 = _GEN_215[7:6] == 2'h0 ? _GEN_193 : valid_0_9; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_994 = _GEN_215[7:6] == 2'h0 ? _GEN_194 : valid_0_10; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_995 = _GEN_215[7:6] == 2'h0 ? _GEN_195 : valid_0_11; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_996 = _GEN_215[7:6] == 2'h0 ? _GEN_196 : valid_0_12; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_997 = _GEN_215[7:6] == 2'h0 ? _GEN_197 : valid_0_13; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_998 = _GEN_215[7:6] == 2'h0 ? _GEN_198 : valid_0_14; // @[i_cache.scala 106:46 27:26]
  wire  _GEN_999 = _GEN_215[7:6] == 2'h0 ? _GEN_199 : valid_0_15; // @[i_cache.scala 106:46 27:26]
  wire [7:0] _GEN_1000 = _GEN_215[7:6] == 2'h0 ? _GEN_216 : _GEN_840; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1001 = _GEN_215[7:6] == 2'h0 ? _GEN_217 : _GEN_841; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1002 = _GEN_215[7:6] == 2'h0 ? _GEN_218 : _GEN_842; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1003 = _GEN_215[7:6] == 2'h0 ? _GEN_219 : _GEN_843; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1004 = _GEN_215[7:6] == 2'h0 ? _GEN_220 : _GEN_844; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1005 = _GEN_215[7:6] == 2'h0 ? _GEN_221 : _GEN_845; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1006 = _GEN_215[7:6] == 2'h0 ? _GEN_222 : _GEN_846; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1007 = _GEN_215[7:6] == 2'h0 ? _GEN_223 : _GEN_847; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1008 = _GEN_215[7:6] == 2'h0 ? _GEN_224 : _GEN_848; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1009 = _GEN_215[7:6] == 2'h0 ? _GEN_225 : _GEN_849; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1010 = _GEN_215[7:6] == 2'h0 ? _GEN_226 : _GEN_850; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1011 = _GEN_215[7:6] == 2'h0 ? _GEN_227 : _GEN_851; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1012 = _GEN_215[7:6] == 2'h0 ? _GEN_228 : _GEN_852; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1013 = _GEN_215[7:6] == 2'h0 ? _GEN_229 : _GEN_853; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1014 = _GEN_215[7:6] == 2'h0 ? _GEN_230 : _GEN_854; // @[i_cache.scala 106:46]
  wire [7:0] _GEN_1015 = _GEN_215[7:6] == 2'h0 ? _GEN_231 : _GEN_855; // @[i_cache.scala 106:46]
  wire [511:0] _GEN_1016 = _GEN_215[7:6] == 2'h0 ? ram_1_0 : _GEN_792; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1017 = _GEN_215[7:6] == 2'h0 ? ram_1_1 : _GEN_793; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1018 = _GEN_215[7:6] == 2'h0 ? ram_1_2 : _GEN_794; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1019 = _GEN_215[7:6] == 2'h0 ? ram_1_3 : _GEN_795; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1020 = _GEN_215[7:6] == 2'h0 ? ram_1_4 : _GEN_796; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1021 = _GEN_215[7:6] == 2'h0 ? ram_1_5 : _GEN_797; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1022 = _GEN_215[7:6] == 2'h0 ? ram_1_6 : _GEN_798; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1023 = _GEN_215[7:6] == 2'h0 ? ram_1_7 : _GEN_799; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1024 = _GEN_215[7:6] == 2'h0 ? ram_1_8 : _GEN_800; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1025 = _GEN_215[7:6] == 2'h0 ? ram_1_9 : _GEN_801; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1026 = _GEN_215[7:6] == 2'h0 ? ram_1_10 : _GEN_802; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1027 = _GEN_215[7:6] == 2'h0 ? ram_1_11 : _GEN_803; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1028 = _GEN_215[7:6] == 2'h0 ? ram_1_12 : _GEN_804; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1029 = _GEN_215[7:6] == 2'h0 ? ram_1_13 : _GEN_805; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1030 = _GEN_215[7:6] == 2'h0 ? ram_1_14 : _GEN_806; // @[i_cache.scala 106:46 20:24]
  wire [511:0] _GEN_1031 = _GEN_215[7:6] == 2'h0 ? ram_1_15 : _GEN_807; // @[i_cache.scala 106:46 20:24]
  wire [31:0] _GEN_1032 = _GEN_215[7:6] == 2'h0 ? tag_1_0 : _GEN_808; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1033 = _GEN_215[7:6] == 2'h0 ? tag_1_1 : _GEN_809; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1034 = _GEN_215[7:6] == 2'h0 ? tag_1_2 : _GEN_810; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1035 = _GEN_215[7:6] == 2'h0 ? tag_1_3 : _GEN_811; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1036 = _GEN_215[7:6] == 2'h0 ? tag_1_4 : _GEN_812; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1037 = _GEN_215[7:6] == 2'h0 ? tag_1_5 : _GEN_813; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1038 = _GEN_215[7:6] == 2'h0 ? tag_1_6 : _GEN_814; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1039 = _GEN_215[7:6] == 2'h0 ? tag_1_7 : _GEN_815; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1040 = _GEN_215[7:6] == 2'h0 ? tag_1_8 : _GEN_816; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1041 = _GEN_215[7:6] == 2'h0 ? tag_1_9 : _GEN_817; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1042 = _GEN_215[7:6] == 2'h0 ? tag_1_10 : _GEN_818; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1043 = _GEN_215[7:6] == 2'h0 ? tag_1_11 : _GEN_819; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1044 = _GEN_215[7:6] == 2'h0 ? tag_1_12 : _GEN_820; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1045 = _GEN_215[7:6] == 2'h0 ? tag_1_13 : _GEN_821; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1046 = _GEN_215[7:6] == 2'h0 ? tag_1_14 : _GEN_822; // @[i_cache.scala 106:46 24:24]
  wire [31:0] _GEN_1047 = _GEN_215[7:6] == 2'h0 ? tag_1_15 : _GEN_823; // @[i_cache.scala 106:46 24:24]
  wire  _GEN_1048 = _GEN_215[7:6] == 2'h0 ? valid_1_0 : _GEN_824; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1049 = _GEN_215[7:6] == 2'h0 ? valid_1_1 : _GEN_825; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1050 = _GEN_215[7:6] == 2'h0 ? valid_1_2 : _GEN_826; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1051 = _GEN_215[7:6] == 2'h0 ? valid_1_3 : _GEN_827; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1052 = _GEN_215[7:6] == 2'h0 ? valid_1_4 : _GEN_828; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1053 = _GEN_215[7:6] == 2'h0 ? valid_1_5 : _GEN_829; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1054 = _GEN_215[7:6] == 2'h0 ? valid_1_6 : _GEN_830; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1055 = _GEN_215[7:6] == 2'h0 ? valid_1_7 : _GEN_831; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1056 = _GEN_215[7:6] == 2'h0 ? valid_1_8 : _GEN_832; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1057 = _GEN_215[7:6] == 2'h0 ? valid_1_9 : _GEN_833; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1058 = _GEN_215[7:6] == 2'h0 ? valid_1_10 : _GEN_834; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1059 = _GEN_215[7:6] == 2'h0 ? valid_1_11 : _GEN_835; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1060 = _GEN_215[7:6] == 2'h0 ? valid_1_12 : _GEN_836; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1061 = _GEN_215[7:6] == 2'h0 ? valid_1_13 : _GEN_837; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1062 = _GEN_215[7:6] == 2'h0 ? valid_1_14 : _GEN_838; // @[i_cache.scala 106:46 28:26]
  wire  _GEN_1063 = _GEN_215[7:6] == 2'h0 ? valid_1_15 : _GEN_839; // @[i_cache.scala 106:46 28:26]
  wire [511:0] _GEN_1064 = _GEN_215[7:6] == 2'h0 ? ram_2_0 : _GEN_856; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1065 = _GEN_215[7:6] == 2'h0 ? ram_2_1 : _GEN_857; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1066 = _GEN_215[7:6] == 2'h0 ? ram_2_2 : _GEN_858; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1067 = _GEN_215[7:6] == 2'h0 ? ram_2_3 : _GEN_859; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1068 = _GEN_215[7:6] == 2'h0 ? ram_2_4 : _GEN_860; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1069 = _GEN_215[7:6] == 2'h0 ? ram_2_5 : _GEN_861; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1070 = _GEN_215[7:6] == 2'h0 ? ram_2_6 : _GEN_862; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1071 = _GEN_215[7:6] == 2'h0 ? ram_2_7 : _GEN_863; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1072 = _GEN_215[7:6] == 2'h0 ? ram_2_8 : _GEN_864; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1073 = _GEN_215[7:6] == 2'h0 ? ram_2_9 : _GEN_865; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1074 = _GEN_215[7:6] == 2'h0 ? ram_2_10 : _GEN_866; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1075 = _GEN_215[7:6] == 2'h0 ? ram_2_11 : _GEN_867; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1076 = _GEN_215[7:6] == 2'h0 ? ram_2_12 : _GEN_868; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1077 = _GEN_215[7:6] == 2'h0 ? ram_2_13 : _GEN_869; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1078 = _GEN_215[7:6] == 2'h0 ? ram_2_14 : _GEN_870; // @[i_cache.scala 106:46 21:24]
  wire [511:0] _GEN_1079 = _GEN_215[7:6] == 2'h0 ? ram_2_15 : _GEN_871; // @[i_cache.scala 106:46 21:24]
  wire [31:0] _GEN_1080 = _GEN_215[7:6] == 2'h0 ? tag_2_0 : _GEN_872; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1081 = _GEN_215[7:6] == 2'h0 ? tag_2_1 : _GEN_873; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1082 = _GEN_215[7:6] == 2'h0 ? tag_2_2 : _GEN_874; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1083 = _GEN_215[7:6] == 2'h0 ? tag_2_3 : _GEN_875; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1084 = _GEN_215[7:6] == 2'h0 ? tag_2_4 : _GEN_876; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1085 = _GEN_215[7:6] == 2'h0 ? tag_2_5 : _GEN_877; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1086 = _GEN_215[7:6] == 2'h0 ? tag_2_6 : _GEN_878; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1087 = _GEN_215[7:6] == 2'h0 ? tag_2_7 : _GEN_879; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1088 = _GEN_215[7:6] == 2'h0 ? tag_2_8 : _GEN_880; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1089 = _GEN_215[7:6] == 2'h0 ? tag_2_9 : _GEN_881; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1090 = _GEN_215[7:6] == 2'h0 ? tag_2_10 : _GEN_882; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1091 = _GEN_215[7:6] == 2'h0 ? tag_2_11 : _GEN_883; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1092 = _GEN_215[7:6] == 2'h0 ? tag_2_12 : _GEN_884; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1093 = _GEN_215[7:6] == 2'h0 ? tag_2_13 : _GEN_885; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1094 = _GEN_215[7:6] == 2'h0 ? tag_2_14 : _GEN_886; // @[i_cache.scala 106:46 25:24]
  wire [31:0] _GEN_1095 = _GEN_215[7:6] == 2'h0 ? tag_2_15 : _GEN_887; // @[i_cache.scala 106:46 25:24]
  wire  _GEN_1096 = _GEN_215[7:6] == 2'h0 ? valid_2_0 : _GEN_888; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1097 = _GEN_215[7:6] == 2'h0 ? valid_2_1 : _GEN_889; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1098 = _GEN_215[7:6] == 2'h0 ? valid_2_2 : _GEN_890; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1099 = _GEN_215[7:6] == 2'h0 ? valid_2_3 : _GEN_891; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1100 = _GEN_215[7:6] == 2'h0 ? valid_2_4 : _GEN_892; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1101 = _GEN_215[7:6] == 2'h0 ? valid_2_5 : _GEN_893; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1102 = _GEN_215[7:6] == 2'h0 ? valid_2_6 : _GEN_894; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1103 = _GEN_215[7:6] == 2'h0 ? valid_2_7 : _GEN_895; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1104 = _GEN_215[7:6] == 2'h0 ? valid_2_8 : _GEN_896; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1105 = _GEN_215[7:6] == 2'h0 ? valid_2_9 : _GEN_897; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1106 = _GEN_215[7:6] == 2'h0 ? valid_2_10 : _GEN_898; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1107 = _GEN_215[7:6] == 2'h0 ? valid_2_11 : _GEN_899; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1108 = _GEN_215[7:6] == 2'h0 ? valid_2_12 : _GEN_900; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1109 = _GEN_215[7:6] == 2'h0 ? valid_2_13 : _GEN_901; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1110 = _GEN_215[7:6] == 2'h0 ? valid_2_14 : _GEN_902; // @[i_cache.scala 106:46 29:26]
  wire  _GEN_1111 = _GEN_215[7:6] == 2'h0 ? valid_2_15 : _GEN_903; // @[i_cache.scala 106:46 29:26]
  wire [511:0] _GEN_1112 = _GEN_215[7:6] == 2'h0 ? ram_3_0 : _GEN_904; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1113 = _GEN_215[7:6] == 2'h0 ? ram_3_1 : _GEN_905; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1114 = _GEN_215[7:6] == 2'h0 ? ram_3_2 : _GEN_906; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1115 = _GEN_215[7:6] == 2'h0 ? ram_3_3 : _GEN_907; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1116 = _GEN_215[7:6] == 2'h0 ? ram_3_4 : _GEN_908; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1117 = _GEN_215[7:6] == 2'h0 ? ram_3_5 : _GEN_909; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1118 = _GEN_215[7:6] == 2'h0 ? ram_3_6 : _GEN_910; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1119 = _GEN_215[7:6] == 2'h0 ? ram_3_7 : _GEN_911; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1120 = _GEN_215[7:6] == 2'h0 ? ram_3_8 : _GEN_912; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1121 = _GEN_215[7:6] == 2'h0 ? ram_3_9 : _GEN_913; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1122 = _GEN_215[7:6] == 2'h0 ? ram_3_10 : _GEN_914; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1123 = _GEN_215[7:6] == 2'h0 ? ram_3_11 : _GEN_915; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1124 = _GEN_215[7:6] == 2'h0 ? ram_3_12 : _GEN_916; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1125 = _GEN_215[7:6] == 2'h0 ? ram_3_13 : _GEN_917; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1126 = _GEN_215[7:6] == 2'h0 ? ram_3_14 : _GEN_918; // @[i_cache.scala 106:46 22:24]
  wire [511:0] _GEN_1127 = _GEN_215[7:6] == 2'h0 ? ram_3_15 : _GEN_919; // @[i_cache.scala 106:46 22:24]
  wire [31:0] _GEN_1128 = _GEN_215[7:6] == 2'h0 ? tag_3_0 : _GEN_920; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1129 = _GEN_215[7:6] == 2'h0 ? tag_3_1 : _GEN_921; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1130 = _GEN_215[7:6] == 2'h0 ? tag_3_2 : _GEN_922; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1131 = _GEN_215[7:6] == 2'h0 ? tag_3_3 : _GEN_923; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1132 = _GEN_215[7:6] == 2'h0 ? tag_3_4 : _GEN_924; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1133 = _GEN_215[7:6] == 2'h0 ? tag_3_5 : _GEN_925; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1134 = _GEN_215[7:6] == 2'h0 ? tag_3_6 : _GEN_926; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1135 = _GEN_215[7:6] == 2'h0 ? tag_3_7 : _GEN_927; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1136 = _GEN_215[7:6] == 2'h0 ? tag_3_8 : _GEN_928; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1137 = _GEN_215[7:6] == 2'h0 ? tag_3_9 : _GEN_929; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1138 = _GEN_215[7:6] == 2'h0 ? tag_3_10 : _GEN_930; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1139 = _GEN_215[7:6] == 2'h0 ? tag_3_11 : _GEN_931; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1140 = _GEN_215[7:6] == 2'h0 ? tag_3_12 : _GEN_932; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1141 = _GEN_215[7:6] == 2'h0 ? tag_3_13 : _GEN_933; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1142 = _GEN_215[7:6] == 2'h0 ? tag_3_14 : _GEN_934; // @[i_cache.scala 106:46 26:24]
  wire [31:0] _GEN_1143 = _GEN_215[7:6] == 2'h0 ? tag_3_15 : _GEN_935; // @[i_cache.scala 106:46 26:24]
  wire  _GEN_1144 = _GEN_215[7:6] == 2'h0 ? valid_3_0 : _GEN_936; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1145 = _GEN_215[7:6] == 2'h0 ? valid_3_1 : _GEN_937; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1146 = _GEN_215[7:6] == 2'h0 ? valid_3_2 : _GEN_938; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1147 = _GEN_215[7:6] == 2'h0 ? valid_3_3 : _GEN_939; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1148 = _GEN_215[7:6] == 2'h0 ? valid_3_4 : _GEN_940; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1149 = _GEN_215[7:6] == 2'h0 ? valid_3_5 : _GEN_941; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1150 = _GEN_215[7:6] == 2'h0 ? valid_3_6 : _GEN_942; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1151 = _GEN_215[7:6] == 2'h0 ? valid_3_7 : _GEN_943; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1152 = _GEN_215[7:6] == 2'h0 ? valid_3_8 : _GEN_944; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1153 = _GEN_215[7:6] == 2'h0 ? valid_3_9 : _GEN_945; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1154 = _GEN_215[7:6] == 2'h0 ? valid_3_10 : _GEN_946; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1155 = _GEN_215[7:6] == 2'h0 ? valid_3_11 : _GEN_947; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1156 = _GEN_215[7:6] == 2'h0 ? valid_3_12 : _GEN_948; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1157 = _GEN_215[7:6] == 2'h0 ? valid_3_13 : _GEN_949; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1158 = _GEN_215[7:6] == 2'h0 ? valid_3_14 : _GEN_950; // @[i_cache.scala 106:46 30:26]
  wire  _GEN_1159 = _GEN_215[7:6] == 2'h0 ? valid_3_15 : _GEN_951; // @[i_cache.scala 106:46 30:26]
  wire [511:0] _GEN_1160 = unuse_way == 3'h4 ? _GEN_360 : _GEN_1112; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1161 = unuse_way == 3'h4 ? _GEN_361 : _GEN_1113; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1162 = unuse_way == 3'h4 ? _GEN_362 : _GEN_1114; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1163 = unuse_way == 3'h4 ? _GEN_363 : _GEN_1115; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1164 = unuse_way == 3'h4 ? _GEN_364 : _GEN_1116; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1165 = unuse_way == 3'h4 ? _GEN_365 : _GEN_1117; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1166 = unuse_way == 3'h4 ? _GEN_366 : _GEN_1118; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1167 = unuse_way == 3'h4 ? _GEN_367 : _GEN_1119; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1168 = unuse_way == 3'h4 ? _GEN_368 : _GEN_1120; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1169 = unuse_way == 3'h4 ? _GEN_369 : _GEN_1121; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1170 = unuse_way == 3'h4 ? _GEN_370 : _GEN_1122; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1171 = unuse_way == 3'h4 ? _GEN_371 : _GEN_1123; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1172 = unuse_way == 3'h4 ? _GEN_372 : _GEN_1124; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1173 = unuse_way == 3'h4 ? _GEN_373 : _GEN_1125; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1174 = unuse_way == 3'h4 ? _GEN_374 : _GEN_1126; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1175 = unuse_way == 3'h4 ? _GEN_375 : _GEN_1127; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1176 = unuse_way == 3'h4 ? _GEN_376 : _GEN_1128; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1177 = unuse_way == 3'h4 ? _GEN_377 : _GEN_1129; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1178 = unuse_way == 3'h4 ? _GEN_378 : _GEN_1130; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1179 = unuse_way == 3'h4 ? _GEN_379 : _GEN_1131; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1180 = unuse_way == 3'h4 ? _GEN_380 : _GEN_1132; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1181 = unuse_way == 3'h4 ? _GEN_381 : _GEN_1133; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1182 = unuse_way == 3'h4 ? _GEN_382 : _GEN_1134; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1183 = unuse_way == 3'h4 ? _GEN_383 : _GEN_1135; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1184 = unuse_way == 3'h4 ? _GEN_384 : _GEN_1136; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1185 = unuse_way == 3'h4 ? _GEN_385 : _GEN_1137; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1186 = unuse_way == 3'h4 ? _GEN_386 : _GEN_1138; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1187 = unuse_way == 3'h4 ? _GEN_387 : _GEN_1139; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1188 = unuse_way == 3'h4 ? _GEN_388 : _GEN_1140; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1189 = unuse_way == 3'h4 ? _GEN_389 : _GEN_1141; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1190 = unuse_way == 3'h4 ? _GEN_390 : _GEN_1142; // @[i_cache.scala 100:40]
  wire [31:0] _GEN_1191 = unuse_way == 3'h4 ? _GEN_391 : _GEN_1143; // @[i_cache.scala 100:40]
  wire  _GEN_1192 = unuse_way == 3'h4 ? _GEN_392 : _GEN_1144; // @[i_cache.scala 100:40]
  wire  _GEN_1193 = unuse_way == 3'h4 ? _GEN_393 : _GEN_1145; // @[i_cache.scala 100:40]
  wire  _GEN_1194 = unuse_way == 3'h4 ? _GEN_394 : _GEN_1146; // @[i_cache.scala 100:40]
  wire  _GEN_1195 = unuse_way == 3'h4 ? _GEN_395 : _GEN_1147; // @[i_cache.scala 100:40]
  wire  _GEN_1196 = unuse_way == 3'h4 ? _GEN_396 : _GEN_1148; // @[i_cache.scala 100:40]
  wire  _GEN_1197 = unuse_way == 3'h4 ? _GEN_397 : _GEN_1149; // @[i_cache.scala 100:40]
  wire  _GEN_1198 = unuse_way == 3'h4 ? _GEN_398 : _GEN_1150; // @[i_cache.scala 100:40]
  wire  _GEN_1199 = unuse_way == 3'h4 ? _GEN_399 : _GEN_1151; // @[i_cache.scala 100:40]
  wire  _GEN_1200 = unuse_way == 3'h4 ? _GEN_400 : _GEN_1152; // @[i_cache.scala 100:40]
  wire  _GEN_1201 = unuse_way == 3'h4 ? _GEN_401 : _GEN_1153; // @[i_cache.scala 100:40]
  wire  _GEN_1202 = unuse_way == 3'h4 ? _GEN_402 : _GEN_1154; // @[i_cache.scala 100:40]
  wire  _GEN_1203 = unuse_way == 3'h4 ? _GEN_403 : _GEN_1155; // @[i_cache.scala 100:40]
  wire  _GEN_1204 = unuse_way == 3'h4 ? _GEN_404 : _GEN_1156; // @[i_cache.scala 100:40]
  wire  _GEN_1205 = unuse_way == 3'h4 ? _GEN_405 : _GEN_1157; // @[i_cache.scala 100:40]
  wire  _GEN_1206 = unuse_way == 3'h4 ? _GEN_406 : _GEN_1158; // @[i_cache.scala 100:40]
  wire  _GEN_1207 = unuse_way == 3'h4 ? _GEN_407 : _GEN_1159; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1208 = unuse_way == 3'h4 ? _GEN_408 : _GEN_1000; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1209 = unuse_way == 3'h4 ? _GEN_409 : _GEN_1001; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1210 = unuse_way == 3'h4 ? _GEN_410 : _GEN_1002; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1211 = unuse_way == 3'h4 ? _GEN_411 : _GEN_1003; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1212 = unuse_way == 3'h4 ? _GEN_412 : _GEN_1004; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1213 = unuse_way == 3'h4 ? _GEN_413 : _GEN_1005; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1214 = unuse_way == 3'h4 ? _GEN_414 : _GEN_1006; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1215 = unuse_way == 3'h4 ? _GEN_415 : _GEN_1007; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1216 = unuse_way == 3'h4 ? _GEN_416 : _GEN_1008; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1217 = unuse_way == 3'h4 ? _GEN_417 : _GEN_1009; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1218 = unuse_way == 3'h4 ? _GEN_418 : _GEN_1010; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1219 = unuse_way == 3'h4 ? _GEN_419 : _GEN_1011; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1220 = unuse_way == 3'h4 ? _GEN_420 : _GEN_1012; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1221 = unuse_way == 3'h4 ? _GEN_421 : _GEN_1013; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1222 = unuse_way == 3'h4 ? _GEN_422 : _GEN_1014; // @[i_cache.scala 100:40]
  wire [7:0] _GEN_1223 = unuse_way == 3'h4 ? _GEN_423 : _GEN_1015; // @[i_cache.scala 100:40]
  wire [511:0] _GEN_1224 = unuse_way == 3'h4 ? ram_0_0 : _GEN_952; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1225 = unuse_way == 3'h4 ? ram_0_1 : _GEN_953; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1226 = unuse_way == 3'h4 ? ram_0_2 : _GEN_954; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1227 = unuse_way == 3'h4 ? ram_0_3 : _GEN_955; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1228 = unuse_way == 3'h4 ? ram_0_4 : _GEN_956; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1229 = unuse_way == 3'h4 ? ram_0_5 : _GEN_957; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1230 = unuse_way == 3'h4 ? ram_0_6 : _GEN_958; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1231 = unuse_way == 3'h4 ? ram_0_7 : _GEN_959; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1232 = unuse_way == 3'h4 ? ram_0_8 : _GEN_960; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1233 = unuse_way == 3'h4 ? ram_0_9 : _GEN_961; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1234 = unuse_way == 3'h4 ? ram_0_10 : _GEN_962; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1235 = unuse_way == 3'h4 ? ram_0_11 : _GEN_963; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1236 = unuse_way == 3'h4 ? ram_0_12 : _GEN_964; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1237 = unuse_way == 3'h4 ? ram_0_13 : _GEN_965; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1238 = unuse_way == 3'h4 ? ram_0_14 : _GEN_966; // @[i_cache.scala 100:40 19:24]
  wire [511:0] _GEN_1239 = unuse_way == 3'h4 ? ram_0_15 : _GEN_967; // @[i_cache.scala 100:40 19:24]
  wire [31:0] _GEN_1240 = unuse_way == 3'h4 ? tag_0_0 : _GEN_968; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1241 = unuse_way == 3'h4 ? tag_0_1 : _GEN_969; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1242 = unuse_way == 3'h4 ? tag_0_2 : _GEN_970; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1243 = unuse_way == 3'h4 ? tag_0_3 : _GEN_971; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1244 = unuse_way == 3'h4 ? tag_0_4 : _GEN_972; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1245 = unuse_way == 3'h4 ? tag_0_5 : _GEN_973; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1246 = unuse_way == 3'h4 ? tag_0_6 : _GEN_974; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1247 = unuse_way == 3'h4 ? tag_0_7 : _GEN_975; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1248 = unuse_way == 3'h4 ? tag_0_8 : _GEN_976; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1249 = unuse_way == 3'h4 ? tag_0_9 : _GEN_977; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1250 = unuse_way == 3'h4 ? tag_0_10 : _GEN_978; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1251 = unuse_way == 3'h4 ? tag_0_11 : _GEN_979; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1252 = unuse_way == 3'h4 ? tag_0_12 : _GEN_980; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1253 = unuse_way == 3'h4 ? tag_0_13 : _GEN_981; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1254 = unuse_way == 3'h4 ? tag_0_14 : _GEN_982; // @[i_cache.scala 100:40 23:24]
  wire [31:0] _GEN_1255 = unuse_way == 3'h4 ? tag_0_15 : _GEN_983; // @[i_cache.scala 100:40 23:24]
  wire  _GEN_1256 = unuse_way == 3'h4 ? valid_0_0 : _GEN_984; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1257 = unuse_way == 3'h4 ? valid_0_1 : _GEN_985; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1258 = unuse_way == 3'h4 ? valid_0_2 : _GEN_986; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1259 = unuse_way == 3'h4 ? valid_0_3 : _GEN_987; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1260 = unuse_way == 3'h4 ? valid_0_4 : _GEN_988; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1261 = unuse_way == 3'h4 ? valid_0_5 : _GEN_989; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1262 = unuse_way == 3'h4 ? valid_0_6 : _GEN_990; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1263 = unuse_way == 3'h4 ? valid_0_7 : _GEN_991; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1264 = unuse_way == 3'h4 ? valid_0_8 : _GEN_992; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1265 = unuse_way == 3'h4 ? valid_0_9 : _GEN_993; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1266 = unuse_way == 3'h4 ? valid_0_10 : _GEN_994; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1267 = unuse_way == 3'h4 ? valid_0_11 : _GEN_995; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1268 = unuse_way == 3'h4 ? valid_0_12 : _GEN_996; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1269 = unuse_way == 3'h4 ? valid_0_13 : _GEN_997; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1270 = unuse_way == 3'h4 ? valid_0_14 : _GEN_998; // @[i_cache.scala 100:40 27:26]
  wire  _GEN_1271 = unuse_way == 3'h4 ? valid_0_15 : _GEN_999; // @[i_cache.scala 100:40 27:26]
  wire [511:0] _GEN_1272 = unuse_way == 3'h4 ? ram_1_0 : _GEN_1016; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1273 = unuse_way == 3'h4 ? ram_1_1 : _GEN_1017; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1274 = unuse_way == 3'h4 ? ram_1_2 : _GEN_1018; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1275 = unuse_way == 3'h4 ? ram_1_3 : _GEN_1019; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1276 = unuse_way == 3'h4 ? ram_1_4 : _GEN_1020; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1277 = unuse_way == 3'h4 ? ram_1_5 : _GEN_1021; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1278 = unuse_way == 3'h4 ? ram_1_6 : _GEN_1022; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1279 = unuse_way == 3'h4 ? ram_1_7 : _GEN_1023; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1280 = unuse_way == 3'h4 ? ram_1_8 : _GEN_1024; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1281 = unuse_way == 3'h4 ? ram_1_9 : _GEN_1025; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1282 = unuse_way == 3'h4 ? ram_1_10 : _GEN_1026; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1283 = unuse_way == 3'h4 ? ram_1_11 : _GEN_1027; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1284 = unuse_way == 3'h4 ? ram_1_12 : _GEN_1028; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1285 = unuse_way == 3'h4 ? ram_1_13 : _GEN_1029; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1286 = unuse_way == 3'h4 ? ram_1_14 : _GEN_1030; // @[i_cache.scala 100:40 20:24]
  wire [511:0] _GEN_1287 = unuse_way == 3'h4 ? ram_1_15 : _GEN_1031; // @[i_cache.scala 100:40 20:24]
  wire [31:0] _GEN_1288 = unuse_way == 3'h4 ? tag_1_0 : _GEN_1032; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1289 = unuse_way == 3'h4 ? tag_1_1 : _GEN_1033; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1290 = unuse_way == 3'h4 ? tag_1_2 : _GEN_1034; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1291 = unuse_way == 3'h4 ? tag_1_3 : _GEN_1035; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1292 = unuse_way == 3'h4 ? tag_1_4 : _GEN_1036; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1293 = unuse_way == 3'h4 ? tag_1_5 : _GEN_1037; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1294 = unuse_way == 3'h4 ? tag_1_6 : _GEN_1038; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1295 = unuse_way == 3'h4 ? tag_1_7 : _GEN_1039; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1296 = unuse_way == 3'h4 ? tag_1_8 : _GEN_1040; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1297 = unuse_way == 3'h4 ? tag_1_9 : _GEN_1041; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1298 = unuse_way == 3'h4 ? tag_1_10 : _GEN_1042; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1299 = unuse_way == 3'h4 ? tag_1_11 : _GEN_1043; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1300 = unuse_way == 3'h4 ? tag_1_12 : _GEN_1044; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1301 = unuse_way == 3'h4 ? tag_1_13 : _GEN_1045; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1302 = unuse_way == 3'h4 ? tag_1_14 : _GEN_1046; // @[i_cache.scala 100:40 24:24]
  wire [31:0] _GEN_1303 = unuse_way == 3'h4 ? tag_1_15 : _GEN_1047; // @[i_cache.scala 100:40 24:24]
  wire  _GEN_1304 = unuse_way == 3'h4 ? valid_1_0 : _GEN_1048; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1305 = unuse_way == 3'h4 ? valid_1_1 : _GEN_1049; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1306 = unuse_way == 3'h4 ? valid_1_2 : _GEN_1050; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1307 = unuse_way == 3'h4 ? valid_1_3 : _GEN_1051; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1308 = unuse_way == 3'h4 ? valid_1_4 : _GEN_1052; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1309 = unuse_way == 3'h4 ? valid_1_5 : _GEN_1053; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1310 = unuse_way == 3'h4 ? valid_1_6 : _GEN_1054; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1311 = unuse_way == 3'h4 ? valid_1_7 : _GEN_1055; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1312 = unuse_way == 3'h4 ? valid_1_8 : _GEN_1056; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1313 = unuse_way == 3'h4 ? valid_1_9 : _GEN_1057; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1314 = unuse_way == 3'h4 ? valid_1_10 : _GEN_1058; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1315 = unuse_way == 3'h4 ? valid_1_11 : _GEN_1059; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1316 = unuse_way == 3'h4 ? valid_1_12 : _GEN_1060; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1317 = unuse_way == 3'h4 ? valid_1_13 : _GEN_1061; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1318 = unuse_way == 3'h4 ? valid_1_14 : _GEN_1062; // @[i_cache.scala 100:40 28:26]
  wire  _GEN_1319 = unuse_way == 3'h4 ? valid_1_15 : _GEN_1063; // @[i_cache.scala 100:40 28:26]
  wire [511:0] _GEN_1320 = unuse_way == 3'h4 ? ram_2_0 : _GEN_1064; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1321 = unuse_way == 3'h4 ? ram_2_1 : _GEN_1065; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1322 = unuse_way == 3'h4 ? ram_2_2 : _GEN_1066; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1323 = unuse_way == 3'h4 ? ram_2_3 : _GEN_1067; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1324 = unuse_way == 3'h4 ? ram_2_4 : _GEN_1068; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1325 = unuse_way == 3'h4 ? ram_2_5 : _GEN_1069; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1326 = unuse_way == 3'h4 ? ram_2_6 : _GEN_1070; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1327 = unuse_way == 3'h4 ? ram_2_7 : _GEN_1071; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1328 = unuse_way == 3'h4 ? ram_2_8 : _GEN_1072; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1329 = unuse_way == 3'h4 ? ram_2_9 : _GEN_1073; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1330 = unuse_way == 3'h4 ? ram_2_10 : _GEN_1074; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1331 = unuse_way == 3'h4 ? ram_2_11 : _GEN_1075; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1332 = unuse_way == 3'h4 ? ram_2_12 : _GEN_1076; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1333 = unuse_way == 3'h4 ? ram_2_13 : _GEN_1077; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1334 = unuse_way == 3'h4 ? ram_2_14 : _GEN_1078; // @[i_cache.scala 100:40 21:24]
  wire [511:0] _GEN_1335 = unuse_way == 3'h4 ? ram_2_15 : _GEN_1079; // @[i_cache.scala 100:40 21:24]
  wire [31:0] _GEN_1336 = unuse_way == 3'h4 ? tag_2_0 : _GEN_1080; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1337 = unuse_way == 3'h4 ? tag_2_1 : _GEN_1081; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1338 = unuse_way == 3'h4 ? tag_2_2 : _GEN_1082; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1339 = unuse_way == 3'h4 ? tag_2_3 : _GEN_1083; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1340 = unuse_way == 3'h4 ? tag_2_4 : _GEN_1084; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1341 = unuse_way == 3'h4 ? tag_2_5 : _GEN_1085; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1342 = unuse_way == 3'h4 ? tag_2_6 : _GEN_1086; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1343 = unuse_way == 3'h4 ? tag_2_7 : _GEN_1087; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1344 = unuse_way == 3'h4 ? tag_2_8 : _GEN_1088; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1345 = unuse_way == 3'h4 ? tag_2_9 : _GEN_1089; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1346 = unuse_way == 3'h4 ? tag_2_10 : _GEN_1090; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1347 = unuse_way == 3'h4 ? tag_2_11 : _GEN_1091; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1348 = unuse_way == 3'h4 ? tag_2_12 : _GEN_1092; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1349 = unuse_way == 3'h4 ? tag_2_13 : _GEN_1093; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1350 = unuse_way == 3'h4 ? tag_2_14 : _GEN_1094; // @[i_cache.scala 100:40 25:24]
  wire [31:0] _GEN_1351 = unuse_way == 3'h4 ? tag_2_15 : _GEN_1095; // @[i_cache.scala 100:40 25:24]
  wire  _GEN_1352 = unuse_way == 3'h4 ? valid_2_0 : _GEN_1096; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1353 = unuse_way == 3'h4 ? valid_2_1 : _GEN_1097; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1354 = unuse_way == 3'h4 ? valid_2_2 : _GEN_1098; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1355 = unuse_way == 3'h4 ? valid_2_3 : _GEN_1099; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1356 = unuse_way == 3'h4 ? valid_2_4 : _GEN_1100; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1357 = unuse_way == 3'h4 ? valid_2_5 : _GEN_1101; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1358 = unuse_way == 3'h4 ? valid_2_6 : _GEN_1102; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1359 = unuse_way == 3'h4 ? valid_2_7 : _GEN_1103; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1360 = unuse_way == 3'h4 ? valid_2_8 : _GEN_1104; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1361 = unuse_way == 3'h4 ? valid_2_9 : _GEN_1105; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1362 = unuse_way == 3'h4 ? valid_2_10 : _GEN_1106; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1363 = unuse_way == 3'h4 ? valid_2_11 : _GEN_1107; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1364 = unuse_way == 3'h4 ? valid_2_12 : _GEN_1108; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1365 = unuse_way == 3'h4 ? valid_2_13 : _GEN_1109; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1366 = unuse_way == 3'h4 ? valid_2_14 : _GEN_1110; // @[i_cache.scala 100:40 29:26]
  wire  _GEN_1367 = unuse_way == 3'h4 ? valid_2_15 : _GEN_1111; // @[i_cache.scala 100:40 29:26]
  wire [511:0] _GEN_1368 = unuse_way == 3'h3 ? _GEN_296 : _GEN_1320; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1369 = unuse_way == 3'h3 ? _GEN_297 : _GEN_1321; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1370 = unuse_way == 3'h3 ? _GEN_298 : _GEN_1322; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1371 = unuse_way == 3'h3 ? _GEN_299 : _GEN_1323; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1372 = unuse_way == 3'h3 ? _GEN_300 : _GEN_1324; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1373 = unuse_way == 3'h3 ? _GEN_301 : _GEN_1325; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1374 = unuse_way == 3'h3 ? _GEN_302 : _GEN_1326; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1375 = unuse_way == 3'h3 ? _GEN_303 : _GEN_1327; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1376 = unuse_way == 3'h3 ? _GEN_304 : _GEN_1328; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1377 = unuse_way == 3'h3 ? _GEN_305 : _GEN_1329; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1378 = unuse_way == 3'h3 ? _GEN_306 : _GEN_1330; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1379 = unuse_way == 3'h3 ? _GEN_307 : _GEN_1331; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1380 = unuse_way == 3'h3 ? _GEN_308 : _GEN_1332; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1381 = unuse_way == 3'h3 ? _GEN_309 : _GEN_1333; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1382 = unuse_way == 3'h3 ? _GEN_310 : _GEN_1334; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1383 = unuse_way == 3'h3 ? _GEN_311 : _GEN_1335; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1384 = unuse_way == 3'h3 ? _GEN_312 : _GEN_1336; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1385 = unuse_way == 3'h3 ? _GEN_313 : _GEN_1337; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1386 = unuse_way == 3'h3 ? _GEN_314 : _GEN_1338; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1387 = unuse_way == 3'h3 ? _GEN_315 : _GEN_1339; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1388 = unuse_way == 3'h3 ? _GEN_316 : _GEN_1340; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1389 = unuse_way == 3'h3 ? _GEN_317 : _GEN_1341; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1390 = unuse_way == 3'h3 ? _GEN_318 : _GEN_1342; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1391 = unuse_way == 3'h3 ? _GEN_319 : _GEN_1343; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1392 = unuse_way == 3'h3 ? _GEN_320 : _GEN_1344; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1393 = unuse_way == 3'h3 ? _GEN_321 : _GEN_1345; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1394 = unuse_way == 3'h3 ? _GEN_322 : _GEN_1346; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1395 = unuse_way == 3'h3 ? _GEN_323 : _GEN_1347; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1396 = unuse_way == 3'h3 ? _GEN_324 : _GEN_1348; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1397 = unuse_way == 3'h3 ? _GEN_325 : _GEN_1349; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1398 = unuse_way == 3'h3 ? _GEN_326 : _GEN_1350; // @[i_cache.scala 95:40]
  wire [31:0] _GEN_1399 = unuse_way == 3'h3 ? _GEN_327 : _GEN_1351; // @[i_cache.scala 95:40]
  wire  _GEN_1400 = unuse_way == 3'h3 ? _GEN_328 : _GEN_1352; // @[i_cache.scala 95:40]
  wire  _GEN_1401 = unuse_way == 3'h3 ? _GEN_329 : _GEN_1353; // @[i_cache.scala 95:40]
  wire  _GEN_1402 = unuse_way == 3'h3 ? _GEN_330 : _GEN_1354; // @[i_cache.scala 95:40]
  wire  _GEN_1403 = unuse_way == 3'h3 ? _GEN_331 : _GEN_1355; // @[i_cache.scala 95:40]
  wire  _GEN_1404 = unuse_way == 3'h3 ? _GEN_332 : _GEN_1356; // @[i_cache.scala 95:40]
  wire  _GEN_1405 = unuse_way == 3'h3 ? _GEN_333 : _GEN_1357; // @[i_cache.scala 95:40]
  wire  _GEN_1406 = unuse_way == 3'h3 ? _GEN_334 : _GEN_1358; // @[i_cache.scala 95:40]
  wire  _GEN_1407 = unuse_way == 3'h3 ? _GEN_335 : _GEN_1359; // @[i_cache.scala 95:40]
  wire  _GEN_1408 = unuse_way == 3'h3 ? _GEN_336 : _GEN_1360; // @[i_cache.scala 95:40]
  wire  _GEN_1409 = unuse_way == 3'h3 ? _GEN_337 : _GEN_1361; // @[i_cache.scala 95:40]
  wire  _GEN_1410 = unuse_way == 3'h3 ? _GEN_338 : _GEN_1362; // @[i_cache.scala 95:40]
  wire  _GEN_1411 = unuse_way == 3'h3 ? _GEN_339 : _GEN_1363; // @[i_cache.scala 95:40]
  wire  _GEN_1412 = unuse_way == 3'h3 ? _GEN_340 : _GEN_1364; // @[i_cache.scala 95:40]
  wire  _GEN_1413 = unuse_way == 3'h3 ? _GEN_341 : _GEN_1365; // @[i_cache.scala 95:40]
  wire  _GEN_1414 = unuse_way == 3'h3 ? _GEN_342 : _GEN_1366; // @[i_cache.scala 95:40]
  wire  _GEN_1415 = unuse_way == 3'h3 ? _GEN_343 : _GEN_1367; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1416 = unuse_way == 3'h3 ? _GEN_344 : _GEN_1208; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1417 = unuse_way == 3'h3 ? _GEN_345 : _GEN_1209; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1418 = unuse_way == 3'h3 ? _GEN_346 : _GEN_1210; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1419 = unuse_way == 3'h3 ? _GEN_347 : _GEN_1211; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1420 = unuse_way == 3'h3 ? _GEN_348 : _GEN_1212; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1421 = unuse_way == 3'h3 ? _GEN_349 : _GEN_1213; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1422 = unuse_way == 3'h3 ? _GEN_350 : _GEN_1214; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1423 = unuse_way == 3'h3 ? _GEN_351 : _GEN_1215; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1424 = unuse_way == 3'h3 ? _GEN_352 : _GEN_1216; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1425 = unuse_way == 3'h3 ? _GEN_353 : _GEN_1217; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1426 = unuse_way == 3'h3 ? _GEN_354 : _GEN_1218; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1427 = unuse_way == 3'h3 ? _GEN_355 : _GEN_1219; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1428 = unuse_way == 3'h3 ? _GEN_356 : _GEN_1220; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1429 = unuse_way == 3'h3 ? _GEN_357 : _GEN_1221; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1430 = unuse_way == 3'h3 ? _GEN_358 : _GEN_1222; // @[i_cache.scala 95:40]
  wire [7:0] _GEN_1431 = unuse_way == 3'h3 ? _GEN_359 : _GEN_1223; // @[i_cache.scala 95:40]
  wire [511:0] _GEN_1432 = unuse_way == 3'h3 ? ram_3_0 : _GEN_1160; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1433 = unuse_way == 3'h3 ? ram_3_1 : _GEN_1161; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1434 = unuse_way == 3'h3 ? ram_3_2 : _GEN_1162; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1435 = unuse_way == 3'h3 ? ram_3_3 : _GEN_1163; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1436 = unuse_way == 3'h3 ? ram_3_4 : _GEN_1164; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1437 = unuse_way == 3'h3 ? ram_3_5 : _GEN_1165; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1438 = unuse_way == 3'h3 ? ram_3_6 : _GEN_1166; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1439 = unuse_way == 3'h3 ? ram_3_7 : _GEN_1167; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1440 = unuse_way == 3'h3 ? ram_3_8 : _GEN_1168; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1441 = unuse_way == 3'h3 ? ram_3_9 : _GEN_1169; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1442 = unuse_way == 3'h3 ? ram_3_10 : _GEN_1170; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1443 = unuse_way == 3'h3 ? ram_3_11 : _GEN_1171; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1444 = unuse_way == 3'h3 ? ram_3_12 : _GEN_1172; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1445 = unuse_way == 3'h3 ? ram_3_13 : _GEN_1173; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1446 = unuse_way == 3'h3 ? ram_3_14 : _GEN_1174; // @[i_cache.scala 22:24 95:40]
  wire [511:0] _GEN_1447 = unuse_way == 3'h3 ? ram_3_15 : _GEN_1175; // @[i_cache.scala 22:24 95:40]
  wire [31:0] _GEN_1448 = unuse_way == 3'h3 ? tag_3_0 : _GEN_1176; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1449 = unuse_way == 3'h3 ? tag_3_1 : _GEN_1177; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1450 = unuse_way == 3'h3 ? tag_3_2 : _GEN_1178; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1451 = unuse_way == 3'h3 ? tag_3_3 : _GEN_1179; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1452 = unuse_way == 3'h3 ? tag_3_4 : _GEN_1180; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1453 = unuse_way == 3'h3 ? tag_3_5 : _GEN_1181; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1454 = unuse_way == 3'h3 ? tag_3_6 : _GEN_1182; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1455 = unuse_way == 3'h3 ? tag_3_7 : _GEN_1183; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1456 = unuse_way == 3'h3 ? tag_3_8 : _GEN_1184; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1457 = unuse_way == 3'h3 ? tag_3_9 : _GEN_1185; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1458 = unuse_way == 3'h3 ? tag_3_10 : _GEN_1186; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1459 = unuse_way == 3'h3 ? tag_3_11 : _GEN_1187; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1460 = unuse_way == 3'h3 ? tag_3_12 : _GEN_1188; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1461 = unuse_way == 3'h3 ? tag_3_13 : _GEN_1189; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1462 = unuse_way == 3'h3 ? tag_3_14 : _GEN_1190; // @[i_cache.scala 26:24 95:40]
  wire [31:0] _GEN_1463 = unuse_way == 3'h3 ? tag_3_15 : _GEN_1191; // @[i_cache.scala 26:24 95:40]
  wire  _GEN_1464 = unuse_way == 3'h3 ? valid_3_0 : _GEN_1192; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1465 = unuse_way == 3'h3 ? valid_3_1 : _GEN_1193; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1466 = unuse_way == 3'h3 ? valid_3_2 : _GEN_1194; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1467 = unuse_way == 3'h3 ? valid_3_3 : _GEN_1195; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1468 = unuse_way == 3'h3 ? valid_3_4 : _GEN_1196; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1469 = unuse_way == 3'h3 ? valid_3_5 : _GEN_1197; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1470 = unuse_way == 3'h3 ? valid_3_6 : _GEN_1198; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1471 = unuse_way == 3'h3 ? valid_3_7 : _GEN_1199; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1472 = unuse_way == 3'h3 ? valid_3_8 : _GEN_1200; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1473 = unuse_way == 3'h3 ? valid_3_9 : _GEN_1201; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1474 = unuse_way == 3'h3 ? valid_3_10 : _GEN_1202; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1475 = unuse_way == 3'h3 ? valid_3_11 : _GEN_1203; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1476 = unuse_way == 3'h3 ? valid_3_12 : _GEN_1204; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1477 = unuse_way == 3'h3 ? valid_3_13 : _GEN_1205; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1478 = unuse_way == 3'h3 ? valid_3_14 : _GEN_1206; // @[i_cache.scala 30:26 95:40]
  wire  _GEN_1479 = unuse_way == 3'h3 ? valid_3_15 : _GEN_1207; // @[i_cache.scala 30:26 95:40]
  wire [511:0] _GEN_1480 = unuse_way == 3'h3 ? ram_0_0 : _GEN_1224; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1481 = unuse_way == 3'h3 ? ram_0_1 : _GEN_1225; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1482 = unuse_way == 3'h3 ? ram_0_2 : _GEN_1226; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1483 = unuse_way == 3'h3 ? ram_0_3 : _GEN_1227; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1484 = unuse_way == 3'h3 ? ram_0_4 : _GEN_1228; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1485 = unuse_way == 3'h3 ? ram_0_5 : _GEN_1229; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1486 = unuse_way == 3'h3 ? ram_0_6 : _GEN_1230; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1487 = unuse_way == 3'h3 ? ram_0_7 : _GEN_1231; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1488 = unuse_way == 3'h3 ? ram_0_8 : _GEN_1232; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1489 = unuse_way == 3'h3 ? ram_0_9 : _GEN_1233; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1490 = unuse_way == 3'h3 ? ram_0_10 : _GEN_1234; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1491 = unuse_way == 3'h3 ? ram_0_11 : _GEN_1235; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1492 = unuse_way == 3'h3 ? ram_0_12 : _GEN_1236; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1493 = unuse_way == 3'h3 ? ram_0_13 : _GEN_1237; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1494 = unuse_way == 3'h3 ? ram_0_14 : _GEN_1238; // @[i_cache.scala 19:24 95:40]
  wire [511:0] _GEN_1495 = unuse_way == 3'h3 ? ram_0_15 : _GEN_1239; // @[i_cache.scala 19:24 95:40]
  wire [31:0] _GEN_1496 = unuse_way == 3'h3 ? tag_0_0 : _GEN_1240; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1497 = unuse_way == 3'h3 ? tag_0_1 : _GEN_1241; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1498 = unuse_way == 3'h3 ? tag_0_2 : _GEN_1242; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1499 = unuse_way == 3'h3 ? tag_0_3 : _GEN_1243; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1500 = unuse_way == 3'h3 ? tag_0_4 : _GEN_1244; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1501 = unuse_way == 3'h3 ? tag_0_5 : _GEN_1245; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1502 = unuse_way == 3'h3 ? tag_0_6 : _GEN_1246; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1503 = unuse_way == 3'h3 ? tag_0_7 : _GEN_1247; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1504 = unuse_way == 3'h3 ? tag_0_8 : _GEN_1248; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1505 = unuse_way == 3'h3 ? tag_0_9 : _GEN_1249; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1506 = unuse_way == 3'h3 ? tag_0_10 : _GEN_1250; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1507 = unuse_way == 3'h3 ? tag_0_11 : _GEN_1251; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1508 = unuse_way == 3'h3 ? tag_0_12 : _GEN_1252; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1509 = unuse_way == 3'h3 ? tag_0_13 : _GEN_1253; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1510 = unuse_way == 3'h3 ? tag_0_14 : _GEN_1254; // @[i_cache.scala 23:24 95:40]
  wire [31:0] _GEN_1511 = unuse_way == 3'h3 ? tag_0_15 : _GEN_1255; // @[i_cache.scala 23:24 95:40]
  wire  _GEN_1512 = unuse_way == 3'h3 ? valid_0_0 : _GEN_1256; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1513 = unuse_way == 3'h3 ? valid_0_1 : _GEN_1257; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1514 = unuse_way == 3'h3 ? valid_0_2 : _GEN_1258; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1515 = unuse_way == 3'h3 ? valid_0_3 : _GEN_1259; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1516 = unuse_way == 3'h3 ? valid_0_4 : _GEN_1260; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1517 = unuse_way == 3'h3 ? valid_0_5 : _GEN_1261; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1518 = unuse_way == 3'h3 ? valid_0_6 : _GEN_1262; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1519 = unuse_way == 3'h3 ? valid_0_7 : _GEN_1263; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1520 = unuse_way == 3'h3 ? valid_0_8 : _GEN_1264; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1521 = unuse_way == 3'h3 ? valid_0_9 : _GEN_1265; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1522 = unuse_way == 3'h3 ? valid_0_10 : _GEN_1266; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1523 = unuse_way == 3'h3 ? valid_0_11 : _GEN_1267; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1524 = unuse_way == 3'h3 ? valid_0_12 : _GEN_1268; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1525 = unuse_way == 3'h3 ? valid_0_13 : _GEN_1269; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1526 = unuse_way == 3'h3 ? valid_0_14 : _GEN_1270; // @[i_cache.scala 27:26 95:40]
  wire  _GEN_1527 = unuse_way == 3'h3 ? valid_0_15 : _GEN_1271; // @[i_cache.scala 27:26 95:40]
  wire [511:0] _GEN_1528 = unuse_way == 3'h3 ? ram_1_0 : _GEN_1272; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1529 = unuse_way == 3'h3 ? ram_1_1 : _GEN_1273; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1530 = unuse_way == 3'h3 ? ram_1_2 : _GEN_1274; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1531 = unuse_way == 3'h3 ? ram_1_3 : _GEN_1275; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1532 = unuse_way == 3'h3 ? ram_1_4 : _GEN_1276; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1533 = unuse_way == 3'h3 ? ram_1_5 : _GEN_1277; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1534 = unuse_way == 3'h3 ? ram_1_6 : _GEN_1278; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1535 = unuse_way == 3'h3 ? ram_1_7 : _GEN_1279; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1536 = unuse_way == 3'h3 ? ram_1_8 : _GEN_1280; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1537 = unuse_way == 3'h3 ? ram_1_9 : _GEN_1281; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1538 = unuse_way == 3'h3 ? ram_1_10 : _GEN_1282; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1539 = unuse_way == 3'h3 ? ram_1_11 : _GEN_1283; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1540 = unuse_way == 3'h3 ? ram_1_12 : _GEN_1284; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1541 = unuse_way == 3'h3 ? ram_1_13 : _GEN_1285; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1542 = unuse_way == 3'h3 ? ram_1_14 : _GEN_1286; // @[i_cache.scala 20:24 95:40]
  wire [511:0] _GEN_1543 = unuse_way == 3'h3 ? ram_1_15 : _GEN_1287; // @[i_cache.scala 20:24 95:40]
  wire [31:0] _GEN_1544 = unuse_way == 3'h3 ? tag_1_0 : _GEN_1288; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1545 = unuse_way == 3'h3 ? tag_1_1 : _GEN_1289; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1546 = unuse_way == 3'h3 ? tag_1_2 : _GEN_1290; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1547 = unuse_way == 3'h3 ? tag_1_3 : _GEN_1291; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1548 = unuse_way == 3'h3 ? tag_1_4 : _GEN_1292; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1549 = unuse_way == 3'h3 ? tag_1_5 : _GEN_1293; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1550 = unuse_way == 3'h3 ? tag_1_6 : _GEN_1294; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1551 = unuse_way == 3'h3 ? tag_1_7 : _GEN_1295; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1552 = unuse_way == 3'h3 ? tag_1_8 : _GEN_1296; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1553 = unuse_way == 3'h3 ? tag_1_9 : _GEN_1297; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1554 = unuse_way == 3'h3 ? tag_1_10 : _GEN_1298; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1555 = unuse_way == 3'h3 ? tag_1_11 : _GEN_1299; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1556 = unuse_way == 3'h3 ? tag_1_12 : _GEN_1300; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1557 = unuse_way == 3'h3 ? tag_1_13 : _GEN_1301; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1558 = unuse_way == 3'h3 ? tag_1_14 : _GEN_1302; // @[i_cache.scala 24:24 95:40]
  wire [31:0] _GEN_1559 = unuse_way == 3'h3 ? tag_1_15 : _GEN_1303; // @[i_cache.scala 24:24 95:40]
  wire  _GEN_1560 = unuse_way == 3'h3 ? valid_1_0 : _GEN_1304; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1561 = unuse_way == 3'h3 ? valid_1_1 : _GEN_1305; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1562 = unuse_way == 3'h3 ? valid_1_2 : _GEN_1306; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1563 = unuse_way == 3'h3 ? valid_1_3 : _GEN_1307; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1564 = unuse_way == 3'h3 ? valid_1_4 : _GEN_1308; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1565 = unuse_way == 3'h3 ? valid_1_5 : _GEN_1309; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1566 = unuse_way == 3'h3 ? valid_1_6 : _GEN_1310; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1567 = unuse_way == 3'h3 ? valid_1_7 : _GEN_1311; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1568 = unuse_way == 3'h3 ? valid_1_8 : _GEN_1312; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1569 = unuse_way == 3'h3 ? valid_1_9 : _GEN_1313; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1570 = unuse_way == 3'h3 ? valid_1_10 : _GEN_1314; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1571 = unuse_way == 3'h3 ? valid_1_11 : _GEN_1315; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1572 = unuse_way == 3'h3 ? valid_1_12 : _GEN_1316; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1573 = unuse_way == 3'h3 ? valid_1_13 : _GEN_1317; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1574 = unuse_way == 3'h3 ? valid_1_14 : _GEN_1318; // @[i_cache.scala 28:26 95:40]
  wire  _GEN_1575 = unuse_way == 3'h3 ? valid_1_15 : _GEN_1319; // @[i_cache.scala 28:26 95:40]
  wire [511:0] _GEN_1576 = unuse_way == 3'h2 ? _GEN_232 : _GEN_1528; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1577 = unuse_way == 3'h2 ? _GEN_233 : _GEN_1529; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1578 = unuse_way == 3'h2 ? _GEN_234 : _GEN_1530; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1579 = unuse_way == 3'h2 ? _GEN_235 : _GEN_1531; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1580 = unuse_way == 3'h2 ? _GEN_236 : _GEN_1532; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1581 = unuse_way == 3'h2 ? _GEN_237 : _GEN_1533; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1582 = unuse_way == 3'h2 ? _GEN_238 : _GEN_1534; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1583 = unuse_way == 3'h2 ? _GEN_239 : _GEN_1535; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1584 = unuse_way == 3'h2 ? _GEN_240 : _GEN_1536; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1585 = unuse_way == 3'h2 ? _GEN_241 : _GEN_1537; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1586 = unuse_way == 3'h2 ? _GEN_242 : _GEN_1538; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1587 = unuse_way == 3'h2 ? _GEN_243 : _GEN_1539; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1588 = unuse_way == 3'h2 ? _GEN_244 : _GEN_1540; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1589 = unuse_way == 3'h2 ? _GEN_245 : _GEN_1541; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1590 = unuse_way == 3'h2 ? _GEN_246 : _GEN_1542; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1591 = unuse_way == 3'h2 ? _GEN_247 : _GEN_1543; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1592 = unuse_way == 3'h2 ? _GEN_248 : _GEN_1544; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1593 = unuse_way == 3'h2 ? _GEN_249 : _GEN_1545; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1594 = unuse_way == 3'h2 ? _GEN_250 : _GEN_1546; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1595 = unuse_way == 3'h2 ? _GEN_251 : _GEN_1547; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1596 = unuse_way == 3'h2 ? _GEN_252 : _GEN_1548; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1597 = unuse_way == 3'h2 ? _GEN_253 : _GEN_1549; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1598 = unuse_way == 3'h2 ? _GEN_254 : _GEN_1550; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1599 = unuse_way == 3'h2 ? _GEN_255 : _GEN_1551; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1600 = unuse_way == 3'h2 ? _GEN_256 : _GEN_1552; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1601 = unuse_way == 3'h2 ? _GEN_257 : _GEN_1553; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1602 = unuse_way == 3'h2 ? _GEN_258 : _GEN_1554; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1603 = unuse_way == 3'h2 ? _GEN_259 : _GEN_1555; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1604 = unuse_way == 3'h2 ? _GEN_260 : _GEN_1556; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1605 = unuse_way == 3'h2 ? _GEN_261 : _GEN_1557; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1606 = unuse_way == 3'h2 ? _GEN_262 : _GEN_1558; // @[i_cache.scala 90:40]
  wire [31:0] _GEN_1607 = unuse_way == 3'h2 ? _GEN_263 : _GEN_1559; // @[i_cache.scala 90:40]
  wire  _GEN_1608 = unuse_way == 3'h2 ? _GEN_264 : _GEN_1560; // @[i_cache.scala 90:40]
  wire  _GEN_1609 = unuse_way == 3'h2 ? _GEN_265 : _GEN_1561; // @[i_cache.scala 90:40]
  wire  _GEN_1610 = unuse_way == 3'h2 ? _GEN_266 : _GEN_1562; // @[i_cache.scala 90:40]
  wire  _GEN_1611 = unuse_way == 3'h2 ? _GEN_267 : _GEN_1563; // @[i_cache.scala 90:40]
  wire  _GEN_1612 = unuse_way == 3'h2 ? _GEN_268 : _GEN_1564; // @[i_cache.scala 90:40]
  wire  _GEN_1613 = unuse_way == 3'h2 ? _GEN_269 : _GEN_1565; // @[i_cache.scala 90:40]
  wire  _GEN_1614 = unuse_way == 3'h2 ? _GEN_270 : _GEN_1566; // @[i_cache.scala 90:40]
  wire  _GEN_1615 = unuse_way == 3'h2 ? _GEN_271 : _GEN_1567; // @[i_cache.scala 90:40]
  wire  _GEN_1616 = unuse_way == 3'h2 ? _GEN_272 : _GEN_1568; // @[i_cache.scala 90:40]
  wire  _GEN_1617 = unuse_way == 3'h2 ? _GEN_273 : _GEN_1569; // @[i_cache.scala 90:40]
  wire  _GEN_1618 = unuse_way == 3'h2 ? _GEN_274 : _GEN_1570; // @[i_cache.scala 90:40]
  wire  _GEN_1619 = unuse_way == 3'h2 ? _GEN_275 : _GEN_1571; // @[i_cache.scala 90:40]
  wire  _GEN_1620 = unuse_way == 3'h2 ? _GEN_276 : _GEN_1572; // @[i_cache.scala 90:40]
  wire  _GEN_1621 = unuse_way == 3'h2 ? _GEN_277 : _GEN_1573; // @[i_cache.scala 90:40]
  wire  _GEN_1622 = unuse_way == 3'h2 ? _GEN_278 : _GEN_1574; // @[i_cache.scala 90:40]
  wire  _GEN_1623 = unuse_way == 3'h2 ? _GEN_279 : _GEN_1575; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1624 = unuse_way == 3'h2 ? _GEN_280 : _GEN_1416; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1625 = unuse_way == 3'h2 ? _GEN_281 : _GEN_1417; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1626 = unuse_way == 3'h2 ? _GEN_282 : _GEN_1418; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1627 = unuse_way == 3'h2 ? _GEN_283 : _GEN_1419; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1628 = unuse_way == 3'h2 ? _GEN_284 : _GEN_1420; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1629 = unuse_way == 3'h2 ? _GEN_285 : _GEN_1421; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1630 = unuse_way == 3'h2 ? _GEN_286 : _GEN_1422; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1631 = unuse_way == 3'h2 ? _GEN_287 : _GEN_1423; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1632 = unuse_way == 3'h2 ? _GEN_288 : _GEN_1424; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1633 = unuse_way == 3'h2 ? _GEN_289 : _GEN_1425; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1634 = unuse_way == 3'h2 ? _GEN_290 : _GEN_1426; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1635 = unuse_way == 3'h2 ? _GEN_291 : _GEN_1427; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1636 = unuse_way == 3'h2 ? _GEN_292 : _GEN_1428; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1637 = unuse_way == 3'h2 ? _GEN_293 : _GEN_1429; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1638 = unuse_way == 3'h2 ? _GEN_294 : _GEN_1430; // @[i_cache.scala 90:40]
  wire [7:0] _GEN_1639 = unuse_way == 3'h2 ? _GEN_295 : _GEN_1431; // @[i_cache.scala 90:40]
  wire [511:0] _GEN_1640 = unuse_way == 3'h2 ? ram_2_0 : _GEN_1368; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1641 = unuse_way == 3'h2 ? ram_2_1 : _GEN_1369; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1642 = unuse_way == 3'h2 ? ram_2_2 : _GEN_1370; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1643 = unuse_way == 3'h2 ? ram_2_3 : _GEN_1371; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1644 = unuse_way == 3'h2 ? ram_2_4 : _GEN_1372; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1645 = unuse_way == 3'h2 ? ram_2_5 : _GEN_1373; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1646 = unuse_way == 3'h2 ? ram_2_6 : _GEN_1374; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1647 = unuse_way == 3'h2 ? ram_2_7 : _GEN_1375; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1648 = unuse_way == 3'h2 ? ram_2_8 : _GEN_1376; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1649 = unuse_way == 3'h2 ? ram_2_9 : _GEN_1377; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1650 = unuse_way == 3'h2 ? ram_2_10 : _GEN_1378; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1651 = unuse_way == 3'h2 ? ram_2_11 : _GEN_1379; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1652 = unuse_way == 3'h2 ? ram_2_12 : _GEN_1380; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1653 = unuse_way == 3'h2 ? ram_2_13 : _GEN_1381; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1654 = unuse_way == 3'h2 ? ram_2_14 : _GEN_1382; // @[i_cache.scala 21:24 90:40]
  wire [511:0] _GEN_1655 = unuse_way == 3'h2 ? ram_2_15 : _GEN_1383; // @[i_cache.scala 21:24 90:40]
  wire [31:0] _GEN_1656 = unuse_way == 3'h2 ? tag_2_0 : _GEN_1384; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1657 = unuse_way == 3'h2 ? tag_2_1 : _GEN_1385; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1658 = unuse_way == 3'h2 ? tag_2_2 : _GEN_1386; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1659 = unuse_way == 3'h2 ? tag_2_3 : _GEN_1387; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1660 = unuse_way == 3'h2 ? tag_2_4 : _GEN_1388; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1661 = unuse_way == 3'h2 ? tag_2_5 : _GEN_1389; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1662 = unuse_way == 3'h2 ? tag_2_6 : _GEN_1390; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1663 = unuse_way == 3'h2 ? tag_2_7 : _GEN_1391; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1664 = unuse_way == 3'h2 ? tag_2_8 : _GEN_1392; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1665 = unuse_way == 3'h2 ? tag_2_9 : _GEN_1393; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1666 = unuse_way == 3'h2 ? tag_2_10 : _GEN_1394; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1667 = unuse_way == 3'h2 ? tag_2_11 : _GEN_1395; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1668 = unuse_way == 3'h2 ? tag_2_12 : _GEN_1396; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1669 = unuse_way == 3'h2 ? tag_2_13 : _GEN_1397; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1670 = unuse_way == 3'h2 ? tag_2_14 : _GEN_1398; // @[i_cache.scala 25:24 90:40]
  wire [31:0] _GEN_1671 = unuse_way == 3'h2 ? tag_2_15 : _GEN_1399; // @[i_cache.scala 25:24 90:40]
  wire  _GEN_1672 = unuse_way == 3'h2 ? valid_2_0 : _GEN_1400; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1673 = unuse_way == 3'h2 ? valid_2_1 : _GEN_1401; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1674 = unuse_way == 3'h2 ? valid_2_2 : _GEN_1402; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1675 = unuse_way == 3'h2 ? valid_2_3 : _GEN_1403; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1676 = unuse_way == 3'h2 ? valid_2_4 : _GEN_1404; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1677 = unuse_way == 3'h2 ? valid_2_5 : _GEN_1405; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1678 = unuse_way == 3'h2 ? valid_2_6 : _GEN_1406; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1679 = unuse_way == 3'h2 ? valid_2_7 : _GEN_1407; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1680 = unuse_way == 3'h2 ? valid_2_8 : _GEN_1408; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1681 = unuse_way == 3'h2 ? valid_2_9 : _GEN_1409; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1682 = unuse_way == 3'h2 ? valid_2_10 : _GEN_1410; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1683 = unuse_way == 3'h2 ? valid_2_11 : _GEN_1411; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1684 = unuse_way == 3'h2 ? valid_2_12 : _GEN_1412; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1685 = unuse_way == 3'h2 ? valid_2_13 : _GEN_1413; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1686 = unuse_way == 3'h2 ? valid_2_14 : _GEN_1414; // @[i_cache.scala 29:26 90:40]
  wire  _GEN_1687 = unuse_way == 3'h2 ? valid_2_15 : _GEN_1415; // @[i_cache.scala 29:26 90:40]
  wire [511:0] _GEN_1688 = unuse_way == 3'h2 ? ram_3_0 : _GEN_1432; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1689 = unuse_way == 3'h2 ? ram_3_1 : _GEN_1433; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1690 = unuse_way == 3'h2 ? ram_3_2 : _GEN_1434; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1691 = unuse_way == 3'h2 ? ram_3_3 : _GEN_1435; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1692 = unuse_way == 3'h2 ? ram_3_4 : _GEN_1436; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1693 = unuse_way == 3'h2 ? ram_3_5 : _GEN_1437; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1694 = unuse_way == 3'h2 ? ram_3_6 : _GEN_1438; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1695 = unuse_way == 3'h2 ? ram_3_7 : _GEN_1439; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1696 = unuse_way == 3'h2 ? ram_3_8 : _GEN_1440; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1697 = unuse_way == 3'h2 ? ram_3_9 : _GEN_1441; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1698 = unuse_way == 3'h2 ? ram_3_10 : _GEN_1442; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1699 = unuse_way == 3'h2 ? ram_3_11 : _GEN_1443; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1700 = unuse_way == 3'h2 ? ram_3_12 : _GEN_1444; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1701 = unuse_way == 3'h2 ? ram_3_13 : _GEN_1445; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1702 = unuse_way == 3'h2 ? ram_3_14 : _GEN_1446; // @[i_cache.scala 22:24 90:40]
  wire [511:0] _GEN_1703 = unuse_way == 3'h2 ? ram_3_15 : _GEN_1447; // @[i_cache.scala 22:24 90:40]
  wire [31:0] _GEN_1704 = unuse_way == 3'h2 ? tag_3_0 : _GEN_1448; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1705 = unuse_way == 3'h2 ? tag_3_1 : _GEN_1449; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1706 = unuse_way == 3'h2 ? tag_3_2 : _GEN_1450; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1707 = unuse_way == 3'h2 ? tag_3_3 : _GEN_1451; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1708 = unuse_way == 3'h2 ? tag_3_4 : _GEN_1452; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1709 = unuse_way == 3'h2 ? tag_3_5 : _GEN_1453; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1710 = unuse_way == 3'h2 ? tag_3_6 : _GEN_1454; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1711 = unuse_way == 3'h2 ? tag_3_7 : _GEN_1455; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1712 = unuse_way == 3'h2 ? tag_3_8 : _GEN_1456; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1713 = unuse_way == 3'h2 ? tag_3_9 : _GEN_1457; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1714 = unuse_way == 3'h2 ? tag_3_10 : _GEN_1458; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1715 = unuse_way == 3'h2 ? tag_3_11 : _GEN_1459; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1716 = unuse_way == 3'h2 ? tag_3_12 : _GEN_1460; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1717 = unuse_way == 3'h2 ? tag_3_13 : _GEN_1461; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1718 = unuse_way == 3'h2 ? tag_3_14 : _GEN_1462; // @[i_cache.scala 26:24 90:40]
  wire [31:0] _GEN_1719 = unuse_way == 3'h2 ? tag_3_15 : _GEN_1463; // @[i_cache.scala 26:24 90:40]
  wire  _GEN_1720 = unuse_way == 3'h2 ? valid_3_0 : _GEN_1464; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1721 = unuse_way == 3'h2 ? valid_3_1 : _GEN_1465; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1722 = unuse_way == 3'h2 ? valid_3_2 : _GEN_1466; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1723 = unuse_way == 3'h2 ? valid_3_3 : _GEN_1467; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1724 = unuse_way == 3'h2 ? valid_3_4 : _GEN_1468; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1725 = unuse_way == 3'h2 ? valid_3_5 : _GEN_1469; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1726 = unuse_way == 3'h2 ? valid_3_6 : _GEN_1470; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1727 = unuse_way == 3'h2 ? valid_3_7 : _GEN_1471; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1728 = unuse_way == 3'h2 ? valid_3_8 : _GEN_1472; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1729 = unuse_way == 3'h2 ? valid_3_9 : _GEN_1473; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1730 = unuse_way == 3'h2 ? valid_3_10 : _GEN_1474; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1731 = unuse_way == 3'h2 ? valid_3_11 : _GEN_1475; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1732 = unuse_way == 3'h2 ? valid_3_12 : _GEN_1476; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1733 = unuse_way == 3'h2 ? valid_3_13 : _GEN_1477; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1734 = unuse_way == 3'h2 ? valid_3_14 : _GEN_1478; // @[i_cache.scala 30:26 90:40]
  wire  _GEN_1735 = unuse_way == 3'h2 ? valid_3_15 : _GEN_1479; // @[i_cache.scala 30:26 90:40]
  wire [511:0] _GEN_1736 = unuse_way == 3'h2 ? ram_0_0 : _GEN_1480; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1737 = unuse_way == 3'h2 ? ram_0_1 : _GEN_1481; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1738 = unuse_way == 3'h2 ? ram_0_2 : _GEN_1482; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1739 = unuse_way == 3'h2 ? ram_0_3 : _GEN_1483; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1740 = unuse_way == 3'h2 ? ram_0_4 : _GEN_1484; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1741 = unuse_way == 3'h2 ? ram_0_5 : _GEN_1485; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1742 = unuse_way == 3'h2 ? ram_0_6 : _GEN_1486; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1743 = unuse_way == 3'h2 ? ram_0_7 : _GEN_1487; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1744 = unuse_way == 3'h2 ? ram_0_8 : _GEN_1488; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1745 = unuse_way == 3'h2 ? ram_0_9 : _GEN_1489; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1746 = unuse_way == 3'h2 ? ram_0_10 : _GEN_1490; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1747 = unuse_way == 3'h2 ? ram_0_11 : _GEN_1491; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1748 = unuse_way == 3'h2 ? ram_0_12 : _GEN_1492; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1749 = unuse_way == 3'h2 ? ram_0_13 : _GEN_1493; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1750 = unuse_way == 3'h2 ? ram_0_14 : _GEN_1494; // @[i_cache.scala 19:24 90:40]
  wire [511:0] _GEN_1751 = unuse_way == 3'h2 ? ram_0_15 : _GEN_1495; // @[i_cache.scala 19:24 90:40]
  wire [31:0] _GEN_1752 = unuse_way == 3'h2 ? tag_0_0 : _GEN_1496; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1753 = unuse_way == 3'h2 ? tag_0_1 : _GEN_1497; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1754 = unuse_way == 3'h2 ? tag_0_2 : _GEN_1498; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1755 = unuse_way == 3'h2 ? tag_0_3 : _GEN_1499; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1756 = unuse_way == 3'h2 ? tag_0_4 : _GEN_1500; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1757 = unuse_way == 3'h2 ? tag_0_5 : _GEN_1501; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1758 = unuse_way == 3'h2 ? tag_0_6 : _GEN_1502; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1759 = unuse_way == 3'h2 ? tag_0_7 : _GEN_1503; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1760 = unuse_way == 3'h2 ? tag_0_8 : _GEN_1504; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1761 = unuse_way == 3'h2 ? tag_0_9 : _GEN_1505; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1762 = unuse_way == 3'h2 ? tag_0_10 : _GEN_1506; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1763 = unuse_way == 3'h2 ? tag_0_11 : _GEN_1507; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1764 = unuse_way == 3'h2 ? tag_0_12 : _GEN_1508; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1765 = unuse_way == 3'h2 ? tag_0_13 : _GEN_1509; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1766 = unuse_way == 3'h2 ? tag_0_14 : _GEN_1510; // @[i_cache.scala 23:24 90:40]
  wire [31:0] _GEN_1767 = unuse_way == 3'h2 ? tag_0_15 : _GEN_1511; // @[i_cache.scala 23:24 90:40]
  wire  _GEN_1768 = unuse_way == 3'h2 ? valid_0_0 : _GEN_1512; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1769 = unuse_way == 3'h2 ? valid_0_1 : _GEN_1513; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1770 = unuse_way == 3'h2 ? valid_0_2 : _GEN_1514; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1771 = unuse_way == 3'h2 ? valid_0_3 : _GEN_1515; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1772 = unuse_way == 3'h2 ? valid_0_4 : _GEN_1516; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1773 = unuse_way == 3'h2 ? valid_0_5 : _GEN_1517; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1774 = unuse_way == 3'h2 ? valid_0_6 : _GEN_1518; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1775 = unuse_way == 3'h2 ? valid_0_7 : _GEN_1519; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1776 = unuse_way == 3'h2 ? valid_0_8 : _GEN_1520; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1777 = unuse_way == 3'h2 ? valid_0_9 : _GEN_1521; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1778 = unuse_way == 3'h2 ? valid_0_10 : _GEN_1522; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1779 = unuse_way == 3'h2 ? valid_0_11 : _GEN_1523; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1780 = unuse_way == 3'h2 ? valid_0_12 : _GEN_1524; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1781 = unuse_way == 3'h2 ? valid_0_13 : _GEN_1525; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1782 = unuse_way == 3'h2 ? valid_0_14 : _GEN_1526; // @[i_cache.scala 27:26 90:40]
  wire  _GEN_1783 = unuse_way == 3'h2 ? valid_0_15 : _GEN_1527; // @[i_cache.scala 27:26 90:40]
  wire [511:0] _GEN_1784 = unuse_way == 3'h1 ? _GEN_152 : _GEN_1736; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1785 = unuse_way == 3'h1 ? _GEN_153 : _GEN_1737; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1786 = unuse_way == 3'h1 ? _GEN_154 : _GEN_1738; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1787 = unuse_way == 3'h1 ? _GEN_155 : _GEN_1739; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1788 = unuse_way == 3'h1 ? _GEN_156 : _GEN_1740; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1789 = unuse_way == 3'h1 ? _GEN_157 : _GEN_1741; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1790 = unuse_way == 3'h1 ? _GEN_158 : _GEN_1742; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1791 = unuse_way == 3'h1 ? _GEN_159 : _GEN_1743; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1792 = unuse_way == 3'h1 ? _GEN_160 : _GEN_1744; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1793 = unuse_way == 3'h1 ? _GEN_161 : _GEN_1745; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1794 = unuse_way == 3'h1 ? _GEN_162 : _GEN_1746; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1795 = unuse_way == 3'h1 ? _GEN_163 : _GEN_1747; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1796 = unuse_way == 3'h1 ? _GEN_164 : _GEN_1748; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1797 = unuse_way == 3'h1 ? _GEN_165 : _GEN_1749; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1798 = unuse_way == 3'h1 ? _GEN_166 : _GEN_1750; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1799 = unuse_way == 3'h1 ? _GEN_167 : _GEN_1751; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1800 = unuse_way == 3'h1 ? _GEN_168 : _GEN_1752; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1801 = unuse_way == 3'h1 ? _GEN_169 : _GEN_1753; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1802 = unuse_way == 3'h1 ? _GEN_170 : _GEN_1754; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1803 = unuse_way == 3'h1 ? _GEN_171 : _GEN_1755; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1804 = unuse_way == 3'h1 ? _GEN_172 : _GEN_1756; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1805 = unuse_way == 3'h1 ? _GEN_173 : _GEN_1757; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1806 = unuse_way == 3'h1 ? _GEN_174 : _GEN_1758; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1807 = unuse_way == 3'h1 ? _GEN_175 : _GEN_1759; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1808 = unuse_way == 3'h1 ? _GEN_176 : _GEN_1760; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1809 = unuse_way == 3'h1 ? _GEN_177 : _GEN_1761; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1810 = unuse_way == 3'h1 ? _GEN_178 : _GEN_1762; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1811 = unuse_way == 3'h1 ? _GEN_179 : _GEN_1763; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1812 = unuse_way == 3'h1 ? _GEN_180 : _GEN_1764; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1813 = unuse_way == 3'h1 ? _GEN_181 : _GEN_1765; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1814 = unuse_way == 3'h1 ? _GEN_182 : _GEN_1766; // @[i_cache.scala 85:34]
  wire [31:0] _GEN_1815 = unuse_way == 3'h1 ? _GEN_183 : _GEN_1767; // @[i_cache.scala 85:34]
  wire  _GEN_1816 = unuse_way == 3'h1 ? _GEN_184 : _GEN_1768; // @[i_cache.scala 85:34]
  wire  _GEN_1817 = unuse_way == 3'h1 ? _GEN_185 : _GEN_1769; // @[i_cache.scala 85:34]
  wire  _GEN_1818 = unuse_way == 3'h1 ? _GEN_186 : _GEN_1770; // @[i_cache.scala 85:34]
  wire  _GEN_1819 = unuse_way == 3'h1 ? _GEN_187 : _GEN_1771; // @[i_cache.scala 85:34]
  wire  _GEN_1820 = unuse_way == 3'h1 ? _GEN_188 : _GEN_1772; // @[i_cache.scala 85:34]
  wire  _GEN_1821 = unuse_way == 3'h1 ? _GEN_189 : _GEN_1773; // @[i_cache.scala 85:34]
  wire  _GEN_1822 = unuse_way == 3'h1 ? _GEN_190 : _GEN_1774; // @[i_cache.scala 85:34]
  wire  _GEN_1823 = unuse_way == 3'h1 ? _GEN_191 : _GEN_1775; // @[i_cache.scala 85:34]
  wire  _GEN_1824 = unuse_way == 3'h1 ? _GEN_192 : _GEN_1776; // @[i_cache.scala 85:34]
  wire  _GEN_1825 = unuse_way == 3'h1 ? _GEN_193 : _GEN_1777; // @[i_cache.scala 85:34]
  wire  _GEN_1826 = unuse_way == 3'h1 ? _GEN_194 : _GEN_1778; // @[i_cache.scala 85:34]
  wire  _GEN_1827 = unuse_way == 3'h1 ? _GEN_195 : _GEN_1779; // @[i_cache.scala 85:34]
  wire  _GEN_1828 = unuse_way == 3'h1 ? _GEN_196 : _GEN_1780; // @[i_cache.scala 85:34]
  wire  _GEN_1829 = unuse_way == 3'h1 ? _GEN_197 : _GEN_1781; // @[i_cache.scala 85:34]
  wire  _GEN_1830 = unuse_way == 3'h1 ? _GEN_198 : _GEN_1782; // @[i_cache.scala 85:34]
  wire  _GEN_1831 = unuse_way == 3'h1 ? _GEN_199 : _GEN_1783; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1832 = unuse_way == 3'h1 ? _GEN_216 : _GEN_1624; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1833 = unuse_way == 3'h1 ? _GEN_217 : _GEN_1625; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1834 = unuse_way == 3'h1 ? _GEN_218 : _GEN_1626; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1835 = unuse_way == 3'h1 ? _GEN_219 : _GEN_1627; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1836 = unuse_way == 3'h1 ? _GEN_220 : _GEN_1628; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1837 = unuse_way == 3'h1 ? _GEN_221 : _GEN_1629; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1838 = unuse_way == 3'h1 ? _GEN_222 : _GEN_1630; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1839 = unuse_way == 3'h1 ? _GEN_223 : _GEN_1631; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1840 = unuse_way == 3'h1 ? _GEN_224 : _GEN_1632; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1841 = unuse_way == 3'h1 ? _GEN_225 : _GEN_1633; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1842 = unuse_way == 3'h1 ? _GEN_226 : _GEN_1634; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1843 = unuse_way == 3'h1 ? _GEN_227 : _GEN_1635; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1844 = unuse_way == 3'h1 ? _GEN_228 : _GEN_1636; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1845 = unuse_way == 3'h1 ? _GEN_229 : _GEN_1637; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1846 = unuse_way == 3'h1 ? _GEN_230 : _GEN_1638; // @[i_cache.scala 85:34]
  wire [7:0] _GEN_1847 = unuse_way == 3'h1 ? _GEN_231 : _GEN_1639; // @[i_cache.scala 85:34]
  wire [511:0] _GEN_1848 = unuse_way == 3'h1 ? ram_1_0 : _GEN_1576; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1849 = unuse_way == 3'h1 ? ram_1_1 : _GEN_1577; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1850 = unuse_way == 3'h1 ? ram_1_2 : _GEN_1578; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1851 = unuse_way == 3'h1 ? ram_1_3 : _GEN_1579; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1852 = unuse_way == 3'h1 ? ram_1_4 : _GEN_1580; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1853 = unuse_way == 3'h1 ? ram_1_5 : _GEN_1581; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1854 = unuse_way == 3'h1 ? ram_1_6 : _GEN_1582; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1855 = unuse_way == 3'h1 ? ram_1_7 : _GEN_1583; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1856 = unuse_way == 3'h1 ? ram_1_8 : _GEN_1584; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1857 = unuse_way == 3'h1 ? ram_1_9 : _GEN_1585; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1858 = unuse_way == 3'h1 ? ram_1_10 : _GEN_1586; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1859 = unuse_way == 3'h1 ? ram_1_11 : _GEN_1587; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1860 = unuse_way == 3'h1 ? ram_1_12 : _GEN_1588; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1861 = unuse_way == 3'h1 ? ram_1_13 : _GEN_1589; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1862 = unuse_way == 3'h1 ? ram_1_14 : _GEN_1590; // @[i_cache.scala 20:24 85:34]
  wire [511:0] _GEN_1863 = unuse_way == 3'h1 ? ram_1_15 : _GEN_1591; // @[i_cache.scala 20:24 85:34]
  wire [31:0] _GEN_1864 = unuse_way == 3'h1 ? tag_1_0 : _GEN_1592; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1865 = unuse_way == 3'h1 ? tag_1_1 : _GEN_1593; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1866 = unuse_way == 3'h1 ? tag_1_2 : _GEN_1594; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1867 = unuse_way == 3'h1 ? tag_1_3 : _GEN_1595; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1868 = unuse_way == 3'h1 ? tag_1_4 : _GEN_1596; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1869 = unuse_way == 3'h1 ? tag_1_5 : _GEN_1597; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1870 = unuse_way == 3'h1 ? tag_1_6 : _GEN_1598; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1871 = unuse_way == 3'h1 ? tag_1_7 : _GEN_1599; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1872 = unuse_way == 3'h1 ? tag_1_8 : _GEN_1600; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1873 = unuse_way == 3'h1 ? tag_1_9 : _GEN_1601; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1874 = unuse_way == 3'h1 ? tag_1_10 : _GEN_1602; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1875 = unuse_way == 3'h1 ? tag_1_11 : _GEN_1603; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1876 = unuse_way == 3'h1 ? tag_1_12 : _GEN_1604; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1877 = unuse_way == 3'h1 ? tag_1_13 : _GEN_1605; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1878 = unuse_way == 3'h1 ? tag_1_14 : _GEN_1606; // @[i_cache.scala 24:24 85:34]
  wire [31:0] _GEN_1879 = unuse_way == 3'h1 ? tag_1_15 : _GEN_1607; // @[i_cache.scala 24:24 85:34]
  wire  _GEN_1880 = unuse_way == 3'h1 ? valid_1_0 : _GEN_1608; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1881 = unuse_way == 3'h1 ? valid_1_1 : _GEN_1609; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1882 = unuse_way == 3'h1 ? valid_1_2 : _GEN_1610; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1883 = unuse_way == 3'h1 ? valid_1_3 : _GEN_1611; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1884 = unuse_way == 3'h1 ? valid_1_4 : _GEN_1612; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1885 = unuse_way == 3'h1 ? valid_1_5 : _GEN_1613; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1886 = unuse_way == 3'h1 ? valid_1_6 : _GEN_1614; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1887 = unuse_way == 3'h1 ? valid_1_7 : _GEN_1615; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1888 = unuse_way == 3'h1 ? valid_1_8 : _GEN_1616; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1889 = unuse_way == 3'h1 ? valid_1_9 : _GEN_1617; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1890 = unuse_way == 3'h1 ? valid_1_10 : _GEN_1618; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1891 = unuse_way == 3'h1 ? valid_1_11 : _GEN_1619; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1892 = unuse_way == 3'h1 ? valid_1_12 : _GEN_1620; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1893 = unuse_way == 3'h1 ? valid_1_13 : _GEN_1621; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1894 = unuse_way == 3'h1 ? valid_1_14 : _GEN_1622; // @[i_cache.scala 28:26 85:34]
  wire  _GEN_1895 = unuse_way == 3'h1 ? valid_1_15 : _GEN_1623; // @[i_cache.scala 28:26 85:34]
  wire [511:0] _GEN_1896 = unuse_way == 3'h1 ? ram_2_0 : _GEN_1640; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1897 = unuse_way == 3'h1 ? ram_2_1 : _GEN_1641; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1898 = unuse_way == 3'h1 ? ram_2_2 : _GEN_1642; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1899 = unuse_way == 3'h1 ? ram_2_3 : _GEN_1643; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1900 = unuse_way == 3'h1 ? ram_2_4 : _GEN_1644; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1901 = unuse_way == 3'h1 ? ram_2_5 : _GEN_1645; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1902 = unuse_way == 3'h1 ? ram_2_6 : _GEN_1646; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1903 = unuse_way == 3'h1 ? ram_2_7 : _GEN_1647; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1904 = unuse_way == 3'h1 ? ram_2_8 : _GEN_1648; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1905 = unuse_way == 3'h1 ? ram_2_9 : _GEN_1649; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1906 = unuse_way == 3'h1 ? ram_2_10 : _GEN_1650; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1907 = unuse_way == 3'h1 ? ram_2_11 : _GEN_1651; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1908 = unuse_way == 3'h1 ? ram_2_12 : _GEN_1652; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1909 = unuse_way == 3'h1 ? ram_2_13 : _GEN_1653; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1910 = unuse_way == 3'h1 ? ram_2_14 : _GEN_1654; // @[i_cache.scala 21:24 85:34]
  wire [511:0] _GEN_1911 = unuse_way == 3'h1 ? ram_2_15 : _GEN_1655; // @[i_cache.scala 21:24 85:34]
  wire [31:0] _GEN_1912 = unuse_way == 3'h1 ? tag_2_0 : _GEN_1656; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1913 = unuse_way == 3'h1 ? tag_2_1 : _GEN_1657; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1914 = unuse_way == 3'h1 ? tag_2_2 : _GEN_1658; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1915 = unuse_way == 3'h1 ? tag_2_3 : _GEN_1659; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1916 = unuse_way == 3'h1 ? tag_2_4 : _GEN_1660; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1917 = unuse_way == 3'h1 ? tag_2_5 : _GEN_1661; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1918 = unuse_way == 3'h1 ? tag_2_6 : _GEN_1662; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1919 = unuse_way == 3'h1 ? tag_2_7 : _GEN_1663; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1920 = unuse_way == 3'h1 ? tag_2_8 : _GEN_1664; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1921 = unuse_way == 3'h1 ? tag_2_9 : _GEN_1665; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1922 = unuse_way == 3'h1 ? tag_2_10 : _GEN_1666; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1923 = unuse_way == 3'h1 ? tag_2_11 : _GEN_1667; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1924 = unuse_way == 3'h1 ? tag_2_12 : _GEN_1668; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1925 = unuse_way == 3'h1 ? tag_2_13 : _GEN_1669; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1926 = unuse_way == 3'h1 ? tag_2_14 : _GEN_1670; // @[i_cache.scala 25:24 85:34]
  wire [31:0] _GEN_1927 = unuse_way == 3'h1 ? tag_2_15 : _GEN_1671; // @[i_cache.scala 25:24 85:34]
  wire  _GEN_1928 = unuse_way == 3'h1 ? valid_2_0 : _GEN_1672; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1929 = unuse_way == 3'h1 ? valid_2_1 : _GEN_1673; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1930 = unuse_way == 3'h1 ? valid_2_2 : _GEN_1674; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1931 = unuse_way == 3'h1 ? valid_2_3 : _GEN_1675; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1932 = unuse_way == 3'h1 ? valid_2_4 : _GEN_1676; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1933 = unuse_way == 3'h1 ? valid_2_5 : _GEN_1677; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1934 = unuse_way == 3'h1 ? valid_2_6 : _GEN_1678; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1935 = unuse_way == 3'h1 ? valid_2_7 : _GEN_1679; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1936 = unuse_way == 3'h1 ? valid_2_8 : _GEN_1680; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1937 = unuse_way == 3'h1 ? valid_2_9 : _GEN_1681; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1938 = unuse_way == 3'h1 ? valid_2_10 : _GEN_1682; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1939 = unuse_way == 3'h1 ? valid_2_11 : _GEN_1683; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1940 = unuse_way == 3'h1 ? valid_2_12 : _GEN_1684; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1941 = unuse_way == 3'h1 ? valid_2_13 : _GEN_1685; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1942 = unuse_way == 3'h1 ? valid_2_14 : _GEN_1686; // @[i_cache.scala 29:26 85:34]
  wire  _GEN_1943 = unuse_way == 3'h1 ? valid_2_15 : _GEN_1687; // @[i_cache.scala 29:26 85:34]
  wire [511:0] _GEN_1944 = unuse_way == 3'h1 ? ram_3_0 : _GEN_1688; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1945 = unuse_way == 3'h1 ? ram_3_1 : _GEN_1689; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1946 = unuse_way == 3'h1 ? ram_3_2 : _GEN_1690; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1947 = unuse_way == 3'h1 ? ram_3_3 : _GEN_1691; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1948 = unuse_way == 3'h1 ? ram_3_4 : _GEN_1692; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1949 = unuse_way == 3'h1 ? ram_3_5 : _GEN_1693; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1950 = unuse_way == 3'h1 ? ram_3_6 : _GEN_1694; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1951 = unuse_way == 3'h1 ? ram_3_7 : _GEN_1695; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1952 = unuse_way == 3'h1 ? ram_3_8 : _GEN_1696; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1953 = unuse_way == 3'h1 ? ram_3_9 : _GEN_1697; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1954 = unuse_way == 3'h1 ? ram_3_10 : _GEN_1698; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1955 = unuse_way == 3'h1 ? ram_3_11 : _GEN_1699; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1956 = unuse_way == 3'h1 ? ram_3_12 : _GEN_1700; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1957 = unuse_way == 3'h1 ? ram_3_13 : _GEN_1701; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1958 = unuse_way == 3'h1 ? ram_3_14 : _GEN_1702; // @[i_cache.scala 22:24 85:34]
  wire [511:0] _GEN_1959 = unuse_way == 3'h1 ? ram_3_15 : _GEN_1703; // @[i_cache.scala 22:24 85:34]
  wire [31:0] _GEN_1960 = unuse_way == 3'h1 ? tag_3_0 : _GEN_1704; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1961 = unuse_way == 3'h1 ? tag_3_1 : _GEN_1705; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1962 = unuse_way == 3'h1 ? tag_3_2 : _GEN_1706; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1963 = unuse_way == 3'h1 ? tag_3_3 : _GEN_1707; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1964 = unuse_way == 3'h1 ? tag_3_4 : _GEN_1708; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1965 = unuse_way == 3'h1 ? tag_3_5 : _GEN_1709; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1966 = unuse_way == 3'h1 ? tag_3_6 : _GEN_1710; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1967 = unuse_way == 3'h1 ? tag_3_7 : _GEN_1711; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1968 = unuse_way == 3'h1 ? tag_3_8 : _GEN_1712; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1969 = unuse_way == 3'h1 ? tag_3_9 : _GEN_1713; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1970 = unuse_way == 3'h1 ? tag_3_10 : _GEN_1714; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1971 = unuse_way == 3'h1 ? tag_3_11 : _GEN_1715; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1972 = unuse_way == 3'h1 ? tag_3_12 : _GEN_1716; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1973 = unuse_way == 3'h1 ? tag_3_13 : _GEN_1717; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1974 = unuse_way == 3'h1 ? tag_3_14 : _GEN_1718; // @[i_cache.scala 26:24 85:34]
  wire [31:0] _GEN_1975 = unuse_way == 3'h1 ? tag_3_15 : _GEN_1719; // @[i_cache.scala 26:24 85:34]
  wire  _GEN_1976 = unuse_way == 3'h1 ? valid_3_0 : _GEN_1720; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1977 = unuse_way == 3'h1 ? valid_3_1 : _GEN_1721; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1978 = unuse_way == 3'h1 ? valid_3_2 : _GEN_1722; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1979 = unuse_way == 3'h1 ? valid_3_3 : _GEN_1723; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1980 = unuse_way == 3'h1 ? valid_3_4 : _GEN_1724; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1981 = unuse_way == 3'h1 ? valid_3_5 : _GEN_1725; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1982 = unuse_way == 3'h1 ? valid_3_6 : _GEN_1726; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1983 = unuse_way == 3'h1 ? valid_3_7 : _GEN_1727; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1984 = unuse_way == 3'h1 ? valid_3_8 : _GEN_1728; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1985 = unuse_way == 3'h1 ? valid_3_9 : _GEN_1729; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1986 = unuse_way == 3'h1 ? valid_3_10 : _GEN_1730; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1987 = unuse_way == 3'h1 ? valid_3_11 : _GEN_1731; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1988 = unuse_way == 3'h1 ? valid_3_12 : _GEN_1732; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1989 = unuse_way == 3'h1 ? valid_3_13 : _GEN_1733; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1990 = unuse_way == 3'h1 ? valid_3_14 : _GEN_1734; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1991 = unuse_way == 3'h1 ? valid_3_15 : _GEN_1735; // @[i_cache.scala 30:26 85:34]
  wire  _GEN_1992 = 3'h4 == state ? 1'h0 : valid_0_0; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1993 = 3'h4 == state ? 1'h0 : valid_0_1; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1994 = 3'h4 == state ? 1'h0 : valid_0_2; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1995 = 3'h4 == state ? 1'h0 : valid_0_3; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1996 = 3'h4 == state ? 1'h0 : valid_0_4; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1997 = 3'h4 == state ? 1'h0 : valid_0_5; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1998 = 3'h4 == state ? 1'h0 : valid_0_6; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_1999 = 3'h4 == state ? 1'h0 : valid_0_7; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2000 = 3'h4 == state ? 1'h0 : valid_0_8; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2001 = 3'h4 == state ? 1'h0 : valid_0_9; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2002 = 3'h4 == state ? 1'h0 : valid_0_10; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2003 = 3'h4 == state ? 1'h0 : valid_0_11; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2004 = 3'h4 == state ? 1'h0 : valid_0_12; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2005 = 3'h4 == state ? 1'h0 : valid_0_13; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2006 = 3'h4 == state ? 1'h0 : valid_0_14; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2007 = 3'h4 == state ? 1'h0 : valid_0_15; // @[i_cache.scala 56:18 130:49 27:26]
  wire  _GEN_2008 = 3'h4 == state ? 1'h0 : valid_1_0; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2009 = 3'h4 == state ? 1'h0 : valid_1_1; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2010 = 3'h4 == state ? 1'h0 : valid_1_2; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2011 = 3'h4 == state ? 1'h0 : valid_1_3; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2012 = 3'h4 == state ? 1'h0 : valid_1_4; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2013 = 3'h4 == state ? 1'h0 : valid_1_5; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2014 = 3'h4 == state ? 1'h0 : valid_1_6; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2015 = 3'h4 == state ? 1'h0 : valid_1_7; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2016 = 3'h4 == state ? 1'h0 : valid_1_8; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2017 = 3'h4 == state ? 1'h0 : valid_1_9; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2018 = 3'h4 == state ? 1'h0 : valid_1_10; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2019 = 3'h4 == state ? 1'h0 : valid_1_11; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2020 = 3'h4 == state ? 1'h0 : valid_1_12; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2021 = 3'h4 == state ? 1'h0 : valid_1_13; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2022 = 3'h4 == state ? 1'h0 : valid_1_14; // @[i_cache.scala 56:18 131:49 28:26]
  wire  _GEN_2023 = 3'h4 == state ? 1'h0 : valid_1_15; // @[i_cache.scala 56:18 131:49 28:26]
  wire [2:0] _GEN_2024 = 3'h4 == state ? 3'h0 : state; // @[i_cache.scala 132:18 56:18 54:24]
  wire [2:0] _GEN_2025 = 3'h3 == state ? 3'h1 : _GEN_2024; // @[i_cache.scala 56:18 84:19]
  wire [511:0] _GEN_2026 = 3'h3 == state ? _GEN_1784 : ram_0_0; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2027 = 3'h3 == state ? _GEN_1785 : ram_0_1; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2028 = 3'h3 == state ? _GEN_1786 : ram_0_2; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2029 = 3'h3 == state ? _GEN_1787 : ram_0_3; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2030 = 3'h3 == state ? _GEN_1788 : ram_0_4; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2031 = 3'h3 == state ? _GEN_1789 : ram_0_5; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2032 = 3'h3 == state ? _GEN_1790 : ram_0_6; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2033 = 3'h3 == state ? _GEN_1791 : ram_0_7; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2034 = 3'h3 == state ? _GEN_1792 : ram_0_8; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2035 = 3'h3 == state ? _GEN_1793 : ram_0_9; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2036 = 3'h3 == state ? _GEN_1794 : ram_0_10; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2037 = 3'h3 == state ? _GEN_1795 : ram_0_11; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2038 = 3'h3 == state ? _GEN_1796 : ram_0_12; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2039 = 3'h3 == state ? _GEN_1797 : ram_0_13; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2040 = 3'h3 == state ? _GEN_1798 : ram_0_14; // @[i_cache.scala 56:18 19:24]
  wire [511:0] _GEN_2041 = 3'h3 == state ? _GEN_1799 : ram_0_15; // @[i_cache.scala 56:18 19:24]
  wire [31:0] _GEN_2042 = 3'h3 == state ? _GEN_1800 : tag_0_0; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2043 = 3'h3 == state ? _GEN_1801 : tag_0_1; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2044 = 3'h3 == state ? _GEN_1802 : tag_0_2; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2045 = 3'h3 == state ? _GEN_1803 : tag_0_3; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2046 = 3'h3 == state ? _GEN_1804 : tag_0_4; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2047 = 3'h3 == state ? _GEN_1805 : tag_0_5; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2048 = 3'h3 == state ? _GEN_1806 : tag_0_6; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2049 = 3'h3 == state ? _GEN_1807 : tag_0_7; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2050 = 3'h3 == state ? _GEN_1808 : tag_0_8; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2051 = 3'h3 == state ? _GEN_1809 : tag_0_9; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2052 = 3'h3 == state ? _GEN_1810 : tag_0_10; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2053 = 3'h3 == state ? _GEN_1811 : tag_0_11; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2054 = 3'h3 == state ? _GEN_1812 : tag_0_12; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2055 = 3'h3 == state ? _GEN_1813 : tag_0_13; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2056 = 3'h3 == state ? _GEN_1814 : tag_0_14; // @[i_cache.scala 56:18 23:24]
  wire [31:0] _GEN_2057 = 3'h3 == state ? _GEN_1815 : tag_0_15; // @[i_cache.scala 56:18 23:24]
  wire  _GEN_2058 = 3'h3 == state ? _GEN_1816 : _GEN_1992; // @[i_cache.scala 56:18]
  wire  _GEN_2059 = 3'h3 == state ? _GEN_1817 : _GEN_1993; // @[i_cache.scala 56:18]
  wire  _GEN_2060 = 3'h3 == state ? _GEN_1818 : _GEN_1994; // @[i_cache.scala 56:18]
  wire  _GEN_2061 = 3'h3 == state ? _GEN_1819 : _GEN_1995; // @[i_cache.scala 56:18]
  wire  _GEN_2062 = 3'h3 == state ? _GEN_1820 : _GEN_1996; // @[i_cache.scala 56:18]
  wire  _GEN_2063 = 3'h3 == state ? _GEN_1821 : _GEN_1997; // @[i_cache.scala 56:18]
  wire  _GEN_2064 = 3'h3 == state ? _GEN_1822 : _GEN_1998; // @[i_cache.scala 56:18]
  wire  _GEN_2065 = 3'h3 == state ? _GEN_1823 : _GEN_1999; // @[i_cache.scala 56:18]
  wire  _GEN_2066 = 3'h3 == state ? _GEN_1824 : _GEN_2000; // @[i_cache.scala 56:18]
  wire  _GEN_2067 = 3'h3 == state ? _GEN_1825 : _GEN_2001; // @[i_cache.scala 56:18]
  wire  _GEN_2068 = 3'h3 == state ? _GEN_1826 : _GEN_2002; // @[i_cache.scala 56:18]
  wire  _GEN_2069 = 3'h3 == state ? _GEN_1827 : _GEN_2003; // @[i_cache.scala 56:18]
  wire  _GEN_2070 = 3'h3 == state ? _GEN_1828 : _GEN_2004; // @[i_cache.scala 56:18]
  wire  _GEN_2071 = 3'h3 == state ? _GEN_1829 : _GEN_2005; // @[i_cache.scala 56:18]
  wire  _GEN_2072 = 3'h3 == state ? _GEN_1830 : _GEN_2006; // @[i_cache.scala 56:18]
  wire  _GEN_2073 = 3'h3 == state ? _GEN_1831 : _GEN_2007; // @[i_cache.scala 56:18]
  wire [7:0] _GEN_2074 = 3'h3 == state ? _GEN_1832 : quene_0; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2075 = 3'h3 == state ? _GEN_1833 : quene_1; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2076 = 3'h3 == state ? _GEN_1834 : quene_2; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2077 = 3'h3 == state ? _GEN_1835 : quene_3; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2078 = 3'h3 == state ? _GEN_1836 : quene_4; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2079 = 3'h3 == state ? _GEN_1837 : quene_5; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2080 = 3'h3 == state ? _GEN_1838 : quene_6; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2081 = 3'h3 == state ? _GEN_1839 : quene_7; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2082 = 3'h3 == state ? _GEN_1840 : quene_8; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2083 = 3'h3 == state ? _GEN_1841 : quene_9; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2084 = 3'h3 == state ? _GEN_1842 : quene_10; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2085 = 3'h3 == state ? _GEN_1843 : quene_11; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2086 = 3'h3 == state ? _GEN_1844 : quene_12; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2087 = 3'h3 == state ? _GEN_1845 : quene_13; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2088 = 3'h3 == state ? _GEN_1846 : quene_14; // @[i_cache.scala 56:18 40:24]
  wire [7:0] _GEN_2089 = 3'h3 == state ? _GEN_1847 : quene_15; // @[i_cache.scala 56:18 40:24]
  wire [511:0] _GEN_2090 = 3'h3 == state ? _GEN_1848 : ram_1_0; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2091 = 3'h3 == state ? _GEN_1849 : ram_1_1; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2092 = 3'h3 == state ? _GEN_1850 : ram_1_2; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2093 = 3'h3 == state ? _GEN_1851 : ram_1_3; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2094 = 3'h3 == state ? _GEN_1852 : ram_1_4; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2095 = 3'h3 == state ? _GEN_1853 : ram_1_5; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2096 = 3'h3 == state ? _GEN_1854 : ram_1_6; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2097 = 3'h3 == state ? _GEN_1855 : ram_1_7; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2098 = 3'h3 == state ? _GEN_1856 : ram_1_8; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2099 = 3'h3 == state ? _GEN_1857 : ram_1_9; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2100 = 3'h3 == state ? _GEN_1858 : ram_1_10; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2101 = 3'h3 == state ? _GEN_1859 : ram_1_11; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2102 = 3'h3 == state ? _GEN_1860 : ram_1_12; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2103 = 3'h3 == state ? _GEN_1861 : ram_1_13; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2104 = 3'h3 == state ? _GEN_1862 : ram_1_14; // @[i_cache.scala 56:18 20:24]
  wire [511:0] _GEN_2105 = 3'h3 == state ? _GEN_1863 : ram_1_15; // @[i_cache.scala 56:18 20:24]
  wire [31:0] _GEN_2106 = 3'h3 == state ? _GEN_1864 : tag_1_0; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2107 = 3'h3 == state ? _GEN_1865 : tag_1_1; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2108 = 3'h3 == state ? _GEN_1866 : tag_1_2; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2109 = 3'h3 == state ? _GEN_1867 : tag_1_3; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2110 = 3'h3 == state ? _GEN_1868 : tag_1_4; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2111 = 3'h3 == state ? _GEN_1869 : tag_1_5; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2112 = 3'h3 == state ? _GEN_1870 : tag_1_6; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2113 = 3'h3 == state ? _GEN_1871 : tag_1_7; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2114 = 3'h3 == state ? _GEN_1872 : tag_1_8; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2115 = 3'h3 == state ? _GEN_1873 : tag_1_9; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2116 = 3'h3 == state ? _GEN_1874 : tag_1_10; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2117 = 3'h3 == state ? _GEN_1875 : tag_1_11; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2118 = 3'h3 == state ? _GEN_1876 : tag_1_12; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2119 = 3'h3 == state ? _GEN_1877 : tag_1_13; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2120 = 3'h3 == state ? _GEN_1878 : tag_1_14; // @[i_cache.scala 56:18 24:24]
  wire [31:0] _GEN_2121 = 3'h3 == state ? _GEN_1879 : tag_1_15; // @[i_cache.scala 56:18 24:24]
  wire  _GEN_2122 = 3'h3 == state ? _GEN_1880 : _GEN_2008; // @[i_cache.scala 56:18]
  wire  _GEN_2123 = 3'h3 == state ? _GEN_1881 : _GEN_2009; // @[i_cache.scala 56:18]
  wire  _GEN_2124 = 3'h3 == state ? _GEN_1882 : _GEN_2010; // @[i_cache.scala 56:18]
  wire  _GEN_2125 = 3'h3 == state ? _GEN_1883 : _GEN_2011; // @[i_cache.scala 56:18]
  wire  _GEN_2126 = 3'h3 == state ? _GEN_1884 : _GEN_2012; // @[i_cache.scala 56:18]
  wire  _GEN_2127 = 3'h3 == state ? _GEN_1885 : _GEN_2013; // @[i_cache.scala 56:18]
  wire  _GEN_2128 = 3'h3 == state ? _GEN_1886 : _GEN_2014; // @[i_cache.scala 56:18]
  wire  _GEN_2129 = 3'h3 == state ? _GEN_1887 : _GEN_2015; // @[i_cache.scala 56:18]
  wire  _GEN_2130 = 3'h3 == state ? _GEN_1888 : _GEN_2016; // @[i_cache.scala 56:18]
  wire  _GEN_2131 = 3'h3 == state ? _GEN_1889 : _GEN_2017; // @[i_cache.scala 56:18]
  wire  _GEN_2132 = 3'h3 == state ? _GEN_1890 : _GEN_2018; // @[i_cache.scala 56:18]
  wire  _GEN_2133 = 3'h3 == state ? _GEN_1891 : _GEN_2019; // @[i_cache.scala 56:18]
  wire  _GEN_2134 = 3'h3 == state ? _GEN_1892 : _GEN_2020; // @[i_cache.scala 56:18]
  wire  _GEN_2135 = 3'h3 == state ? _GEN_1893 : _GEN_2021; // @[i_cache.scala 56:18]
  wire  _GEN_2136 = 3'h3 == state ? _GEN_1894 : _GEN_2022; // @[i_cache.scala 56:18]
  wire  _GEN_2137 = 3'h3 == state ? _GEN_1895 : _GEN_2023; // @[i_cache.scala 56:18]
  wire [511:0] _GEN_2138 = 3'h3 == state ? _GEN_1896 : ram_2_0; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2139 = 3'h3 == state ? _GEN_1897 : ram_2_1; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2140 = 3'h3 == state ? _GEN_1898 : ram_2_2; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2141 = 3'h3 == state ? _GEN_1899 : ram_2_3; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2142 = 3'h3 == state ? _GEN_1900 : ram_2_4; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2143 = 3'h3 == state ? _GEN_1901 : ram_2_5; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2144 = 3'h3 == state ? _GEN_1902 : ram_2_6; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2145 = 3'h3 == state ? _GEN_1903 : ram_2_7; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2146 = 3'h3 == state ? _GEN_1904 : ram_2_8; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2147 = 3'h3 == state ? _GEN_1905 : ram_2_9; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2148 = 3'h3 == state ? _GEN_1906 : ram_2_10; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2149 = 3'h3 == state ? _GEN_1907 : ram_2_11; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2150 = 3'h3 == state ? _GEN_1908 : ram_2_12; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2151 = 3'h3 == state ? _GEN_1909 : ram_2_13; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2152 = 3'h3 == state ? _GEN_1910 : ram_2_14; // @[i_cache.scala 56:18 21:24]
  wire [511:0] _GEN_2153 = 3'h3 == state ? _GEN_1911 : ram_2_15; // @[i_cache.scala 56:18 21:24]
  wire [31:0] _GEN_2154 = 3'h3 == state ? _GEN_1912 : tag_2_0; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2155 = 3'h3 == state ? _GEN_1913 : tag_2_1; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2156 = 3'h3 == state ? _GEN_1914 : tag_2_2; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2157 = 3'h3 == state ? _GEN_1915 : tag_2_3; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2158 = 3'h3 == state ? _GEN_1916 : tag_2_4; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2159 = 3'h3 == state ? _GEN_1917 : tag_2_5; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2160 = 3'h3 == state ? _GEN_1918 : tag_2_6; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2161 = 3'h3 == state ? _GEN_1919 : tag_2_7; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2162 = 3'h3 == state ? _GEN_1920 : tag_2_8; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2163 = 3'h3 == state ? _GEN_1921 : tag_2_9; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2164 = 3'h3 == state ? _GEN_1922 : tag_2_10; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2165 = 3'h3 == state ? _GEN_1923 : tag_2_11; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2166 = 3'h3 == state ? _GEN_1924 : tag_2_12; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2167 = 3'h3 == state ? _GEN_1925 : tag_2_13; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2168 = 3'h3 == state ? _GEN_1926 : tag_2_14; // @[i_cache.scala 56:18 25:24]
  wire [31:0] _GEN_2169 = 3'h3 == state ? _GEN_1927 : tag_2_15; // @[i_cache.scala 56:18 25:24]
  wire  _GEN_2170 = 3'h3 == state ? _GEN_1928 : valid_2_0; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2171 = 3'h3 == state ? _GEN_1929 : valid_2_1; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2172 = 3'h3 == state ? _GEN_1930 : valid_2_2; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2173 = 3'h3 == state ? _GEN_1931 : valid_2_3; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2174 = 3'h3 == state ? _GEN_1932 : valid_2_4; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2175 = 3'h3 == state ? _GEN_1933 : valid_2_5; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2176 = 3'h3 == state ? _GEN_1934 : valid_2_6; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2177 = 3'h3 == state ? _GEN_1935 : valid_2_7; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2178 = 3'h3 == state ? _GEN_1936 : valid_2_8; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2179 = 3'h3 == state ? _GEN_1937 : valid_2_9; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2180 = 3'h3 == state ? _GEN_1938 : valid_2_10; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2181 = 3'h3 == state ? _GEN_1939 : valid_2_11; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2182 = 3'h3 == state ? _GEN_1940 : valid_2_12; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2183 = 3'h3 == state ? _GEN_1941 : valid_2_13; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2184 = 3'h3 == state ? _GEN_1942 : valid_2_14; // @[i_cache.scala 56:18 29:26]
  wire  _GEN_2185 = 3'h3 == state ? _GEN_1943 : valid_2_15; // @[i_cache.scala 56:18 29:26]
  wire [511:0] _GEN_2186 = 3'h3 == state ? _GEN_1944 : ram_3_0; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2187 = 3'h3 == state ? _GEN_1945 : ram_3_1; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2188 = 3'h3 == state ? _GEN_1946 : ram_3_2; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2189 = 3'h3 == state ? _GEN_1947 : ram_3_3; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2190 = 3'h3 == state ? _GEN_1948 : ram_3_4; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2191 = 3'h3 == state ? _GEN_1949 : ram_3_5; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2192 = 3'h3 == state ? _GEN_1950 : ram_3_6; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2193 = 3'h3 == state ? _GEN_1951 : ram_3_7; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2194 = 3'h3 == state ? _GEN_1952 : ram_3_8; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2195 = 3'h3 == state ? _GEN_1953 : ram_3_9; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2196 = 3'h3 == state ? _GEN_1954 : ram_3_10; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2197 = 3'h3 == state ? _GEN_1955 : ram_3_11; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2198 = 3'h3 == state ? _GEN_1956 : ram_3_12; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2199 = 3'h3 == state ? _GEN_1957 : ram_3_13; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2200 = 3'h3 == state ? _GEN_1958 : ram_3_14; // @[i_cache.scala 56:18 22:24]
  wire [511:0] _GEN_2201 = 3'h3 == state ? _GEN_1959 : ram_3_15; // @[i_cache.scala 56:18 22:24]
  wire [31:0] _GEN_2202 = 3'h3 == state ? _GEN_1960 : tag_3_0; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2203 = 3'h3 == state ? _GEN_1961 : tag_3_1; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2204 = 3'h3 == state ? _GEN_1962 : tag_3_2; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2205 = 3'h3 == state ? _GEN_1963 : tag_3_3; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2206 = 3'h3 == state ? _GEN_1964 : tag_3_4; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2207 = 3'h3 == state ? _GEN_1965 : tag_3_5; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2208 = 3'h3 == state ? _GEN_1966 : tag_3_6; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2209 = 3'h3 == state ? _GEN_1967 : tag_3_7; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2210 = 3'h3 == state ? _GEN_1968 : tag_3_8; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2211 = 3'h3 == state ? _GEN_1969 : tag_3_9; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2212 = 3'h3 == state ? _GEN_1970 : tag_3_10; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2213 = 3'h3 == state ? _GEN_1971 : tag_3_11; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2214 = 3'h3 == state ? _GEN_1972 : tag_3_12; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2215 = 3'h3 == state ? _GEN_1973 : tag_3_13; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2216 = 3'h3 == state ? _GEN_1974 : tag_3_14; // @[i_cache.scala 56:18 26:24]
  wire [31:0] _GEN_2217 = 3'h3 == state ? _GEN_1975 : tag_3_15; // @[i_cache.scala 56:18 26:24]
  wire  _GEN_2218 = 3'h3 == state ? _GEN_1976 : valid_3_0; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2219 = 3'h3 == state ? _GEN_1977 : valid_3_1; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2220 = 3'h3 == state ? _GEN_1978 : valid_3_2; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2221 = 3'h3 == state ? _GEN_1979 : valid_3_3; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2222 = 3'h3 == state ? _GEN_1980 : valid_3_4; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2223 = 3'h3 == state ? _GEN_1981 : valid_3_5; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2224 = 3'h3 == state ? _GEN_1982 : valid_3_6; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2225 = 3'h3 == state ? _GEN_1983 : valid_3_7; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2226 = 3'h3 == state ? _GEN_1984 : valid_3_8; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2227 = 3'h3 == state ? _GEN_1985 : valid_3_9; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2228 = 3'h3 == state ? _GEN_1986 : valid_3_10; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2229 = 3'h3 == state ? _GEN_1987 : valid_3_11; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2230 = 3'h3 == state ? _GEN_1988 : valid_3_12; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2231 = 3'h3 == state ? _GEN_1989 : valid_3_13; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2232 = 3'h3 == state ? _GEN_1990 : valid_3_14; // @[i_cache.scala 56:18 30:26]
  wire  _GEN_2233 = 3'h3 == state ? _GEN_1991 : valid_3_15; // @[i_cache.scala 56:18 30:26]
  wire [511:0] _GEN_2889 = 4'h1 == index ? ram_0_1 : ram_0_0; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2890 = 4'h2 == index ? ram_0_2 : _GEN_2889; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2891 = 4'h3 == index ? ram_0_3 : _GEN_2890; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2892 = 4'h4 == index ? ram_0_4 : _GEN_2891; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2893 = 4'h5 == index ? ram_0_5 : _GEN_2892; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2894 = 4'h6 == index ? ram_0_6 : _GEN_2893; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2895 = 4'h7 == index ? ram_0_7 : _GEN_2894; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2896 = 4'h8 == index ? ram_0_8 : _GEN_2895; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2897 = 4'h9 == index ? ram_0_9 : _GEN_2896; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2898 = 4'ha == index ? ram_0_10 : _GEN_2897; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2899 = 4'hb == index ? ram_0_11 : _GEN_2898; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2900 = 4'hc == index ? ram_0_12 : _GEN_2899; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2901 = 4'hd == index ? ram_0_13 : _GEN_2900; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2902 = 4'he == index ? ram_0_14 : _GEN_2901; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _GEN_2903 = 4'hf == index ? ram_0_15 : _GEN_2902; // @[i_cache.scala 153:{55,55}]
  wire [511:0] _io_to_ifu_rdata_T = _GEN_2903 >> shift_bit; // @[i_cache.scala 153:55]
  wire [511:0] _GEN_2905 = 4'h1 == index ? ram_1_1 : ram_1_0; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2906 = 4'h2 == index ? ram_1_2 : _GEN_2905; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2907 = 4'h3 == index ? ram_1_3 : _GEN_2906; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2908 = 4'h4 == index ? ram_1_4 : _GEN_2907; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2909 = 4'h5 == index ? ram_1_5 : _GEN_2908; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2910 = 4'h6 == index ? ram_1_6 : _GEN_2909; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2911 = 4'h7 == index ? ram_1_7 : _GEN_2910; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2912 = 4'h8 == index ? ram_1_8 : _GEN_2911; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2913 = 4'h9 == index ? ram_1_9 : _GEN_2912; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2914 = 4'ha == index ? ram_1_10 : _GEN_2913; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2915 = 4'hb == index ? ram_1_11 : _GEN_2914; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2916 = 4'hc == index ? ram_1_12 : _GEN_2915; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2917 = 4'hd == index ? ram_1_13 : _GEN_2916; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2918 = 4'he == index ? ram_1_14 : _GEN_2917; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _GEN_2919 = 4'hf == index ? ram_1_15 : _GEN_2918; // @[i_cache.scala 153:{95,95}]
  wire [511:0] _io_to_ifu_rdata_T_1 = _GEN_2919 >> shift_bit; // @[i_cache.scala 153:95]
  wire [511:0] _GEN_2921 = 4'h1 == index ? ram_2_1 : ram_2_0; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2922 = 4'h2 == index ? ram_2_2 : _GEN_2921; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2923 = 4'h3 == index ? ram_2_3 : _GEN_2922; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2924 = 4'h4 == index ? ram_2_4 : _GEN_2923; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2925 = 4'h5 == index ? ram_2_5 : _GEN_2924; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2926 = 4'h6 == index ? ram_2_6 : _GEN_2925; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2927 = 4'h7 == index ? ram_2_7 : _GEN_2926; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2928 = 4'h8 == index ? ram_2_8 : _GEN_2927; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2929 = 4'h9 == index ? ram_2_9 : _GEN_2928; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2930 = 4'ha == index ? ram_2_10 : _GEN_2929; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2931 = 4'hb == index ? ram_2_11 : _GEN_2930; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2932 = 4'hc == index ? ram_2_12 : _GEN_2931; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2933 = 4'hd == index ? ram_2_13 : _GEN_2932; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2934 = 4'he == index ? ram_2_14 : _GEN_2933; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _GEN_2935 = 4'hf == index ? ram_2_15 : _GEN_2934; // @[i_cache.scala 153:{135,135}]
  wire [511:0] _io_to_ifu_rdata_T_2 = _GEN_2935 >> shift_bit; // @[i_cache.scala 153:135]
  wire [511:0] _GEN_2937 = 4'h1 == index ? ram_3_1 : ram_3_0; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2938 = 4'h2 == index ? ram_3_2 : _GEN_2937; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2939 = 4'h3 == index ? ram_3_3 : _GEN_2938; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2940 = 4'h4 == index ? ram_3_4 : _GEN_2939; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2941 = 4'h5 == index ? ram_3_5 : _GEN_2940; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2942 = 4'h6 == index ? ram_3_6 : _GEN_2941; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2943 = 4'h7 == index ? ram_3_7 : _GEN_2942; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2944 = 4'h8 == index ? ram_3_8 : _GEN_2943; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2945 = 4'h9 == index ? ram_3_9 : _GEN_2944; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2946 = 4'ha == index ? ram_3_10 : _GEN_2945; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2947 = 4'hb == index ? ram_3_11 : _GEN_2946; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2948 = 4'hc == index ? ram_3_12 : _GEN_2947; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2949 = 4'hd == index ? ram_3_13 : _GEN_2948; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2950 = 4'he == index ? ram_3_14 : _GEN_2949; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _GEN_2951 = 4'hf == index ? ram_3_15 : _GEN_2950; // @[i_cache.scala 153:{162,162}]
  wire [511:0] _io_to_ifu_rdata_T_3 = _GEN_2951 >> shift_bit; // @[i_cache.scala 153:162]
  wire [511:0] _io_to_ifu_rdata_T_4 = way2_hit ? _io_to_ifu_rdata_T_2 : _io_to_ifu_rdata_T_3; // @[i_cache.scala 153:112]
  wire [511:0] _io_to_ifu_rdata_T_5 = way1_hit ? _io_to_ifu_rdata_T_1 : _io_to_ifu_rdata_T_4; // @[i_cache.scala 153:72]
  wire [511:0] _io_to_ifu_rdata_T_6 = way0_hit ? _io_to_ifu_rdata_T : _io_to_ifu_rdata_T_5; // @[i_cache.scala 153:32]
  wire  _T_19 = state == 3'h2; // @[i_cache.scala 160:21]
  wire [63:0] _GEN_3105 = {{32'd0}, io_from_ifu_araddr}; // @[i_cache.scala 169:49]
  wire [63:0] _io_to_axi_araddr_T = _GEN_3105 & 64'hffffffffffffffc0; // @[i_cache.scala 169:49]
  wire [63:0] _GEN_2954 = state == 3'h2 ? _io_to_axi_araddr_T : {{32'd0}, io_from_ifu_araddr}; // @[i_cache.scala 160:29 169:26 193:26]
  wire [2:0] _GEN_2955 = state == 3'h2 ? 3'h7 : 3'h0; // @[i_cache.scala 160:29 170:25 195:25]
  wire [63:0] _GEN_2959 = state == 3'h1 ? {{32'd0}, io_from_ifu_araddr} : _GEN_2954; // @[i_cache.scala 136:25 138:26]
  wire [2:0] _GEN_2960 = state == 3'h1 ? 3'h0 : _GEN_2955; // @[i_cache.scala 136:25 139:25]
  wire [511:0] _GEN_2964 = state == 3'h1 ? _io_to_ifu_rdata_T_6 : 512'h0; // @[i_cache.scala 136:25 153:25]
  assign io_to_ifu_rdata = _GEN_2964[63:0];
  assign io_to_ifu_rlast = state == 3'h1 & _T_4; // @[i_cache.scala 136:25 156:25]
  assign io_to_ifu_rvalid = state == 3'h1 & _T_4; // @[i_cache.scala 136:25 155:26]
  assign io_to_axi_araddr = _GEN_2959[31:0];
  assign io_to_axi_arlen = {{5'd0}, _GEN_2960};
  assign io_to_axi_arvalid = state == 3'h1 ? 1'h0 : _T_19; // @[i_cache.scala 136:25 137:27]
  assign io_to_axi_rready = state == 3'h1 ? 1'h0 : io_from_ifu_rready; // @[i_cache.scala 136:25 142:26]
  assign io_cache_init = state == 3'h4; // @[i_cache.scala 209:27]
  always @(posedge clock) begin
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_0 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_0 <= _GEN_2026;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_1 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_1 <= _GEN_2027;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_2 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_2 <= _GEN_2028;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_3 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_3 <= _GEN_2029;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_4 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_4 <= _GEN_2030;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_5 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_5 <= _GEN_2031;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_6 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_6 <= _GEN_2032;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_7 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_7 <= _GEN_2033;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_8 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_8 <= _GEN_2034;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_9 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_9 <= _GEN_2035;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_10 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_10 <= _GEN_2036;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_11 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_11 <= _GEN_2037;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_12 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_12 <= _GEN_2038;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_13 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_13 <= _GEN_2039;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_14 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_14 <= _GEN_2040;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_15 <= 512'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_0_15 <= _GEN_2041;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_0 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_0 <= _GEN_2090;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_1 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_1 <= _GEN_2091;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_2 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_2 <= _GEN_2092;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_3 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_3 <= _GEN_2093;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_4 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_4 <= _GEN_2094;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_5 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_5 <= _GEN_2095;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_6 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_6 <= _GEN_2096;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_7 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_7 <= _GEN_2097;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_8 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_8 <= _GEN_2098;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_9 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_9 <= _GEN_2099;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_10 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_10 <= _GEN_2100;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_11 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_11 <= _GEN_2101;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_12 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_12 <= _GEN_2102;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_13 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_13 <= _GEN_2103;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_14 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_14 <= _GEN_2104;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_15 <= 512'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_1_15 <= _GEN_2105;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_0 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_0 <= _GEN_2138;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_1 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_1 <= _GEN_2139;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_2 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_2 <= _GEN_2140;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_3 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_3 <= _GEN_2141;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_4 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_4 <= _GEN_2142;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_5 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_5 <= _GEN_2143;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_6 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_6 <= _GEN_2144;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_7 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_7 <= _GEN_2145;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_8 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_8 <= _GEN_2146;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_9 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_9 <= _GEN_2147;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_10 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_10 <= _GEN_2148;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_11 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_11 <= _GEN_2149;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_12 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_12 <= _GEN_2150;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_13 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_13 <= _GEN_2151;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_14 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_14 <= _GEN_2152;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_15 <= 512'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_2_15 <= _GEN_2153;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_0 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_0 <= _GEN_2186;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_1 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_1 <= _GEN_2187;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_2 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_2 <= _GEN_2188;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_3 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_3 <= _GEN_2189;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_4 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_4 <= _GEN_2190;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_5 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_5 <= _GEN_2191;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_6 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_6 <= _GEN_2192;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_7 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_7 <= _GEN_2193;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_8 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_8 <= _GEN_2194;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_9 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_9 <= _GEN_2195;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_10 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_10 <= _GEN_2196;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_11 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_11 <= _GEN_2197;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_12 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_12 <= _GEN_2198;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_13 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_13 <= _GEN_2199;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_14 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_14 <= _GEN_2200;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_15 <= 512'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          ram_3_15 <= _GEN_2201;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_0 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_0 <= _GEN_2042;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_1 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_1 <= _GEN_2043;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_2 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_2 <= _GEN_2044;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_3 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_3 <= _GEN_2045;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_4 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_4 <= _GEN_2046;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_5 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_5 <= _GEN_2047;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_6 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_6 <= _GEN_2048;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_7 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_7 <= _GEN_2049;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_8 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_8 <= _GEN_2050;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_9 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_9 <= _GEN_2051;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_10 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_10 <= _GEN_2052;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_11 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_11 <= _GEN_2053;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_12 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_12 <= _GEN_2054;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_13 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_13 <= _GEN_2055;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_14 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_14 <= _GEN_2056;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_15 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_0_15 <= _GEN_2057;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_0 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_0 <= _GEN_2106;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_1 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_1 <= _GEN_2107;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_2 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_2 <= _GEN_2108;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_3 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_3 <= _GEN_2109;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_4 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_4 <= _GEN_2110;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_5 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_5 <= _GEN_2111;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_6 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_6 <= _GEN_2112;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_7 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_7 <= _GEN_2113;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_8 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_8 <= _GEN_2114;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_9 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_9 <= _GEN_2115;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_10 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_10 <= _GEN_2116;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_11 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_11 <= _GEN_2117;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_12 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_12 <= _GEN_2118;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_13 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_13 <= _GEN_2119;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_14 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_14 <= _GEN_2120;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_15 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_1_15 <= _GEN_2121;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_0 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_0 <= _GEN_2154;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_1 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_1 <= _GEN_2155;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_2 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_2 <= _GEN_2156;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_3 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_3 <= _GEN_2157;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_4 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_4 <= _GEN_2158;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_5 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_5 <= _GEN_2159;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_6 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_6 <= _GEN_2160;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_7 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_7 <= _GEN_2161;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_8 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_8 <= _GEN_2162;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_9 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_9 <= _GEN_2163;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_10 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_10 <= _GEN_2164;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_11 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_11 <= _GEN_2165;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_12 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_12 <= _GEN_2166;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_13 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_13 <= _GEN_2167;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_14 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_14 <= _GEN_2168;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_15 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_2_15 <= _GEN_2169;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_0 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_0 <= _GEN_2202;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_1 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_1 <= _GEN_2203;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_2 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_2 <= _GEN_2204;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_3 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_3 <= _GEN_2205;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_4 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_4 <= _GEN_2206;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_5 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_5 <= _GEN_2207;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_6 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_6 <= _GEN_2208;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_7 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_7 <= _GEN_2209;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_8 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_8 <= _GEN_2210;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_9 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_9 <= _GEN_2211;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_10 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_10 <= _GEN_2212;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_11 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_11 <= _GEN_2213;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_12 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_12 <= _GEN_2214;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_13 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_13 <= _GEN_2215;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_14 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_14 <= _GEN_2216;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_15 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          tag_3_15 <= _GEN_2217;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_0 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_0 <= _GEN_2058;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_1 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_1 <= _GEN_2059;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_2 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_2 <= _GEN_2060;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_3 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_3 <= _GEN_2061;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_4 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_4 <= _GEN_2062;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_5 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_5 <= _GEN_2063;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_6 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_6 <= _GEN_2064;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_7 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_7 <= _GEN_2065;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_8 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_8 <= _GEN_2066;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_9 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_9 <= _GEN_2067;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_10 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_10 <= _GEN_2068;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_11 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_11 <= _GEN_2069;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_12 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_12 <= _GEN_2070;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_13 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_13 <= _GEN_2071;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_14 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_14 <= _GEN_2072;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_15 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_0_15 <= _GEN_2073;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_0 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_0 <= _GEN_2122;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_1 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_1 <= _GEN_2123;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_2 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_2 <= _GEN_2124;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_3 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_3 <= _GEN_2125;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_4 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_4 <= _GEN_2126;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_5 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_5 <= _GEN_2127;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_6 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_6 <= _GEN_2128;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_7 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_7 <= _GEN_2129;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_8 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_8 <= _GEN_2130;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_9 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_9 <= _GEN_2131;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_10 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_10 <= _GEN_2132;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_11 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_11 <= _GEN_2133;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_12 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_12 <= _GEN_2134;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_13 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_13 <= _GEN_2135;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_14 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_14 <= _GEN_2136;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_15 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_1_15 <= _GEN_2137;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_0 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_0 <= _GEN_2170;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_1 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_1 <= _GEN_2171;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_2 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_2 <= _GEN_2172;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_3 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_3 <= _GEN_2173;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_4 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_4 <= _GEN_2174;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_5 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_5 <= _GEN_2175;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_6 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_6 <= _GEN_2176;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_7 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_7 <= _GEN_2177;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_8 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_8 <= _GEN_2178;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_9 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_9 <= _GEN_2179;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_10 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_10 <= _GEN_2180;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_11 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_11 <= _GEN_2181;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_12 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_12 <= _GEN_2182;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_13 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_13 <= _GEN_2183;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_14 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_14 <= _GEN_2184;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_15 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_2_15 <= _GEN_2185;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_0 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_0 <= _GEN_2218;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_1 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_1 <= _GEN_2219;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_2 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_2 <= _GEN_2220;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_3 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_3 <= _GEN_2221;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_4 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_4 <= _GEN_2222;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_5 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_5 <= _GEN_2223;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_6 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_6 <= _GEN_2224;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_7 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_7 <= _GEN_2225;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_8 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_8 <= _GEN_2226;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_9 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_9 <= _GEN_2227;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_10 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_10 <= _GEN_2228;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_11 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_11 <= _GEN_2229;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_12 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_12 <= _GEN_2230;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_13 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_13 <= _GEN_2231;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_14 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_14 <= _GEN_2232;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_15 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          valid_3_15 <= _GEN_2233;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_0 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_0 <= _GEN_142;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_1 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_1 <= _GEN_143;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_2 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_2 <= _GEN_144;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_3 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_3 <= _GEN_145;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_4 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_4 <= _GEN_146;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_5 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_5 <= _GEN_147;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_6 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_6 <= _GEN_148;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 38:31]
      receive_data_7 <= 64'h0; // @[i_cache.scala 38:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (3'h2 == state) begin // @[i_cache.scala 56:18]
          receive_data_7 <= _GEN_149;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 39:30]
      receive_num <= 3'h0; // @[i_cache.scala 39:30]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (3'h1 == state) begin // @[i_cache.scala 56:18]
        if (!(way0_hit | way1_hit | way2_hit | way3_hit)) begin // @[i_cache.scala 65:57]
          receive_num <= 3'h0; // @[i_cache.scala 71:29]
        end
      end else if (3'h2 == state) begin // @[i_cache.scala 56:18]
        receive_num <= _GEN_150;
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_0 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_0 <= _GEN_2074;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_1 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_1 <= _GEN_2075;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_2 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_2 <= _GEN_2076;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_3 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_3 <= _GEN_2077;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_4 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_4 <= _GEN_2078;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_5 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_5 <= _GEN_2079;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_6 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_6 <= _GEN_2080;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_7 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_7 <= _GEN_2081;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_8 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_8 <= _GEN_2082;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_9 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_9 <= _GEN_2083;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_10 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_10 <= _GEN_2084;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_11 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_11 <= _GEN_2085;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_12 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_12 <= _GEN_2086;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_13 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_13 <= _GEN_2087;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_14 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_14 <= _GEN_2088;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:24]
      quene_15 <= 8'h0; // @[i_cache.scala 40:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 56:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 56:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 56:18]
          quene_15 <= _GEN_2089;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 54:24]
      state <= 3'h0; // @[i_cache.scala 54:24]
    end else if (3'h0 == state) begin // @[i_cache.scala 56:18]
      if (io_clear_cache) begin // @[i_cache.scala 58:33]
        state <= 3'h4; // @[i_cache.scala 59:23]
      end else if (io_from_ifu_arvalid) begin // @[i_cache.scala 60:44]
        state <= 3'h1; // @[i_cache.scala 61:23]
      end
    end else if (3'h1 == state) begin // @[i_cache.scala 56:18]
      if (way0_hit | way1_hit | way2_hit | way3_hit) begin // @[i_cache.scala 65:57]
        state <= _GEN_130;
      end else begin
        state <= 3'h2; // @[i_cache.scala 70:23]
      end
    end else if (3'h2 == state) begin // @[i_cache.scala 56:18]
      state <= _GEN_151;
    end else begin
      state <= _GEN_2025;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  ram_0_0 = _RAND_0[511:0];
  _RAND_1 = {16{`RANDOM}};
  ram_0_1 = _RAND_1[511:0];
  _RAND_2 = {16{`RANDOM}};
  ram_0_2 = _RAND_2[511:0];
  _RAND_3 = {16{`RANDOM}};
  ram_0_3 = _RAND_3[511:0];
  _RAND_4 = {16{`RANDOM}};
  ram_0_4 = _RAND_4[511:0];
  _RAND_5 = {16{`RANDOM}};
  ram_0_5 = _RAND_5[511:0];
  _RAND_6 = {16{`RANDOM}};
  ram_0_6 = _RAND_6[511:0];
  _RAND_7 = {16{`RANDOM}};
  ram_0_7 = _RAND_7[511:0];
  _RAND_8 = {16{`RANDOM}};
  ram_0_8 = _RAND_8[511:0];
  _RAND_9 = {16{`RANDOM}};
  ram_0_9 = _RAND_9[511:0];
  _RAND_10 = {16{`RANDOM}};
  ram_0_10 = _RAND_10[511:0];
  _RAND_11 = {16{`RANDOM}};
  ram_0_11 = _RAND_11[511:0];
  _RAND_12 = {16{`RANDOM}};
  ram_0_12 = _RAND_12[511:0];
  _RAND_13 = {16{`RANDOM}};
  ram_0_13 = _RAND_13[511:0];
  _RAND_14 = {16{`RANDOM}};
  ram_0_14 = _RAND_14[511:0];
  _RAND_15 = {16{`RANDOM}};
  ram_0_15 = _RAND_15[511:0];
  _RAND_16 = {16{`RANDOM}};
  ram_1_0 = _RAND_16[511:0];
  _RAND_17 = {16{`RANDOM}};
  ram_1_1 = _RAND_17[511:0];
  _RAND_18 = {16{`RANDOM}};
  ram_1_2 = _RAND_18[511:0];
  _RAND_19 = {16{`RANDOM}};
  ram_1_3 = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  ram_1_4 = _RAND_20[511:0];
  _RAND_21 = {16{`RANDOM}};
  ram_1_5 = _RAND_21[511:0];
  _RAND_22 = {16{`RANDOM}};
  ram_1_6 = _RAND_22[511:0];
  _RAND_23 = {16{`RANDOM}};
  ram_1_7 = _RAND_23[511:0];
  _RAND_24 = {16{`RANDOM}};
  ram_1_8 = _RAND_24[511:0];
  _RAND_25 = {16{`RANDOM}};
  ram_1_9 = _RAND_25[511:0];
  _RAND_26 = {16{`RANDOM}};
  ram_1_10 = _RAND_26[511:0];
  _RAND_27 = {16{`RANDOM}};
  ram_1_11 = _RAND_27[511:0];
  _RAND_28 = {16{`RANDOM}};
  ram_1_12 = _RAND_28[511:0];
  _RAND_29 = {16{`RANDOM}};
  ram_1_13 = _RAND_29[511:0];
  _RAND_30 = {16{`RANDOM}};
  ram_1_14 = _RAND_30[511:0];
  _RAND_31 = {16{`RANDOM}};
  ram_1_15 = _RAND_31[511:0];
  _RAND_32 = {16{`RANDOM}};
  ram_2_0 = _RAND_32[511:0];
  _RAND_33 = {16{`RANDOM}};
  ram_2_1 = _RAND_33[511:0];
  _RAND_34 = {16{`RANDOM}};
  ram_2_2 = _RAND_34[511:0];
  _RAND_35 = {16{`RANDOM}};
  ram_2_3 = _RAND_35[511:0];
  _RAND_36 = {16{`RANDOM}};
  ram_2_4 = _RAND_36[511:0];
  _RAND_37 = {16{`RANDOM}};
  ram_2_5 = _RAND_37[511:0];
  _RAND_38 = {16{`RANDOM}};
  ram_2_6 = _RAND_38[511:0];
  _RAND_39 = {16{`RANDOM}};
  ram_2_7 = _RAND_39[511:0];
  _RAND_40 = {16{`RANDOM}};
  ram_2_8 = _RAND_40[511:0];
  _RAND_41 = {16{`RANDOM}};
  ram_2_9 = _RAND_41[511:0];
  _RAND_42 = {16{`RANDOM}};
  ram_2_10 = _RAND_42[511:0];
  _RAND_43 = {16{`RANDOM}};
  ram_2_11 = _RAND_43[511:0];
  _RAND_44 = {16{`RANDOM}};
  ram_2_12 = _RAND_44[511:0];
  _RAND_45 = {16{`RANDOM}};
  ram_2_13 = _RAND_45[511:0];
  _RAND_46 = {16{`RANDOM}};
  ram_2_14 = _RAND_46[511:0];
  _RAND_47 = {16{`RANDOM}};
  ram_2_15 = _RAND_47[511:0];
  _RAND_48 = {16{`RANDOM}};
  ram_3_0 = _RAND_48[511:0];
  _RAND_49 = {16{`RANDOM}};
  ram_3_1 = _RAND_49[511:0];
  _RAND_50 = {16{`RANDOM}};
  ram_3_2 = _RAND_50[511:0];
  _RAND_51 = {16{`RANDOM}};
  ram_3_3 = _RAND_51[511:0];
  _RAND_52 = {16{`RANDOM}};
  ram_3_4 = _RAND_52[511:0];
  _RAND_53 = {16{`RANDOM}};
  ram_3_5 = _RAND_53[511:0];
  _RAND_54 = {16{`RANDOM}};
  ram_3_6 = _RAND_54[511:0];
  _RAND_55 = {16{`RANDOM}};
  ram_3_7 = _RAND_55[511:0];
  _RAND_56 = {16{`RANDOM}};
  ram_3_8 = _RAND_56[511:0];
  _RAND_57 = {16{`RANDOM}};
  ram_3_9 = _RAND_57[511:0];
  _RAND_58 = {16{`RANDOM}};
  ram_3_10 = _RAND_58[511:0];
  _RAND_59 = {16{`RANDOM}};
  ram_3_11 = _RAND_59[511:0];
  _RAND_60 = {16{`RANDOM}};
  ram_3_12 = _RAND_60[511:0];
  _RAND_61 = {16{`RANDOM}};
  ram_3_13 = _RAND_61[511:0];
  _RAND_62 = {16{`RANDOM}};
  ram_3_14 = _RAND_62[511:0];
  _RAND_63 = {16{`RANDOM}};
  ram_3_15 = _RAND_63[511:0];
  _RAND_64 = {1{`RANDOM}};
  tag_0_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  tag_0_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  tag_0_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  tag_0_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  tag_0_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  tag_0_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  tag_0_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  tag_0_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  tag_0_8 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  tag_0_9 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  tag_0_10 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  tag_0_11 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  tag_0_12 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  tag_0_13 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  tag_0_14 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  tag_0_15 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  tag_1_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  tag_1_1 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  tag_1_2 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  tag_1_3 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  tag_1_4 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  tag_1_5 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  tag_1_6 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  tag_1_7 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  tag_1_8 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  tag_1_9 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  tag_1_10 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  tag_1_11 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  tag_1_12 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  tag_1_13 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  tag_1_14 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  tag_1_15 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  tag_2_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  tag_2_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  tag_2_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  tag_2_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  tag_2_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  tag_2_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  tag_2_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  tag_2_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  tag_2_8 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  tag_2_9 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  tag_2_10 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  tag_2_11 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  tag_2_12 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  tag_2_13 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  tag_2_14 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  tag_2_15 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  tag_3_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  tag_3_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  tag_3_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  tag_3_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  tag_3_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  tag_3_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  tag_3_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  tag_3_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  tag_3_8 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  tag_3_9 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  tag_3_10 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  tag_3_11 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  tag_3_12 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  tag_3_13 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  tag_3_14 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  tag_3_15 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_1_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_1_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_1_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_1_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_1_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_1_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_1_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_1_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_1_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_1_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_1_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_1_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_1_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_1_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_1_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_1_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_2_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_2_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_2_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_2_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_2_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_2_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_2_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_2_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_2_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_2_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_2_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_2_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_2_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_2_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_2_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_2_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_3_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_3_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_3_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_3_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_3_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_3_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_3_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_3_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_3_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_3_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_3_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_3_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_3_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_3_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_3_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_3_15 = _RAND_191[0:0];
  _RAND_192 = {2{`RANDOM}};
  receive_data_0 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  receive_data_1 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  receive_data_2 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  receive_data_3 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  receive_data_4 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  receive_data_5 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  receive_data_6 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  receive_data_7 = _RAND_199[63:0];
  _RAND_200 = {1{`RANDOM}};
  receive_num = _RAND_200[2:0];
  _RAND_201 = {1{`RANDOM}};
  quene_0 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  quene_1 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  quene_2 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  quene_3 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  quene_4 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  quene_5 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  quene_6 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  quene_7 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  quene_8 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  quene_9 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  quene_10 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  quene_11 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  quene_12 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  quene_13 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  quene_14 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  quene_15 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  state = _RAND_217[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [63:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_wready,
  output [31:0] io_to_axi_araddr,
  output [7:0]  io_to_axi_arlen,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output [7:0]  io_to_axi_awlen,
  output        io_to_axi_awvalid,
  output [63:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rlast,
  input         io_from_axi_rvalid,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [511:0] _RAND_2;
  reg [511:0] _RAND_3;
  reg [511:0] _RAND_4;
  reg [511:0] _RAND_5;
  reg [511:0] _RAND_6;
  reg [511:0] _RAND_7;
  reg [511:0] _RAND_8;
  reg [511:0] _RAND_9;
  reg [511:0] _RAND_10;
  reg [511:0] _RAND_11;
  reg [511:0] _RAND_12;
  reg [511:0] _RAND_13;
  reg [511:0] _RAND_14;
  reg [511:0] _RAND_15;
  reg [511:0] _RAND_16;
  reg [511:0] _RAND_17;
  reg [511:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [511:0] _RAND_21;
  reg [511:0] _RAND_22;
  reg [511:0] _RAND_23;
  reg [511:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [511:0] _RAND_26;
  reg [511:0] _RAND_27;
  reg [511:0] _RAND_28;
  reg [511:0] _RAND_29;
  reg [511:0] _RAND_30;
  reg [511:0] _RAND_31;
  reg [511:0] _RAND_32;
  reg [511:0] _RAND_33;
  reg [511:0] _RAND_34;
  reg [511:0] _RAND_35;
  reg [511:0] _RAND_36;
  reg [511:0] _RAND_37;
  reg [511:0] _RAND_38;
  reg [511:0] _RAND_39;
  reg [511:0] _RAND_40;
  reg [511:0] _RAND_41;
  reg [511:0] _RAND_42;
  reg [511:0] _RAND_43;
  reg [511:0] _RAND_44;
  reg [511:0] _RAND_45;
  reg [511:0] _RAND_46;
  reg [511:0] _RAND_47;
  reg [511:0] _RAND_48;
  reg [511:0] _RAND_49;
  reg [511:0] _RAND_50;
  reg [511:0] _RAND_51;
  reg [511:0] _RAND_52;
  reg [511:0] _RAND_53;
  reg [511:0] _RAND_54;
  reg [511:0] _RAND_55;
  reg [511:0] _RAND_56;
  reg [511:0] _RAND_57;
  reg [511:0] _RAND_58;
  reg [511:0] _RAND_59;
  reg [511:0] _RAND_60;
  reg [511:0] _RAND_61;
  reg [511:0] _RAND_62;
  reg [511:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [511:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [63:0] _RAND_258;
  reg [63:0] _RAND_259;
  reg [63:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [63:0] _RAND_263;
  reg [63:0] _RAND_264;
  reg [63:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] ram_0_0; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_1; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_2; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_3; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_4; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_5; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_6; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_7; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_8; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_9; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_10; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_11; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_12; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_13; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_14; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_15; // @[d_cache.scala 19:24]
  reg [511:0] ram_1_0; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_1; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_2; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_3; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_4; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_5; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_6; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_7; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_8; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_9; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_10; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_11; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_12; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_13; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_14; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_15; // @[d_cache.scala 20:24]
  reg [511:0] ram_2_0; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_1; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_2; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_3; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_4; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_5; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_6; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_7; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_8; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_9; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_10; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_11; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_12; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_13; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_14; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_15; // @[d_cache.scala 21:24]
  reg [511:0] ram_3_0; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_1; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_2; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_3; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_4; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_5; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_6; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_7; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_8; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_9; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_10; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_11; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_12; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_13; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_14; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_15; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_0; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 24:24]
  reg [31:0] tag_1_0; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_1; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_2; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_3; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_4; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_5; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_6; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_7; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_8; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_9; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_10; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_11; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_12; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_13; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_14; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_15; // @[d_cache.scala 25:24]
  reg [31:0] tag_2_0; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_1; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_2; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_3; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_4; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_5; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_6; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_7; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_8; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_9; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_10; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_11; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_12; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_13; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_14; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_15; // @[d_cache.scala 26:24]
  reg [31:0] tag_3_0; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_1; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_2; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_3; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_4; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_5; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_6; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_7; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_8; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_9; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_10; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_11; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_12; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_13; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_14; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_15; // @[d_cache.scala 27:24]
  reg  valid_0_0; // @[d_cache.scala 29:26]
  reg  valid_0_1; // @[d_cache.scala 29:26]
  reg  valid_0_2; // @[d_cache.scala 29:26]
  reg  valid_0_3; // @[d_cache.scala 29:26]
  reg  valid_0_4; // @[d_cache.scala 29:26]
  reg  valid_0_5; // @[d_cache.scala 29:26]
  reg  valid_0_6; // @[d_cache.scala 29:26]
  reg  valid_0_7; // @[d_cache.scala 29:26]
  reg  valid_0_8; // @[d_cache.scala 29:26]
  reg  valid_0_9; // @[d_cache.scala 29:26]
  reg  valid_0_10; // @[d_cache.scala 29:26]
  reg  valid_0_11; // @[d_cache.scala 29:26]
  reg  valid_0_12; // @[d_cache.scala 29:26]
  reg  valid_0_13; // @[d_cache.scala 29:26]
  reg  valid_0_14; // @[d_cache.scala 29:26]
  reg  valid_0_15; // @[d_cache.scala 29:26]
  reg  valid_1_0; // @[d_cache.scala 30:26]
  reg  valid_1_1; // @[d_cache.scala 30:26]
  reg  valid_1_2; // @[d_cache.scala 30:26]
  reg  valid_1_3; // @[d_cache.scala 30:26]
  reg  valid_1_4; // @[d_cache.scala 30:26]
  reg  valid_1_5; // @[d_cache.scala 30:26]
  reg  valid_1_6; // @[d_cache.scala 30:26]
  reg  valid_1_7; // @[d_cache.scala 30:26]
  reg  valid_1_8; // @[d_cache.scala 30:26]
  reg  valid_1_9; // @[d_cache.scala 30:26]
  reg  valid_1_10; // @[d_cache.scala 30:26]
  reg  valid_1_11; // @[d_cache.scala 30:26]
  reg  valid_1_12; // @[d_cache.scala 30:26]
  reg  valid_1_13; // @[d_cache.scala 30:26]
  reg  valid_1_14; // @[d_cache.scala 30:26]
  reg  valid_1_15; // @[d_cache.scala 30:26]
  reg  valid_2_0; // @[d_cache.scala 31:26]
  reg  valid_2_1; // @[d_cache.scala 31:26]
  reg  valid_2_2; // @[d_cache.scala 31:26]
  reg  valid_2_3; // @[d_cache.scala 31:26]
  reg  valid_2_4; // @[d_cache.scala 31:26]
  reg  valid_2_5; // @[d_cache.scala 31:26]
  reg  valid_2_6; // @[d_cache.scala 31:26]
  reg  valid_2_7; // @[d_cache.scala 31:26]
  reg  valid_2_8; // @[d_cache.scala 31:26]
  reg  valid_2_9; // @[d_cache.scala 31:26]
  reg  valid_2_10; // @[d_cache.scala 31:26]
  reg  valid_2_11; // @[d_cache.scala 31:26]
  reg  valid_2_12; // @[d_cache.scala 31:26]
  reg  valid_2_13; // @[d_cache.scala 31:26]
  reg  valid_2_14; // @[d_cache.scala 31:26]
  reg  valid_2_15; // @[d_cache.scala 31:26]
  reg  valid_3_0; // @[d_cache.scala 32:26]
  reg  valid_3_1; // @[d_cache.scala 32:26]
  reg  valid_3_2; // @[d_cache.scala 32:26]
  reg  valid_3_3; // @[d_cache.scala 32:26]
  reg  valid_3_4; // @[d_cache.scala 32:26]
  reg  valid_3_5; // @[d_cache.scala 32:26]
  reg  valid_3_6; // @[d_cache.scala 32:26]
  reg  valid_3_7; // @[d_cache.scala 32:26]
  reg  valid_3_8; // @[d_cache.scala 32:26]
  reg  valid_3_9; // @[d_cache.scala 32:26]
  reg  valid_3_10; // @[d_cache.scala 32:26]
  reg  valid_3_11; // @[d_cache.scala 32:26]
  reg  valid_3_12; // @[d_cache.scala 32:26]
  reg  valid_3_13; // @[d_cache.scala 32:26]
  reg  valid_3_14; // @[d_cache.scala 32:26]
  reg  valid_3_15; // @[d_cache.scala 32:26]
  reg  dirty_0_0; // @[d_cache.scala 34:26]
  reg  dirty_0_1; // @[d_cache.scala 34:26]
  reg  dirty_0_2; // @[d_cache.scala 34:26]
  reg  dirty_0_3; // @[d_cache.scala 34:26]
  reg  dirty_0_4; // @[d_cache.scala 34:26]
  reg  dirty_0_5; // @[d_cache.scala 34:26]
  reg  dirty_0_6; // @[d_cache.scala 34:26]
  reg  dirty_0_7; // @[d_cache.scala 34:26]
  reg  dirty_0_8; // @[d_cache.scala 34:26]
  reg  dirty_0_9; // @[d_cache.scala 34:26]
  reg  dirty_0_10; // @[d_cache.scala 34:26]
  reg  dirty_0_11; // @[d_cache.scala 34:26]
  reg  dirty_0_12; // @[d_cache.scala 34:26]
  reg  dirty_0_13; // @[d_cache.scala 34:26]
  reg  dirty_0_14; // @[d_cache.scala 34:26]
  reg  dirty_0_15; // @[d_cache.scala 34:26]
  reg  dirty_1_0; // @[d_cache.scala 35:26]
  reg  dirty_1_1; // @[d_cache.scala 35:26]
  reg  dirty_1_2; // @[d_cache.scala 35:26]
  reg  dirty_1_3; // @[d_cache.scala 35:26]
  reg  dirty_1_4; // @[d_cache.scala 35:26]
  reg  dirty_1_5; // @[d_cache.scala 35:26]
  reg  dirty_1_6; // @[d_cache.scala 35:26]
  reg  dirty_1_7; // @[d_cache.scala 35:26]
  reg  dirty_1_8; // @[d_cache.scala 35:26]
  reg  dirty_1_9; // @[d_cache.scala 35:26]
  reg  dirty_1_10; // @[d_cache.scala 35:26]
  reg  dirty_1_11; // @[d_cache.scala 35:26]
  reg  dirty_1_12; // @[d_cache.scala 35:26]
  reg  dirty_1_13; // @[d_cache.scala 35:26]
  reg  dirty_1_14; // @[d_cache.scala 35:26]
  reg  dirty_1_15; // @[d_cache.scala 35:26]
  reg  dirty_2_0; // @[d_cache.scala 36:26]
  reg  dirty_2_1; // @[d_cache.scala 36:26]
  reg  dirty_2_2; // @[d_cache.scala 36:26]
  reg  dirty_2_3; // @[d_cache.scala 36:26]
  reg  dirty_2_4; // @[d_cache.scala 36:26]
  reg  dirty_2_5; // @[d_cache.scala 36:26]
  reg  dirty_2_6; // @[d_cache.scala 36:26]
  reg  dirty_2_7; // @[d_cache.scala 36:26]
  reg  dirty_2_8; // @[d_cache.scala 36:26]
  reg  dirty_2_9; // @[d_cache.scala 36:26]
  reg  dirty_2_10; // @[d_cache.scala 36:26]
  reg  dirty_2_11; // @[d_cache.scala 36:26]
  reg  dirty_2_12; // @[d_cache.scala 36:26]
  reg  dirty_2_13; // @[d_cache.scala 36:26]
  reg  dirty_2_14; // @[d_cache.scala 36:26]
  reg  dirty_2_15; // @[d_cache.scala 36:26]
  reg  dirty_3_0; // @[d_cache.scala 37:26]
  reg  dirty_3_1; // @[d_cache.scala 37:26]
  reg  dirty_3_2; // @[d_cache.scala 37:26]
  reg  dirty_3_3; // @[d_cache.scala 37:26]
  reg  dirty_3_4; // @[d_cache.scala 37:26]
  reg  dirty_3_5; // @[d_cache.scala 37:26]
  reg  dirty_3_6; // @[d_cache.scala 37:26]
  reg  dirty_3_7; // @[d_cache.scala 37:26]
  reg  dirty_3_8; // @[d_cache.scala 37:26]
  reg  dirty_3_9; // @[d_cache.scala 37:26]
  reg  dirty_3_10; // @[d_cache.scala 37:26]
  reg  dirty_3_11; // @[d_cache.scala 37:26]
  reg  dirty_3_12; // @[d_cache.scala 37:26]
  reg  dirty_3_13; // @[d_cache.scala 37:26]
  reg  dirty_3_14; // @[d_cache.scala 37:26]
  reg  dirty_3_15; // @[d_cache.scala 37:26]
  reg [511:0] write_back_data; // @[d_cache.scala 44:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 45:34]
  reg [63:0] receive_data_0; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_1; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_2; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_3; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_4; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_5; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_6; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_7; // @[d_cache.scala 50:31]
  reg [2:0] receive_num; // @[d_cache.scala 51:30]
  reg [7:0] quene_0; // @[d_cache.scala 52:24]
  reg [7:0] quene_1; // @[d_cache.scala 52:24]
  reg [7:0] quene_2; // @[d_cache.scala 52:24]
  reg [7:0] quene_3; // @[d_cache.scala 52:24]
  reg [7:0] quene_4; // @[d_cache.scala 52:24]
  reg [7:0] quene_5; // @[d_cache.scala 52:24]
  reg [7:0] quene_6; // @[d_cache.scala 52:24]
  reg [7:0] quene_7; // @[d_cache.scala 52:24]
  reg [7:0] quene_8; // @[d_cache.scala 52:24]
  reg [7:0] quene_9; // @[d_cache.scala 52:24]
  reg [7:0] quene_10; // @[d_cache.scala 52:24]
  reg [7:0] quene_11; // @[d_cache.scala 52:24]
  reg [7:0] quene_12; // @[d_cache.scala 52:24]
  reg [7:0] quene_13; // @[d_cache.scala 52:24]
  reg [7:0] quene_14; // @[d_cache.scala 52:24]
  reg [7:0] quene_15; // @[d_cache.scala 52:24]
  wire [5:0] offset = io_from_lsu_araddr[5:0]; // @[d_cache.scala 54:36]
  wire [3:0] index = io_from_lsu_araddr[9:6]; // @[d_cache.scala 55:35]
  wire [21:0] tag = io_from_lsu_araddr[31:10]; // @[d_cache.scala 56:33]
  wire [8:0] shift_bit = {offset, 3'h0}; // @[d_cache.scala 58:28]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 71:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 70:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 69:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 68:20]
  wire [31:0] _GEN_1 = 4'h1 == index ? tag_0_1 : tag_0_0; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_2 = 4'h2 == index ? tag_0_2 : _GEN_1; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_3 = 4'h3 == index ? tag_0_3 : _GEN_2; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_4 = 4'h4 == index ? tag_0_4 : _GEN_3; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_5 = 4'h5 == index ? tag_0_5 : _GEN_4; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_6 = 4'h6 == index ? tag_0_6 : _GEN_5; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_7 = 4'h7 == index ? tag_0_7 : _GEN_6; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_8 = 4'h8 == index ? tag_0_8 : _GEN_7; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_9 = 4'h9 == index ? tag_0_9 : _GEN_8; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_10 = 4'ha == index ? tag_0_10 : _GEN_9; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_11 = 4'hb == index ? tag_0_11 : _GEN_10; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_12 = 4'hc == index ? tag_0_12 : _GEN_11; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_13 = 4'hd == index ? tag_0_13 : _GEN_12; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_14 = 4'he == index ? tag_0_14 : _GEN_13; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_15 = 4'hf == index ? tag_0_15 : _GEN_14; // @[d_cache.scala 73:{31,31}]
  wire [31:0] _GEN_5341 = {{10'd0}, tag}; // @[d_cache.scala 73:31]
  wire  _GEN_17 = 4'h1 == index ? valid_0_1 : valid_0_0; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_18 = 4'h2 == index ? valid_0_2 : _GEN_17; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_19 = 4'h3 == index ? valid_0_3 : _GEN_18; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_20 = 4'h4 == index ? valid_0_4 : _GEN_19; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_21 = 4'h5 == index ? valid_0_5 : _GEN_20; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_22 = 4'h6 == index ? valid_0_6 : _GEN_21; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_23 = 4'h7 == index ? valid_0_7 : _GEN_22; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_24 = 4'h8 == index ? valid_0_8 : _GEN_23; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_25 = 4'h9 == index ? valid_0_9 : _GEN_24; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_26 = 4'ha == index ? valid_0_10 : _GEN_25; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_27 = 4'hb == index ? valid_0_11 : _GEN_26; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_28 = 4'hc == index ? valid_0_12 : _GEN_27; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_29 = 4'hd == index ? valid_0_13 : _GEN_28; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_30 = 4'he == index ? valid_0_14 : _GEN_29; // @[d_cache.scala 73:{57,57}]
  wire  _GEN_31 = 4'hf == index ? valid_0_15 : _GEN_30; // @[d_cache.scala 73:{57,57}]
  wire  way0_hit = _GEN_15 == _GEN_5341 & _GEN_31; // @[d_cache.scala 73:40]
  wire [31:0] _GEN_33 = 4'h1 == index ? tag_1_1 : tag_1_0; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_34 = 4'h2 == index ? tag_1_2 : _GEN_33; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_35 = 4'h3 == index ? tag_1_3 : _GEN_34; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_36 = 4'h4 == index ? tag_1_4 : _GEN_35; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_37 = 4'h5 == index ? tag_1_5 : _GEN_36; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_38 = 4'h6 == index ? tag_1_6 : _GEN_37; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_39 = 4'h7 == index ? tag_1_7 : _GEN_38; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_40 = 4'h8 == index ? tag_1_8 : _GEN_39; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_41 = 4'h9 == index ? tag_1_9 : _GEN_40; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_42 = 4'ha == index ? tag_1_10 : _GEN_41; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_43 = 4'hb == index ? tag_1_11 : _GEN_42; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_44 = 4'hc == index ? tag_1_12 : _GEN_43; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_45 = 4'hd == index ? tag_1_13 : _GEN_44; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_46 = 4'he == index ? tag_1_14 : _GEN_45; // @[d_cache.scala 75:{31,31}]
  wire [31:0] _GEN_47 = 4'hf == index ? tag_1_15 : _GEN_46; // @[d_cache.scala 75:{31,31}]
  wire  _GEN_49 = 4'h1 == index ? valid_1_1 : valid_1_0; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_50 = 4'h2 == index ? valid_1_2 : _GEN_49; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_51 = 4'h3 == index ? valid_1_3 : _GEN_50; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_52 = 4'h4 == index ? valid_1_4 : _GEN_51; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_53 = 4'h5 == index ? valid_1_5 : _GEN_52; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_54 = 4'h6 == index ? valid_1_6 : _GEN_53; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_55 = 4'h7 == index ? valid_1_7 : _GEN_54; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_56 = 4'h8 == index ? valid_1_8 : _GEN_55; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_57 = 4'h9 == index ? valid_1_9 : _GEN_56; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_58 = 4'ha == index ? valid_1_10 : _GEN_57; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_59 = 4'hb == index ? valid_1_11 : _GEN_58; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_60 = 4'hc == index ? valid_1_12 : _GEN_59; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_61 = 4'hd == index ? valid_1_13 : _GEN_60; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_62 = 4'he == index ? valid_1_14 : _GEN_61; // @[d_cache.scala 75:{57,57}]
  wire  _GEN_63 = 4'hf == index ? valid_1_15 : _GEN_62; // @[d_cache.scala 75:{57,57}]
  wire  way1_hit = _GEN_47 == _GEN_5341 & _GEN_63; // @[d_cache.scala 75:40]
  wire [31:0] _GEN_65 = 4'h1 == index ? tag_2_1 : tag_2_0; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_66 = 4'h2 == index ? tag_2_2 : _GEN_65; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_67 = 4'h3 == index ? tag_2_3 : _GEN_66; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_68 = 4'h4 == index ? tag_2_4 : _GEN_67; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_69 = 4'h5 == index ? tag_2_5 : _GEN_68; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_70 = 4'h6 == index ? tag_2_6 : _GEN_69; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_71 = 4'h7 == index ? tag_2_7 : _GEN_70; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_72 = 4'h8 == index ? tag_2_8 : _GEN_71; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_73 = 4'h9 == index ? tag_2_9 : _GEN_72; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_74 = 4'ha == index ? tag_2_10 : _GEN_73; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_75 = 4'hb == index ? tag_2_11 : _GEN_74; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_76 = 4'hc == index ? tag_2_12 : _GEN_75; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_77 = 4'hd == index ? tag_2_13 : _GEN_76; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_78 = 4'he == index ? tag_2_14 : _GEN_77; // @[d_cache.scala 76:{31,31}]
  wire [31:0] _GEN_79 = 4'hf == index ? tag_2_15 : _GEN_78; // @[d_cache.scala 76:{31,31}]
  wire  _GEN_81 = 4'h1 == index ? valid_2_1 : valid_2_0; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_82 = 4'h2 == index ? valid_2_2 : _GEN_81; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_83 = 4'h3 == index ? valid_2_3 : _GEN_82; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_84 = 4'h4 == index ? valid_2_4 : _GEN_83; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_85 = 4'h5 == index ? valid_2_5 : _GEN_84; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_86 = 4'h6 == index ? valid_2_6 : _GEN_85; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_87 = 4'h7 == index ? valid_2_7 : _GEN_86; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_88 = 4'h8 == index ? valid_2_8 : _GEN_87; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_89 = 4'h9 == index ? valid_2_9 : _GEN_88; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_90 = 4'ha == index ? valid_2_10 : _GEN_89; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_91 = 4'hb == index ? valid_2_11 : _GEN_90; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_92 = 4'hc == index ? valid_2_12 : _GEN_91; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_93 = 4'hd == index ? valid_2_13 : _GEN_92; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_94 = 4'he == index ? valid_2_14 : _GEN_93; // @[d_cache.scala 76:{57,57}]
  wire  _GEN_95 = 4'hf == index ? valid_2_15 : _GEN_94; // @[d_cache.scala 76:{57,57}]
  wire  way2_hit = _GEN_79 == _GEN_5341 & _GEN_95; // @[d_cache.scala 76:40]
  wire [31:0] _GEN_97 = 4'h1 == index ? tag_3_1 : tag_3_0; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_98 = 4'h2 == index ? tag_3_2 : _GEN_97; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_99 = 4'h3 == index ? tag_3_3 : _GEN_98; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_100 = 4'h4 == index ? tag_3_4 : _GEN_99; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_101 = 4'h5 == index ? tag_3_5 : _GEN_100; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_102 = 4'h6 == index ? tag_3_6 : _GEN_101; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_103 = 4'h7 == index ? tag_3_7 : _GEN_102; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_104 = 4'h8 == index ? tag_3_8 : _GEN_103; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_105 = 4'h9 == index ? tag_3_9 : _GEN_104; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_106 = 4'ha == index ? tag_3_10 : _GEN_105; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_107 = 4'hb == index ? tag_3_11 : _GEN_106; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_108 = 4'hc == index ? tag_3_12 : _GEN_107; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_109 = 4'hd == index ? tag_3_13 : _GEN_108; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_110 = 4'he == index ? tag_3_14 : _GEN_109; // @[d_cache.scala 77:{31,31}]
  wire [31:0] _GEN_111 = 4'hf == index ? tag_3_15 : _GEN_110; // @[d_cache.scala 77:{31,31}]
  wire  _GEN_113 = 4'h1 == index ? valid_3_1 : valid_3_0; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_114 = 4'h2 == index ? valid_3_2 : _GEN_113; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_115 = 4'h3 == index ? valid_3_3 : _GEN_114; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_116 = 4'h4 == index ? valid_3_4 : _GEN_115; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_117 = 4'h5 == index ? valid_3_5 : _GEN_116; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_118 = 4'h6 == index ? valid_3_6 : _GEN_117; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_119 = 4'h7 == index ? valid_3_7 : _GEN_118; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_120 = 4'h8 == index ? valid_3_8 : _GEN_119; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_121 = 4'h9 == index ? valid_3_9 : _GEN_120; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_122 = 4'ha == index ? valid_3_10 : _GEN_121; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_123 = 4'hb == index ? valid_3_11 : _GEN_122; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_124 = 4'hc == index ? valid_3_12 : _GEN_123; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_125 = 4'hd == index ? valid_3_13 : _GEN_124; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_126 = 4'he == index ? valid_3_14 : _GEN_125; // @[d_cache.scala 77:{57,57}]
  wire  _GEN_127 = 4'hf == index ? valid_3_15 : _GEN_126; // @[d_cache.scala 77:{57,57}]
  wire  way3_hit = _GEN_111 == _GEN_5341 & _GEN_127; // @[d_cache.scala 77:40]
  wire [2:0] _unuse_way_T_4 = ~_GEN_127 ? 3'h4 : 3'h0; // @[d_cache.scala 80:108]
  wire [2:0] _unuse_way_T_5 = ~_GEN_95 ? 3'h3 : _unuse_way_T_4; // @[d_cache.scala 80:79]
  wire [2:0] _unuse_way_T_6 = ~_GEN_63 ? 3'h2 : _unuse_way_T_5; // @[d_cache.scala 80:50]
  wire [2:0] unuse_way = ~_GEN_31 ? 3'h1 : _unuse_way_T_6; // @[d_cache.scala 80:21]
  reg [3:0] state; // @[d_cache.scala 82:24]
  wire  _T_1 = io_from_lsu_araddr >= 32'ha0000000; // @[d_cache.scala 90:41]
  wire [3:0] _GEN_129 = _T_1 ? 4'h8 : 4'h2; // @[d_cache.scala 96:58 97:27 99:27]
  wire  _T_6 = way0_hit | way1_hit | way2_hit | way3_hit; // @[d_cache.scala 105:46]
  wire [63:0] _ram_0_T = io_from_lsu_wdata & wmask; // @[d_cache.scala 117:53]
  wire [574:0] _GEN_5704 = {{511'd0}, _ram_0_T}; // @[d_cache.scala 117:62]
  wire [574:0] _ram_0_T_1 = _GEN_5704 << shift_bit; // @[d_cache.scala 117:62]
  wire [574:0] _GEN_5705 = {{511'd0}, wmask}; // @[d_cache.scala 117:102]
  wire [574:0] _ram_0_T_2 = _GEN_5705 << shift_bit; // @[d_cache.scala 117:102]
  wire [574:0] _ram_0_T_3 = ~_ram_0_T_2; // @[d_cache.scala 117:94]
  wire [511:0] _GEN_136 = 4'h1 == index ? ram_0_1 : ram_0_0; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_137 = 4'h2 == index ? ram_0_2 : _GEN_136; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_138 = 4'h3 == index ? ram_0_3 : _GEN_137; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_139 = 4'h4 == index ? ram_0_4 : _GEN_138; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_140 = 4'h5 == index ? ram_0_5 : _GEN_139; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_141 = 4'h6 == index ? ram_0_6 : _GEN_140; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_142 = 4'h7 == index ? ram_0_7 : _GEN_141; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_143 = 4'h8 == index ? ram_0_8 : _GEN_142; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_144 = 4'h9 == index ? ram_0_9 : _GEN_143; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_145 = 4'ha == index ? ram_0_10 : _GEN_144; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_146 = 4'hb == index ? ram_0_11 : _GEN_145; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_147 = 4'hc == index ? ram_0_12 : _GEN_146; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_148 = 4'hd == index ? ram_0_13 : _GEN_147; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_149 = 4'he == index ? ram_0_14 : _GEN_148; // @[d_cache.scala 117:{92,92}]
  wire [511:0] _GEN_150 = 4'hf == index ? ram_0_15 : _GEN_149; // @[d_cache.scala 117:{92,92}]
  wire [574:0] _GEN_5350 = {{63'd0}, _GEN_150}; // @[d_cache.scala 117:92]
  wire [574:0] _ram_0_T_4 = _GEN_5350 & _ram_0_T_3; // @[d_cache.scala 117:92]
  wire [574:0] _ram_0_T_5 = _ram_0_T_1 | _ram_0_T_4; // @[d_cache.scala 117:76]
  wire [511:0] _GEN_151 = 4'h0 == index ? _ram_0_T_5[511:0] : ram_0_0; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_152 = 4'h1 == index ? _ram_0_T_5[511:0] : ram_0_1; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_153 = 4'h2 == index ? _ram_0_T_5[511:0] : ram_0_2; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_154 = 4'h3 == index ? _ram_0_T_5[511:0] : ram_0_3; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_155 = 4'h4 == index ? _ram_0_T_5[511:0] : ram_0_4; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_156 = 4'h5 == index ? _ram_0_T_5[511:0] : ram_0_5; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_157 = 4'h6 == index ? _ram_0_T_5[511:0] : ram_0_6; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_158 = 4'h7 == index ? _ram_0_T_5[511:0] : ram_0_7; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_159 = 4'h8 == index ? _ram_0_T_5[511:0] : ram_0_8; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_160 = 4'h9 == index ? _ram_0_T_5[511:0] : ram_0_9; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_161 = 4'ha == index ? _ram_0_T_5[511:0] : ram_0_10; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_162 = 4'hb == index ? _ram_0_T_5[511:0] : ram_0_11; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_163 = 4'hc == index ? _ram_0_T_5[511:0] : ram_0_12; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_164 = 4'hd == index ? _ram_0_T_5[511:0] : ram_0_13; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_165 = 4'he == index ? _ram_0_T_5[511:0] : ram_0_14; // @[d_cache.scala 117:{30,30} 19:24]
  wire [511:0] _GEN_166 = 4'hf == index ? _ram_0_T_5[511:0] : ram_0_15; // @[d_cache.scala 117:{30,30} 19:24]
  wire  _GEN_5351 = 4'h0 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_167 = 4'h0 == index | dirty_0_0; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5356 = 4'h1 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_168 = 4'h1 == index | dirty_0_1; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5357 = 4'h2 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_169 = 4'h2 == index | dirty_0_2; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5361 = 4'h3 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_170 = 4'h3 == index | dirty_0_3; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5365 = 4'h4 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_171 = 4'h4 == index | dirty_0_4; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5367 = 4'h5 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_172 = 4'h5 == index | dirty_0_5; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5369 = 4'h6 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_173 = 4'h6 == index | dirty_0_6; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5370 = 4'h7 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_174 = 4'h7 == index | dirty_0_7; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5374 = 4'h8 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_175 = 4'h8 == index | dirty_0_8; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5375 = 4'h9 == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_176 = 4'h9 == index | dirty_0_9; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5380 = 4'ha == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_177 = 4'ha == index | dirty_0_10; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5381 = 4'hb == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_178 = 4'hb == index | dirty_0_11; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5384 = 4'hc == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_179 = 4'hc == index | dirty_0_12; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5388 = 4'hd == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_180 = 4'hd == index | dirty_0_13; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5390 = 4'he == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_181 = 4'he == index | dirty_0_14; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_5392 = 4'hf == index; // @[d_cache.scala 118:{32,32} 34:26]
  wire  _GEN_182 = 4'hf == index | dirty_0_15; // @[d_cache.scala 118:{32,32} 34:26]
  wire [511:0] _GEN_184 = 4'h1 == index ? ram_1_1 : ram_1_0; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_185 = 4'h2 == index ? ram_1_2 : _GEN_184; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_186 = 4'h3 == index ? ram_1_3 : _GEN_185; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_187 = 4'h4 == index ? ram_1_4 : _GEN_186; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_188 = 4'h5 == index ? ram_1_5 : _GEN_187; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_189 = 4'h6 == index ? ram_1_6 : _GEN_188; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_190 = 4'h7 == index ? ram_1_7 : _GEN_189; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_191 = 4'h8 == index ? ram_1_8 : _GEN_190; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_192 = 4'h9 == index ? ram_1_9 : _GEN_191; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_193 = 4'ha == index ? ram_1_10 : _GEN_192; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_194 = 4'hb == index ? ram_1_11 : _GEN_193; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_195 = 4'hc == index ? ram_1_12 : _GEN_194; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_196 = 4'hd == index ? ram_1_13 : _GEN_195; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_197 = 4'he == index ? ram_1_14 : _GEN_196; // @[d_cache.scala 121:{92,92}]
  wire [511:0] _GEN_198 = 4'hf == index ? ram_1_15 : _GEN_197; // @[d_cache.scala 121:{92,92}]
  wire [574:0] _GEN_5393 = {{63'd0}, _GEN_198}; // @[d_cache.scala 121:92]
  wire [574:0] _ram_1_T_4 = _GEN_5393 & _ram_0_T_3; // @[d_cache.scala 121:92]
  wire [574:0] _ram_1_T_5 = _ram_0_T_1 | _ram_1_T_4; // @[d_cache.scala 121:76]
  wire [511:0] _GEN_199 = 4'h0 == index ? _ram_1_T_5[511:0] : ram_1_0; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_200 = 4'h1 == index ? _ram_1_T_5[511:0] : ram_1_1; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_201 = 4'h2 == index ? _ram_1_T_5[511:0] : ram_1_2; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_202 = 4'h3 == index ? _ram_1_T_5[511:0] : ram_1_3; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_203 = 4'h4 == index ? _ram_1_T_5[511:0] : ram_1_4; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_204 = 4'h5 == index ? _ram_1_T_5[511:0] : ram_1_5; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_205 = 4'h6 == index ? _ram_1_T_5[511:0] : ram_1_6; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_206 = 4'h7 == index ? _ram_1_T_5[511:0] : ram_1_7; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_207 = 4'h8 == index ? _ram_1_T_5[511:0] : ram_1_8; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_208 = 4'h9 == index ? _ram_1_T_5[511:0] : ram_1_9; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_209 = 4'ha == index ? _ram_1_T_5[511:0] : ram_1_10; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_210 = 4'hb == index ? _ram_1_T_5[511:0] : ram_1_11; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_211 = 4'hc == index ? _ram_1_T_5[511:0] : ram_1_12; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_212 = 4'hd == index ? _ram_1_T_5[511:0] : ram_1_13; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_213 = 4'he == index ? _ram_1_T_5[511:0] : ram_1_14; // @[d_cache.scala 121:{30,30} 20:24]
  wire [511:0] _GEN_214 = 4'hf == index ? _ram_1_T_5[511:0] : ram_1_15; // @[d_cache.scala 121:{30,30} 20:24]
  wire  _GEN_215 = _GEN_5351 | dirty_1_0; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_216 = _GEN_5356 | dirty_1_1; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_217 = _GEN_5357 | dirty_1_2; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_218 = _GEN_5361 | dirty_1_3; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_219 = _GEN_5365 | dirty_1_4; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_220 = _GEN_5367 | dirty_1_5; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_221 = _GEN_5369 | dirty_1_6; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_222 = _GEN_5370 | dirty_1_7; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_223 = _GEN_5374 | dirty_1_8; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_224 = _GEN_5375 | dirty_1_9; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_225 = _GEN_5380 | dirty_1_10; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_226 = _GEN_5381 | dirty_1_11; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_227 = _GEN_5384 | dirty_1_12; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_228 = _GEN_5388 | dirty_1_13; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_229 = _GEN_5390 | dirty_1_14; // @[d_cache.scala 122:{32,32} 35:26]
  wire  _GEN_230 = _GEN_5392 | dirty_1_15; // @[d_cache.scala 122:{32,32} 35:26]
  wire [511:0] _GEN_232 = 4'h1 == index ? ram_2_1 : ram_2_0; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_233 = 4'h2 == index ? ram_2_2 : _GEN_232; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_234 = 4'h3 == index ? ram_2_3 : _GEN_233; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_235 = 4'h4 == index ? ram_2_4 : _GEN_234; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_236 = 4'h5 == index ? ram_2_5 : _GEN_235; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_237 = 4'h6 == index ? ram_2_6 : _GEN_236; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_238 = 4'h7 == index ? ram_2_7 : _GEN_237; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_239 = 4'h8 == index ? ram_2_8 : _GEN_238; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_240 = 4'h9 == index ? ram_2_9 : _GEN_239; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_241 = 4'ha == index ? ram_2_10 : _GEN_240; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_242 = 4'hb == index ? ram_2_11 : _GEN_241; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_243 = 4'hc == index ? ram_2_12 : _GEN_242; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_244 = 4'hd == index ? ram_2_13 : _GEN_243; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_245 = 4'he == index ? ram_2_14 : _GEN_244; // @[d_cache.scala 125:{92,92}]
  wire [511:0] _GEN_246 = 4'hf == index ? ram_2_15 : _GEN_245; // @[d_cache.scala 125:{92,92}]
  wire [574:0] _GEN_5442 = {{63'd0}, _GEN_246}; // @[d_cache.scala 125:92]
  wire [574:0] _ram_2_T_4 = _GEN_5442 & _ram_0_T_3; // @[d_cache.scala 125:92]
  wire [574:0] _ram_2_T_5 = _ram_0_T_1 | _ram_2_T_4; // @[d_cache.scala 125:76]
  wire [511:0] _GEN_247 = 4'h0 == index ? _ram_2_T_5[511:0] : ram_2_0; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_248 = 4'h1 == index ? _ram_2_T_5[511:0] : ram_2_1; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_249 = 4'h2 == index ? _ram_2_T_5[511:0] : ram_2_2; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_250 = 4'h3 == index ? _ram_2_T_5[511:0] : ram_2_3; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_251 = 4'h4 == index ? _ram_2_T_5[511:0] : ram_2_4; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_252 = 4'h5 == index ? _ram_2_T_5[511:0] : ram_2_5; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_253 = 4'h6 == index ? _ram_2_T_5[511:0] : ram_2_6; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_254 = 4'h7 == index ? _ram_2_T_5[511:0] : ram_2_7; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_255 = 4'h8 == index ? _ram_2_T_5[511:0] : ram_2_8; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_256 = 4'h9 == index ? _ram_2_T_5[511:0] : ram_2_9; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_257 = 4'ha == index ? _ram_2_T_5[511:0] : ram_2_10; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_258 = 4'hb == index ? _ram_2_T_5[511:0] : ram_2_11; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_259 = 4'hc == index ? _ram_2_T_5[511:0] : ram_2_12; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_260 = 4'hd == index ? _ram_2_T_5[511:0] : ram_2_13; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_261 = 4'he == index ? _ram_2_T_5[511:0] : ram_2_14; // @[d_cache.scala 125:{30,30} 21:24]
  wire [511:0] _GEN_262 = 4'hf == index ? _ram_2_T_5[511:0] : ram_2_15; // @[d_cache.scala 125:{30,30} 21:24]
  wire  _GEN_263 = _GEN_5351 | dirty_2_0; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_264 = _GEN_5356 | dirty_2_1; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_265 = _GEN_5357 | dirty_2_2; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_266 = _GEN_5361 | dirty_2_3; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_267 = _GEN_5365 | dirty_2_4; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_268 = _GEN_5367 | dirty_2_5; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_269 = _GEN_5369 | dirty_2_6; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_270 = _GEN_5370 | dirty_2_7; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_271 = _GEN_5374 | dirty_2_8; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_272 = _GEN_5375 | dirty_2_9; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_273 = _GEN_5380 | dirty_2_10; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_274 = _GEN_5381 | dirty_2_11; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_275 = _GEN_5384 | dirty_2_12; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_276 = _GEN_5388 | dirty_2_13; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_277 = _GEN_5390 | dirty_2_14; // @[d_cache.scala 126:{32,32} 36:26]
  wire  _GEN_278 = _GEN_5392 | dirty_2_15; // @[d_cache.scala 126:{32,32} 36:26]
  wire [511:0] _GEN_280 = 4'h1 == index ? ram_3_1 : ram_3_0; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_281 = 4'h2 == index ? ram_3_2 : _GEN_280; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_282 = 4'h3 == index ? ram_3_3 : _GEN_281; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_283 = 4'h4 == index ? ram_3_4 : _GEN_282; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_284 = 4'h5 == index ? ram_3_5 : _GEN_283; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_285 = 4'h6 == index ? ram_3_6 : _GEN_284; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_286 = 4'h7 == index ? ram_3_7 : _GEN_285; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_287 = 4'h8 == index ? ram_3_8 : _GEN_286; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_288 = 4'h9 == index ? ram_3_9 : _GEN_287; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_289 = 4'ha == index ? ram_3_10 : _GEN_288; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_290 = 4'hb == index ? ram_3_11 : _GEN_289; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_291 = 4'hc == index ? ram_3_12 : _GEN_290; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_292 = 4'hd == index ? ram_3_13 : _GEN_291; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_293 = 4'he == index ? ram_3_14 : _GEN_292; // @[d_cache.scala 129:{92,92}]
  wire [511:0] _GEN_294 = 4'hf == index ? ram_3_15 : _GEN_293; // @[d_cache.scala 129:{92,92}]
  wire [574:0] _GEN_5480 = {{63'd0}, _GEN_294}; // @[d_cache.scala 129:92]
  wire [574:0] _ram_3_T_4 = _GEN_5480 & _ram_0_T_3; // @[d_cache.scala 129:92]
  wire [574:0] _ram_3_T_5 = _ram_0_T_1 | _ram_3_T_4; // @[d_cache.scala 129:76]
  wire [511:0] _GEN_295 = 4'h0 == index ? _ram_3_T_5[511:0] : ram_3_0; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_296 = 4'h1 == index ? _ram_3_T_5[511:0] : ram_3_1; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_297 = 4'h2 == index ? _ram_3_T_5[511:0] : ram_3_2; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_298 = 4'h3 == index ? _ram_3_T_5[511:0] : ram_3_3; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_299 = 4'h4 == index ? _ram_3_T_5[511:0] : ram_3_4; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_300 = 4'h5 == index ? _ram_3_T_5[511:0] : ram_3_5; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_301 = 4'h6 == index ? _ram_3_T_5[511:0] : ram_3_6; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_302 = 4'h7 == index ? _ram_3_T_5[511:0] : ram_3_7; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_303 = 4'h8 == index ? _ram_3_T_5[511:0] : ram_3_8; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_304 = 4'h9 == index ? _ram_3_T_5[511:0] : ram_3_9; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_305 = 4'ha == index ? _ram_3_T_5[511:0] : ram_3_10; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_306 = 4'hb == index ? _ram_3_T_5[511:0] : ram_3_11; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_307 = 4'hc == index ? _ram_3_T_5[511:0] : ram_3_12; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_308 = 4'hd == index ? _ram_3_T_5[511:0] : ram_3_13; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_309 = 4'he == index ? _ram_3_T_5[511:0] : ram_3_14; // @[d_cache.scala 129:{30,30} 22:24]
  wire [511:0] _GEN_310 = 4'hf == index ? _ram_3_T_5[511:0] : ram_3_15; // @[d_cache.scala 129:{30,30} 22:24]
  wire  _GEN_311 = _GEN_5351 | dirty_3_0; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_312 = _GEN_5356 | dirty_3_1; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_313 = _GEN_5357 | dirty_3_2; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_314 = _GEN_5361 | dirty_3_3; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_315 = _GEN_5365 | dirty_3_4; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_316 = _GEN_5367 | dirty_3_5; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_317 = _GEN_5369 | dirty_3_6; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_318 = _GEN_5370 | dirty_3_7; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_319 = _GEN_5374 | dirty_3_8; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_320 = _GEN_5375 | dirty_3_9; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_321 = _GEN_5380 | dirty_3_10; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_322 = _GEN_5381 | dirty_3_11; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_323 = _GEN_5384 | dirty_3_12; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_324 = _GEN_5388 | dirty_3_13; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_325 = _GEN_5390 | dirty_3_14; // @[d_cache.scala 130:{32,32} 37:26]
  wire  _GEN_326 = _GEN_5392 | dirty_3_15; // @[d_cache.scala 130:{32,32} 37:26]
  wire [3:0] _GEN_327 = way3_hit ? 4'h0 : 4'h4; // @[d_cache.scala 127:33 128:23 132:23]
  wire [511:0] _GEN_328 = way3_hit ? _GEN_295 : ram_3_0; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_329 = way3_hit ? _GEN_296 : ram_3_1; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_330 = way3_hit ? _GEN_297 : ram_3_2; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_331 = way3_hit ? _GEN_298 : ram_3_3; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_332 = way3_hit ? _GEN_299 : ram_3_4; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_333 = way3_hit ? _GEN_300 : ram_3_5; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_334 = way3_hit ? _GEN_301 : ram_3_6; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_335 = way3_hit ? _GEN_302 : ram_3_7; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_336 = way3_hit ? _GEN_303 : ram_3_8; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_337 = way3_hit ? _GEN_304 : ram_3_9; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_338 = way3_hit ? _GEN_305 : ram_3_10; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_339 = way3_hit ? _GEN_306 : ram_3_11; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_340 = way3_hit ? _GEN_307 : ram_3_12; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_341 = way3_hit ? _GEN_308 : ram_3_13; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_342 = way3_hit ? _GEN_309 : ram_3_14; // @[d_cache.scala 127:33 22:24]
  wire [511:0] _GEN_343 = way3_hit ? _GEN_310 : ram_3_15; // @[d_cache.scala 127:33 22:24]
  wire  _GEN_344 = way3_hit ? _GEN_311 : dirty_3_0; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_345 = way3_hit ? _GEN_312 : dirty_3_1; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_346 = way3_hit ? _GEN_313 : dirty_3_2; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_347 = way3_hit ? _GEN_314 : dirty_3_3; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_348 = way3_hit ? _GEN_315 : dirty_3_4; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_349 = way3_hit ? _GEN_316 : dirty_3_5; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_350 = way3_hit ? _GEN_317 : dirty_3_6; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_351 = way3_hit ? _GEN_318 : dirty_3_7; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_352 = way3_hit ? _GEN_319 : dirty_3_8; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_353 = way3_hit ? _GEN_320 : dirty_3_9; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_354 = way3_hit ? _GEN_321 : dirty_3_10; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_355 = way3_hit ? _GEN_322 : dirty_3_11; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_356 = way3_hit ? _GEN_323 : dirty_3_12; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_357 = way3_hit ? _GEN_324 : dirty_3_13; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_358 = way3_hit ? _GEN_325 : dirty_3_14; // @[d_cache.scala 127:33 37:26]
  wire  _GEN_359 = way3_hit ? _GEN_326 : dirty_3_15; // @[d_cache.scala 127:33 37:26]
  wire [3:0] _GEN_360 = way2_hit ? 4'h0 : _GEN_327; // @[d_cache.scala 123:33 124:23]
  wire [511:0] _GEN_361 = way2_hit ? _GEN_247 : ram_2_0; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_362 = way2_hit ? _GEN_248 : ram_2_1; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_363 = way2_hit ? _GEN_249 : ram_2_2; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_364 = way2_hit ? _GEN_250 : ram_2_3; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_365 = way2_hit ? _GEN_251 : ram_2_4; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_366 = way2_hit ? _GEN_252 : ram_2_5; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_367 = way2_hit ? _GEN_253 : ram_2_6; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_368 = way2_hit ? _GEN_254 : ram_2_7; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_369 = way2_hit ? _GEN_255 : ram_2_8; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_370 = way2_hit ? _GEN_256 : ram_2_9; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_371 = way2_hit ? _GEN_257 : ram_2_10; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_372 = way2_hit ? _GEN_258 : ram_2_11; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_373 = way2_hit ? _GEN_259 : ram_2_12; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_374 = way2_hit ? _GEN_260 : ram_2_13; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_375 = way2_hit ? _GEN_261 : ram_2_14; // @[d_cache.scala 123:33 21:24]
  wire [511:0] _GEN_376 = way2_hit ? _GEN_262 : ram_2_15; // @[d_cache.scala 123:33 21:24]
  wire  _GEN_377 = way2_hit ? _GEN_263 : dirty_2_0; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_378 = way2_hit ? _GEN_264 : dirty_2_1; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_379 = way2_hit ? _GEN_265 : dirty_2_2; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_380 = way2_hit ? _GEN_266 : dirty_2_3; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_381 = way2_hit ? _GEN_267 : dirty_2_4; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_382 = way2_hit ? _GEN_268 : dirty_2_5; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_383 = way2_hit ? _GEN_269 : dirty_2_6; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_384 = way2_hit ? _GEN_270 : dirty_2_7; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_385 = way2_hit ? _GEN_271 : dirty_2_8; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_386 = way2_hit ? _GEN_272 : dirty_2_9; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_387 = way2_hit ? _GEN_273 : dirty_2_10; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_388 = way2_hit ? _GEN_274 : dirty_2_11; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_389 = way2_hit ? _GEN_275 : dirty_2_12; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_390 = way2_hit ? _GEN_276 : dirty_2_13; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_391 = way2_hit ? _GEN_277 : dirty_2_14; // @[d_cache.scala 123:33 36:26]
  wire  _GEN_392 = way2_hit ? _GEN_278 : dirty_2_15; // @[d_cache.scala 123:33 36:26]
  wire [511:0] _GEN_393 = way2_hit ? ram_3_0 : _GEN_328; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_394 = way2_hit ? ram_3_1 : _GEN_329; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_395 = way2_hit ? ram_3_2 : _GEN_330; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_396 = way2_hit ? ram_3_3 : _GEN_331; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_397 = way2_hit ? ram_3_4 : _GEN_332; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_398 = way2_hit ? ram_3_5 : _GEN_333; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_399 = way2_hit ? ram_3_6 : _GEN_334; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_400 = way2_hit ? ram_3_7 : _GEN_335; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_401 = way2_hit ? ram_3_8 : _GEN_336; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_402 = way2_hit ? ram_3_9 : _GEN_337; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_403 = way2_hit ? ram_3_10 : _GEN_338; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_404 = way2_hit ? ram_3_11 : _GEN_339; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_405 = way2_hit ? ram_3_12 : _GEN_340; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_406 = way2_hit ? ram_3_13 : _GEN_341; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_407 = way2_hit ? ram_3_14 : _GEN_342; // @[d_cache.scala 123:33 22:24]
  wire [511:0] _GEN_408 = way2_hit ? ram_3_15 : _GEN_343; // @[d_cache.scala 123:33 22:24]
  wire  _GEN_409 = way2_hit ? dirty_3_0 : _GEN_344; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_410 = way2_hit ? dirty_3_1 : _GEN_345; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_411 = way2_hit ? dirty_3_2 : _GEN_346; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_412 = way2_hit ? dirty_3_3 : _GEN_347; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_413 = way2_hit ? dirty_3_4 : _GEN_348; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_414 = way2_hit ? dirty_3_5 : _GEN_349; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_415 = way2_hit ? dirty_3_6 : _GEN_350; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_416 = way2_hit ? dirty_3_7 : _GEN_351; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_417 = way2_hit ? dirty_3_8 : _GEN_352; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_418 = way2_hit ? dirty_3_9 : _GEN_353; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_419 = way2_hit ? dirty_3_10 : _GEN_354; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_420 = way2_hit ? dirty_3_11 : _GEN_355; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_421 = way2_hit ? dirty_3_12 : _GEN_356; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_422 = way2_hit ? dirty_3_13 : _GEN_357; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_423 = way2_hit ? dirty_3_14 : _GEN_358; // @[d_cache.scala 123:33 37:26]
  wire  _GEN_424 = way2_hit ? dirty_3_15 : _GEN_359; // @[d_cache.scala 123:33 37:26]
  wire [3:0] _GEN_425 = way1_hit ? 4'h0 : _GEN_360; // @[d_cache.scala 119:33 120:23]
  wire [511:0] _GEN_426 = way1_hit ? _GEN_199 : ram_1_0; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_427 = way1_hit ? _GEN_200 : ram_1_1; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_428 = way1_hit ? _GEN_201 : ram_1_2; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_429 = way1_hit ? _GEN_202 : ram_1_3; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_430 = way1_hit ? _GEN_203 : ram_1_4; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_431 = way1_hit ? _GEN_204 : ram_1_5; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_432 = way1_hit ? _GEN_205 : ram_1_6; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_433 = way1_hit ? _GEN_206 : ram_1_7; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_434 = way1_hit ? _GEN_207 : ram_1_8; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_435 = way1_hit ? _GEN_208 : ram_1_9; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_436 = way1_hit ? _GEN_209 : ram_1_10; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_437 = way1_hit ? _GEN_210 : ram_1_11; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_438 = way1_hit ? _GEN_211 : ram_1_12; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_439 = way1_hit ? _GEN_212 : ram_1_13; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_440 = way1_hit ? _GEN_213 : ram_1_14; // @[d_cache.scala 119:33 20:24]
  wire [511:0] _GEN_441 = way1_hit ? _GEN_214 : ram_1_15; // @[d_cache.scala 119:33 20:24]
  wire  _GEN_442 = way1_hit ? _GEN_215 : dirty_1_0; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_443 = way1_hit ? _GEN_216 : dirty_1_1; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_444 = way1_hit ? _GEN_217 : dirty_1_2; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_445 = way1_hit ? _GEN_218 : dirty_1_3; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_446 = way1_hit ? _GEN_219 : dirty_1_4; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_447 = way1_hit ? _GEN_220 : dirty_1_5; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_448 = way1_hit ? _GEN_221 : dirty_1_6; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_449 = way1_hit ? _GEN_222 : dirty_1_7; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_450 = way1_hit ? _GEN_223 : dirty_1_8; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_451 = way1_hit ? _GEN_224 : dirty_1_9; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_452 = way1_hit ? _GEN_225 : dirty_1_10; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_453 = way1_hit ? _GEN_226 : dirty_1_11; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_454 = way1_hit ? _GEN_227 : dirty_1_12; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_455 = way1_hit ? _GEN_228 : dirty_1_13; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_456 = way1_hit ? _GEN_229 : dirty_1_14; // @[d_cache.scala 119:33 35:26]
  wire  _GEN_457 = way1_hit ? _GEN_230 : dirty_1_15; // @[d_cache.scala 119:33 35:26]
  wire [511:0] _GEN_458 = way1_hit ? ram_2_0 : _GEN_361; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_459 = way1_hit ? ram_2_1 : _GEN_362; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_460 = way1_hit ? ram_2_2 : _GEN_363; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_461 = way1_hit ? ram_2_3 : _GEN_364; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_462 = way1_hit ? ram_2_4 : _GEN_365; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_463 = way1_hit ? ram_2_5 : _GEN_366; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_464 = way1_hit ? ram_2_6 : _GEN_367; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_465 = way1_hit ? ram_2_7 : _GEN_368; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_466 = way1_hit ? ram_2_8 : _GEN_369; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_467 = way1_hit ? ram_2_9 : _GEN_370; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_468 = way1_hit ? ram_2_10 : _GEN_371; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_469 = way1_hit ? ram_2_11 : _GEN_372; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_470 = way1_hit ? ram_2_12 : _GEN_373; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_471 = way1_hit ? ram_2_13 : _GEN_374; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_472 = way1_hit ? ram_2_14 : _GEN_375; // @[d_cache.scala 119:33 21:24]
  wire [511:0] _GEN_473 = way1_hit ? ram_2_15 : _GEN_376; // @[d_cache.scala 119:33 21:24]
  wire  _GEN_474 = way1_hit ? dirty_2_0 : _GEN_377; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_475 = way1_hit ? dirty_2_1 : _GEN_378; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_476 = way1_hit ? dirty_2_2 : _GEN_379; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_477 = way1_hit ? dirty_2_3 : _GEN_380; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_478 = way1_hit ? dirty_2_4 : _GEN_381; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_479 = way1_hit ? dirty_2_5 : _GEN_382; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_480 = way1_hit ? dirty_2_6 : _GEN_383; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_481 = way1_hit ? dirty_2_7 : _GEN_384; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_482 = way1_hit ? dirty_2_8 : _GEN_385; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_483 = way1_hit ? dirty_2_9 : _GEN_386; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_484 = way1_hit ? dirty_2_10 : _GEN_387; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_485 = way1_hit ? dirty_2_11 : _GEN_388; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_486 = way1_hit ? dirty_2_12 : _GEN_389; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_487 = way1_hit ? dirty_2_13 : _GEN_390; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_488 = way1_hit ? dirty_2_14 : _GEN_391; // @[d_cache.scala 119:33 36:26]
  wire  _GEN_489 = way1_hit ? dirty_2_15 : _GEN_392; // @[d_cache.scala 119:33 36:26]
  wire [511:0] _GEN_490 = way1_hit ? ram_3_0 : _GEN_393; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_491 = way1_hit ? ram_3_1 : _GEN_394; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_492 = way1_hit ? ram_3_2 : _GEN_395; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_493 = way1_hit ? ram_3_3 : _GEN_396; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_494 = way1_hit ? ram_3_4 : _GEN_397; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_495 = way1_hit ? ram_3_5 : _GEN_398; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_496 = way1_hit ? ram_3_6 : _GEN_399; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_497 = way1_hit ? ram_3_7 : _GEN_400; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_498 = way1_hit ? ram_3_8 : _GEN_401; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_499 = way1_hit ? ram_3_9 : _GEN_402; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_500 = way1_hit ? ram_3_10 : _GEN_403; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_501 = way1_hit ? ram_3_11 : _GEN_404; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_502 = way1_hit ? ram_3_12 : _GEN_405; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_503 = way1_hit ? ram_3_13 : _GEN_406; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_504 = way1_hit ? ram_3_14 : _GEN_407; // @[d_cache.scala 119:33 22:24]
  wire [511:0] _GEN_505 = way1_hit ? ram_3_15 : _GEN_408; // @[d_cache.scala 119:33 22:24]
  wire  _GEN_506 = way1_hit ? dirty_3_0 : _GEN_409; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_507 = way1_hit ? dirty_3_1 : _GEN_410; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_508 = way1_hit ? dirty_3_2 : _GEN_411; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_509 = way1_hit ? dirty_3_3 : _GEN_412; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_510 = way1_hit ? dirty_3_4 : _GEN_413; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_511 = way1_hit ? dirty_3_5 : _GEN_414; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_512 = way1_hit ? dirty_3_6 : _GEN_415; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_513 = way1_hit ? dirty_3_7 : _GEN_416; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_514 = way1_hit ? dirty_3_8 : _GEN_417; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_515 = way1_hit ? dirty_3_9 : _GEN_418; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_516 = way1_hit ? dirty_3_10 : _GEN_419; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_517 = way1_hit ? dirty_3_11 : _GEN_420; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_518 = way1_hit ? dirty_3_12 : _GEN_421; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_519 = way1_hit ? dirty_3_13 : _GEN_422; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_520 = way1_hit ? dirty_3_14 : _GEN_423; // @[d_cache.scala 119:33 37:26]
  wire  _GEN_521 = way1_hit ? dirty_3_15 : _GEN_424; // @[d_cache.scala 119:33 37:26]
  wire [3:0] _GEN_522 = way0_hit ? 4'h0 : _GEN_425; // @[d_cache.scala 115:27 116:23]
  wire [511:0] _GEN_523 = way0_hit ? _GEN_151 : ram_0_0; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_524 = way0_hit ? _GEN_152 : ram_0_1; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_525 = way0_hit ? _GEN_153 : ram_0_2; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_526 = way0_hit ? _GEN_154 : ram_0_3; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_527 = way0_hit ? _GEN_155 : ram_0_4; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_528 = way0_hit ? _GEN_156 : ram_0_5; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_529 = way0_hit ? _GEN_157 : ram_0_6; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_530 = way0_hit ? _GEN_158 : ram_0_7; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_531 = way0_hit ? _GEN_159 : ram_0_8; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_532 = way0_hit ? _GEN_160 : ram_0_9; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_533 = way0_hit ? _GEN_161 : ram_0_10; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_534 = way0_hit ? _GEN_162 : ram_0_11; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_535 = way0_hit ? _GEN_163 : ram_0_12; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_536 = way0_hit ? _GEN_164 : ram_0_13; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_537 = way0_hit ? _GEN_165 : ram_0_14; // @[d_cache.scala 115:27 19:24]
  wire [511:0] _GEN_538 = way0_hit ? _GEN_166 : ram_0_15; // @[d_cache.scala 115:27 19:24]
  wire  _GEN_539 = way0_hit ? _GEN_167 : dirty_0_0; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_540 = way0_hit ? _GEN_168 : dirty_0_1; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_541 = way0_hit ? _GEN_169 : dirty_0_2; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_542 = way0_hit ? _GEN_170 : dirty_0_3; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_543 = way0_hit ? _GEN_171 : dirty_0_4; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_544 = way0_hit ? _GEN_172 : dirty_0_5; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_545 = way0_hit ? _GEN_173 : dirty_0_6; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_546 = way0_hit ? _GEN_174 : dirty_0_7; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_547 = way0_hit ? _GEN_175 : dirty_0_8; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_548 = way0_hit ? _GEN_176 : dirty_0_9; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_549 = way0_hit ? _GEN_177 : dirty_0_10; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_550 = way0_hit ? _GEN_178 : dirty_0_11; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_551 = way0_hit ? _GEN_179 : dirty_0_12; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_552 = way0_hit ? _GEN_180 : dirty_0_13; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_553 = way0_hit ? _GEN_181 : dirty_0_14; // @[d_cache.scala 115:27 34:26]
  wire  _GEN_554 = way0_hit ? _GEN_182 : dirty_0_15; // @[d_cache.scala 115:27 34:26]
  wire [511:0] _GEN_555 = way0_hit ? ram_1_0 : _GEN_426; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_556 = way0_hit ? ram_1_1 : _GEN_427; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_557 = way0_hit ? ram_1_2 : _GEN_428; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_558 = way0_hit ? ram_1_3 : _GEN_429; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_559 = way0_hit ? ram_1_4 : _GEN_430; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_560 = way0_hit ? ram_1_5 : _GEN_431; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_561 = way0_hit ? ram_1_6 : _GEN_432; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_562 = way0_hit ? ram_1_7 : _GEN_433; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_563 = way0_hit ? ram_1_8 : _GEN_434; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_564 = way0_hit ? ram_1_9 : _GEN_435; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_565 = way0_hit ? ram_1_10 : _GEN_436; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_566 = way0_hit ? ram_1_11 : _GEN_437; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_567 = way0_hit ? ram_1_12 : _GEN_438; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_568 = way0_hit ? ram_1_13 : _GEN_439; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_569 = way0_hit ? ram_1_14 : _GEN_440; // @[d_cache.scala 115:27 20:24]
  wire [511:0] _GEN_570 = way0_hit ? ram_1_15 : _GEN_441; // @[d_cache.scala 115:27 20:24]
  wire  _GEN_571 = way0_hit ? dirty_1_0 : _GEN_442; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_572 = way0_hit ? dirty_1_1 : _GEN_443; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_573 = way0_hit ? dirty_1_2 : _GEN_444; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_574 = way0_hit ? dirty_1_3 : _GEN_445; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_575 = way0_hit ? dirty_1_4 : _GEN_446; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_576 = way0_hit ? dirty_1_5 : _GEN_447; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_577 = way0_hit ? dirty_1_6 : _GEN_448; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_578 = way0_hit ? dirty_1_7 : _GEN_449; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_579 = way0_hit ? dirty_1_8 : _GEN_450; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_580 = way0_hit ? dirty_1_9 : _GEN_451; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_581 = way0_hit ? dirty_1_10 : _GEN_452; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_582 = way0_hit ? dirty_1_11 : _GEN_453; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_583 = way0_hit ? dirty_1_12 : _GEN_454; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_584 = way0_hit ? dirty_1_13 : _GEN_455; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_585 = way0_hit ? dirty_1_14 : _GEN_456; // @[d_cache.scala 115:27 35:26]
  wire  _GEN_586 = way0_hit ? dirty_1_15 : _GEN_457; // @[d_cache.scala 115:27 35:26]
  wire [511:0] _GEN_587 = way0_hit ? ram_2_0 : _GEN_458; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_588 = way0_hit ? ram_2_1 : _GEN_459; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_589 = way0_hit ? ram_2_2 : _GEN_460; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_590 = way0_hit ? ram_2_3 : _GEN_461; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_591 = way0_hit ? ram_2_4 : _GEN_462; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_592 = way0_hit ? ram_2_5 : _GEN_463; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_593 = way0_hit ? ram_2_6 : _GEN_464; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_594 = way0_hit ? ram_2_7 : _GEN_465; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_595 = way0_hit ? ram_2_8 : _GEN_466; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_596 = way0_hit ? ram_2_9 : _GEN_467; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_597 = way0_hit ? ram_2_10 : _GEN_468; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_598 = way0_hit ? ram_2_11 : _GEN_469; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_599 = way0_hit ? ram_2_12 : _GEN_470; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_600 = way0_hit ? ram_2_13 : _GEN_471; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_601 = way0_hit ? ram_2_14 : _GEN_472; // @[d_cache.scala 115:27 21:24]
  wire [511:0] _GEN_602 = way0_hit ? ram_2_15 : _GEN_473; // @[d_cache.scala 115:27 21:24]
  wire  _GEN_603 = way0_hit ? dirty_2_0 : _GEN_474; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_604 = way0_hit ? dirty_2_1 : _GEN_475; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_605 = way0_hit ? dirty_2_2 : _GEN_476; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_606 = way0_hit ? dirty_2_3 : _GEN_477; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_607 = way0_hit ? dirty_2_4 : _GEN_478; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_608 = way0_hit ? dirty_2_5 : _GEN_479; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_609 = way0_hit ? dirty_2_6 : _GEN_480; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_610 = way0_hit ? dirty_2_7 : _GEN_481; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_611 = way0_hit ? dirty_2_8 : _GEN_482; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_612 = way0_hit ? dirty_2_9 : _GEN_483; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_613 = way0_hit ? dirty_2_10 : _GEN_484; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_614 = way0_hit ? dirty_2_11 : _GEN_485; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_615 = way0_hit ? dirty_2_12 : _GEN_486; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_616 = way0_hit ? dirty_2_13 : _GEN_487; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_617 = way0_hit ? dirty_2_14 : _GEN_488; // @[d_cache.scala 115:27 36:26]
  wire  _GEN_618 = way0_hit ? dirty_2_15 : _GEN_489; // @[d_cache.scala 115:27 36:26]
  wire [511:0] _GEN_619 = way0_hit ? ram_3_0 : _GEN_490; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_620 = way0_hit ? ram_3_1 : _GEN_491; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_621 = way0_hit ? ram_3_2 : _GEN_492; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_622 = way0_hit ? ram_3_3 : _GEN_493; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_623 = way0_hit ? ram_3_4 : _GEN_494; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_624 = way0_hit ? ram_3_5 : _GEN_495; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_625 = way0_hit ? ram_3_6 : _GEN_496; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_626 = way0_hit ? ram_3_7 : _GEN_497; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_627 = way0_hit ? ram_3_8 : _GEN_498; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_628 = way0_hit ? ram_3_9 : _GEN_499; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_629 = way0_hit ? ram_3_10 : _GEN_500; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_630 = way0_hit ? ram_3_11 : _GEN_501; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_631 = way0_hit ? ram_3_12 : _GEN_502; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_632 = way0_hit ? ram_3_13 : _GEN_503; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_633 = way0_hit ? ram_3_14 : _GEN_504; // @[d_cache.scala 115:27 22:24]
  wire [511:0] _GEN_634 = way0_hit ? ram_3_15 : _GEN_505; // @[d_cache.scala 115:27 22:24]
  wire  _GEN_635 = way0_hit ? dirty_3_0 : _GEN_506; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_636 = way0_hit ? dirty_3_1 : _GEN_507; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_637 = way0_hit ? dirty_3_2 : _GEN_508; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_638 = way0_hit ? dirty_3_3 : _GEN_509; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_639 = way0_hit ? dirty_3_4 : _GEN_510; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_640 = way0_hit ? dirty_3_5 : _GEN_511; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_641 = way0_hit ? dirty_3_6 : _GEN_512; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_642 = way0_hit ? dirty_3_7 : _GEN_513; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_643 = way0_hit ? dirty_3_8 : _GEN_514; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_644 = way0_hit ? dirty_3_9 : _GEN_515; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_645 = way0_hit ? dirty_3_10 : _GEN_516; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_646 = way0_hit ? dirty_3_11 : _GEN_517; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_647 = way0_hit ? dirty_3_12 : _GEN_518; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_648 = way0_hit ? dirty_3_13 : _GEN_519; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_649 = way0_hit ? dirty_3_14 : _GEN_520; // @[d_cache.scala 115:27 37:26]
  wire  _GEN_650 = way0_hit ? dirty_3_15 : _GEN_521; // @[d_cache.scala 115:27 37:26]
  wire [63:0] _GEN_651 = 3'h0 == receive_num ? io_from_axi_rdata : receive_data_0; // @[d_cache.scala 137:{43,43} 50:31]
  wire [63:0] _GEN_652 = 3'h1 == receive_num ? io_from_axi_rdata : receive_data_1; // @[d_cache.scala 137:{43,43} 50:31]
  wire [63:0] _GEN_653 = 3'h2 == receive_num ? io_from_axi_rdata : receive_data_2; // @[d_cache.scala 137:{43,43} 50:31]
  wire [63:0] _GEN_654 = 3'h3 == receive_num ? io_from_axi_rdata : receive_data_3; // @[d_cache.scala 137:{43,43} 50:31]
  wire [63:0] _GEN_655 = 3'h4 == receive_num ? io_from_axi_rdata : receive_data_4; // @[d_cache.scala 137:{43,43} 50:31]
  wire [63:0] _GEN_656 = 3'h5 == receive_num ? io_from_axi_rdata : receive_data_5; // @[d_cache.scala 137:{43,43} 50:31]
  wire [63:0] _GEN_657 = 3'h6 == receive_num ? io_from_axi_rdata : receive_data_6; // @[d_cache.scala 137:{43,43} 50:31]
  wire [63:0] _GEN_658 = 3'h7 == receive_num ? io_from_axi_rdata : receive_data_7; // @[d_cache.scala 137:{43,43} 50:31]
  wire [2:0] _receive_num_T_1 = receive_num + 3'h1; // @[d_cache.scala 138:44]
  wire [3:0] _GEN_659 = io_from_axi_rlast ? 4'h5 : state; // @[d_cache.scala 139:40 140:27 82:24]
  wire [63:0] _GEN_660 = io_from_axi_rvalid ? _GEN_651 : receive_data_0; // @[d_cache.scala 136:37 50:31]
  wire [63:0] _GEN_661 = io_from_axi_rvalid ? _GEN_652 : receive_data_1; // @[d_cache.scala 136:37 50:31]
  wire [63:0] _GEN_662 = io_from_axi_rvalid ? _GEN_653 : receive_data_2; // @[d_cache.scala 136:37 50:31]
  wire [63:0] _GEN_663 = io_from_axi_rvalid ? _GEN_654 : receive_data_3; // @[d_cache.scala 136:37 50:31]
  wire [63:0] _GEN_664 = io_from_axi_rvalid ? _GEN_655 : receive_data_4; // @[d_cache.scala 136:37 50:31]
  wire [63:0] _GEN_665 = io_from_axi_rvalid ? _GEN_656 : receive_data_5; // @[d_cache.scala 136:37 50:31]
  wire [63:0] _GEN_666 = io_from_axi_rvalid ? _GEN_657 : receive_data_6; // @[d_cache.scala 136:37 50:31]
  wire [63:0] _GEN_667 = io_from_axi_rvalid ? _GEN_658 : receive_data_7; // @[d_cache.scala 136:37 50:31]
  wire [2:0] _GEN_668 = io_from_axi_rvalid ? _receive_num_T_1 : receive_num; // @[d_cache.scala 136:37 138:29 51:30]
  wire [3:0] _GEN_669 = io_from_axi_rvalid ? _GEN_659 : state; // @[d_cache.scala 136:37 82:24]
  wire [3:0] _GEN_670 = io_from_axi_bvalid ? 4'h0 : state; // @[d_cache.scala 145:37 146:23 82:24]
  wire [511:0] _ram_0_T_6 = {receive_data_7,receive_data_6,receive_data_5,receive_data_4,receive_data_3,receive_data_2,
    receive_data_1,receive_data_0}; // @[Cat.scala 31:58]
  wire [511:0] _GEN_671 = 4'h0 == index ? _ram_0_T_6 : ram_0_0; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_672 = 4'h1 == index ? _ram_0_T_6 : ram_0_1; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_673 = 4'h2 == index ? _ram_0_T_6 : ram_0_2; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_674 = 4'h3 == index ? _ram_0_T_6 : ram_0_3; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_675 = 4'h4 == index ? _ram_0_T_6 : ram_0_4; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_676 = 4'h5 == index ? _ram_0_T_6 : ram_0_5; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_677 = 4'h6 == index ? _ram_0_T_6 : ram_0_6; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_678 = 4'h7 == index ? _ram_0_T_6 : ram_0_7; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_679 = 4'h8 == index ? _ram_0_T_6 : ram_0_8; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_680 = 4'h9 == index ? _ram_0_T_6 : ram_0_9; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_681 = 4'ha == index ? _ram_0_T_6 : ram_0_10; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_682 = 4'hb == index ? _ram_0_T_6 : ram_0_11; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_683 = 4'hc == index ? _ram_0_T_6 : ram_0_12; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_684 = 4'hd == index ? _ram_0_T_6 : ram_0_13; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_685 = 4'he == index ? _ram_0_T_6 : ram_0_14; // @[d_cache.scala 152:{30,30} 19:24]
  wire [511:0] _GEN_686 = 4'hf == index ? _ram_0_T_6 : ram_0_15; // @[d_cache.scala 152:{30,30} 19:24]
  wire [31:0] _GEN_687 = 4'h0 == index ? _GEN_5341 : tag_0_0; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_688 = 4'h1 == index ? _GEN_5341 : tag_0_1; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_689 = 4'h2 == index ? _GEN_5341 : tag_0_2; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_690 = 4'h3 == index ? _GEN_5341 : tag_0_3; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_691 = 4'h4 == index ? _GEN_5341 : tag_0_4; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_692 = 4'h5 == index ? _GEN_5341 : tag_0_5; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_693 = 4'h6 == index ? _GEN_5341 : tag_0_6; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_694 = 4'h7 == index ? _GEN_5341 : tag_0_7; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_695 = 4'h8 == index ? _GEN_5341 : tag_0_8; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_696 = 4'h9 == index ? _GEN_5341 : tag_0_9; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_697 = 4'ha == index ? _GEN_5341 : tag_0_10; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_698 = 4'hb == index ? _GEN_5341 : tag_0_11; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_699 = 4'hc == index ? _GEN_5341 : tag_0_12; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_700 = 4'hd == index ? _GEN_5341 : tag_0_13; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_701 = 4'he == index ? _GEN_5341 : tag_0_14; // @[d_cache.scala 153:{30,30} 24:24]
  wire [31:0] _GEN_702 = 4'hf == index ? _GEN_5341 : tag_0_15; // @[d_cache.scala 153:{30,30} 24:24]
  wire  _GEN_703 = _GEN_5351 | valid_0_0; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_704 = _GEN_5356 | valid_0_1; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_705 = _GEN_5357 | valid_0_2; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_706 = _GEN_5361 | valid_0_3; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_707 = _GEN_5365 | valid_0_4; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_708 = _GEN_5367 | valid_0_5; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_709 = _GEN_5369 | valid_0_6; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_710 = _GEN_5370 | valid_0_7; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_711 = _GEN_5374 | valid_0_8; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_712 = _GEN_5375 | valid_0_9; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_713 = _GEN_5380 | valid_0_10; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_714 = _GEN_5381 | valid_0_11; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_715 = _GEN_5384 | valid_0_12; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_716 = _GEN_5388 | valid_0_13; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_717 = _GEN_5390 | valid_0_14; // @[d_cache.scala 154:{32,32} 29:26]
  wire  _GEN_718 = _GEN_5392 | valid_0_15; // @[d_cache.scala 154:{32,32} 29:26]
  wire [7:0] _GEN_720 = 4'h1 == index ? quene_1 : quene_0; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_721 = 4'h2 == index ? quene_2 : _GEN_720; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_722 = 4'h3 == index ? quene_3 : _GEN_721; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_723 = 4'h4 == index ? quene_4 : _GEN_722; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_724 = 4'h5 == index ? quene_5 : _GEN_723; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_725 = 4'h6 == index ? quene_6 : _GEN_724; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_726 = 4'h7 == index ? quene_7 : _GEN_725; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_727 = 4'h8 == index ? quene_8 : _GEN_726; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_728 = 4'h9 == index ? quene_9 : _GEN_727; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_729 = 4'ha == index ? quene_10 : _GEN_728; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_730 = 4'hb == index ? quene_11 : _GEN_729; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_731 = 4'hc == index ? quene_12 : _GEN_730; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_732 = 4'hd == index ? quene_13 : _GEN_731; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_733 = 4'he == index ? quene_14 : _GEN_732; // @[d_cache.scala 155:{46,46}]
  wire [7:0] _GEN_734 = 4'hf == index ? quene_15 : _GEN_733; // @[d_cache.scala 155:{46,46}]
  wire [9:0] _GEN_5513 = {_GEN_734, 2'h0}; // @[d_cache.scala 155:46]
  wire [10:0] _quene_T = {{1'd0}, _GEN_5513}; // @[d_cache.scala 155:46]
  wire [7:0] _GEN_735 = 4'h0 == index ? _quene_T[7:0] : quene_0; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_736 = 4'h1 == index ? _quene_T[7:0] : quene_1; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_737 = 4'h2 == index ? _quene_T[7:0] : quene_2; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_738 = 4'h3 == index ? _quene_T[7:0] : quene_3; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_739 = 4'h4 == index ? _quene_T[7:0] : quene_4; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_740 = 4'h5 == index ? _quene_T[7:0] : quene_5; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_741 = 4'h6 == index ? _quene_T[7:0] : quene_6; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_742 = 4'h7 == index ? _quene_T[7:0] : quene_7; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_743 = 4'h8 == index ? _quene_T[7:0] : quene_8; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_744 = 4'h9 == index ? _quene_T[7:0] : quene_9; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_745 = 4'ha == index ? _quene_T[7:0] : quene_10; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_746 = 4'hb == index ? _quene_T[7:0] : quene_11; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_747 = 4'hc == index ? _quene_T[7:0] : quene_12; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_748 = 4'hd == index ? _quene_T[7:0] : quene_13; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_749 = 4'he == index ? _quene_T[7:0] : quene_14; // @[d_cache.scala 155:{30,30} 52:24]
  wire [7:0] _GEN_750 = 4'hf == index ? _quene_T[7:0] : quene_15; // @[d_cache.scala 155:{30,30} 52:24]
  wire [511:0] _GEN_751 = 4'h0 == index ? _ram_0_T_6 : ram_1_0; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_752 = 4'h1 == index ? _ram_0_T_6 : ram_1_1; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_753 = 4'h2 == index ? _ram_0_T_6 : ram_1_2; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_754 = 4'h3 == index ? _ram_0_T_6 : ram_1_3; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_755 = 4'h4 == index ? _ram_0_T_6 : ram_1_4; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_756 = 4'h5 == index ? _ram_0_T_6 : ram_1_5; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_757 = 4'h6 == index ? _ram_0_T_6 : ram_1_6; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_758 = 4'h7 == index ? _ram_0_T_6 : ram_1_7; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_759 = 4'h8 == index ? _ram_0_T_6 : ram_1_8; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_760 = 4'h9 == index ? _ram_0_T_6 : ram_1_9; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_761 = 4'ha == index ? _ram_0_T_6 : ram_1_10; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_762 = 4'hb == index ? _ram_0_T_6 : ram_1_11; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_763 = 4'hc == index ? _ram_0_T_6 : ram_1_12; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_764 = 4'hd == index ? _ram_0_T_6 : ram_1_13; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_765 = 4'he == index ? _ram_0_T_6 : ram_1_14; // @[d_cache.scala 158:{30,30} 20:24]
  wire [511:0] _GEN_766 = 4'hf == index ? _ram_0_T_6 : ram_1_15; // @[d_cache.scala 158:{30,30} 20:24]
  wire [31:0] _GEN_767 = 4'h0 == index ? _GEN_5341 : tag_1_0; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_768 = 4'h1 == index ? _GEN_5341 : tag_1_1; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_769 = 4'h2 == index ? _GEN_5341 : tag_1_2; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_770 = 4'h3 == index ? _GEN_5341 : tag_1_3; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_771 = 4'h4 == index ? _GEN_5341 : tag_1_4; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_772 = 4'h5 == index ? _GEN_5341 : tag_1_5; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_773 = 4'h6 == index ? _GEN_5341 : tag_1_6; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_774 = 4'h7 == index ? _GEN_5341 : tag_1_7; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_775 = 4'h8 == index ? _GEN_5341 : tag_1_8; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_776 = 4'h9 == index ? _GEN_5341 : tag_1_9; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_777 = 4'ha == index ? _GEN_5341 : tag_1_10; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_778 = 4'hb == index ? _GEN_5341 : tag_1_11; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_779 = 4'hc == index ? _GEN_5341 : tag_1_12; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_780 = 4'hd == index ? _GEN_5341 : tag_1_13; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_781 = 4'he == index ? _GEN_5341 : tag_1_14; // @[d_cache.scala 159:{30,30} 25:24]
  wire [31:0] _GEN_782 = 4'hf == index ? _GEN_5341 : tag_1_15; // @[d_cache.scala 159:{30,30} 25:24]
  wire  _GEN_783 = _GEN_5351 | valid_1_0; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_784 = _GEN_5356 | valid_1_1; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_785 = _GEN_5357 | valid_1_2; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_786 = _GEN_5361 | valid_1_3; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_787 = _GEN_5365 | valid_1_4; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_788 = _GEN_5367 | valid_1_5; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_789 = _GEN_5369 | valid_1_6; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_790 = _GEN_5370 | valid_1_7; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_791 = _GEN_5374 | valid_1_8; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_792 = _GEN_5375 | valid_1_9; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_793 = _GEN_5380 | valid_1_10; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_794 = _GEN_5381 | valid_1_11; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_795 = _GEN_5384 | valid_1_12; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_796 = _GEN_5388 | valid_1_13; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_797 = _GEN_5390 | valid_1_14; // @[d_cache.scala 160:{32,32} 30:26]
  wire  _GEN_798 = _GEN_5392 | valid_1_15; // @[d_cache.scala 160:{32,32} 30:26]
  wire [10:0] _quene_T_2 = _quene_T | 11'h1; // @[d_cache.scala 161:55]
  wire [7:0] _GEN_799 = 4'h0 == index ? _quene_T_2[7:0] : quene_0; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_800 = 4'h1 == index ? _quene_T_2[7:0] : quene_1; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_801 = 4'h2 == index ? _quene_T_2[7:0] : quene_2; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_802 = 4'h3 == index ? _quene_T_2[7:0] : quene_3; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_803 = 4'h4 == index ? _quene_T_2[7:0] : quene_4; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_804 = 4'h5 == index ? _quene_T_2[7:0] : quene_5; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_805 = 4'h6 == index ? _quene_T_2[7:0] : quene_6; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_806 = 4'h7 == index ? _quene_T_2[7:0] : quene_7; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_807 = 4'h8 == index ? _quene_T_2[7:0] : quene_8; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_808 = 4'h9 == index ? _quene_T_2[7:0] : quene_9; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_809 = 4'ha == index ? _quene_T_2[7:0] : quene_10; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_810 = 4'hb == index ? _quene_T_2[7:0] : quene_11; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_811 = 4'hc == index ? _quene_T_2[7:0] : quene_12; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_812 = 4'hd == index ? _quene_T_2[7:0] : quene_13; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_813 = 4'he == index ? _quene_T_2[7:0] : quene_14; // @[d_cache.scala 161:{30,30} 52:24]
  wire [7:0] _GEN_814 = 4'hf == index ? _quene_T_2[7:0] : quene_15; // @[d_cache.scala 161:{30,30} 52:24]
  wire [511:0] _GEN_815 = 4'h0 == index ? _ram_0_T_6 : ram_2_0; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_816 = 4'h1 == index ? _ram_0_T_6 : ram_2_1; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_817 = 4'h2 == index ? _ram_0_T_6 : ram_2_2; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_818 = 4'h3 == index ? _ram_0_T_6 : ram_2_3; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_819 = 4'h4 == index ? _ram_0_T_6 : ram_2_4; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_820 = 4'h5 == index ? _ram_0_T_6 : ram_2_5; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_821 = 4'h6 == index ? _ram_0_T_6 : ram_2_6; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_822 = 4'h7 == index ? _ram_0_T_6 : ram_2_7; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_823 = 4'h8 == index ? _ram_0_T_6 : ram_2_8; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_824 = 4'h9 == index ? _ram_0_T_6 : ram_2_9; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_825 = 4'ha == index ? _ram_0_T_6 : ram_2_10; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_826 = 4'hb == index ? _ram_0_T_6 : ram_2_11; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_827 = 4'hc == index ? _ram_0_T_6 : ram_2_12; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_828 = 4'hd == index ? _ram_0_T_6 : ram_2_13; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_829 = 4'he == index ? _ram_0_T_6 : ram_2_14; // @[d_cache.scala 164:{30,30} 21:24]
  wire [511:0] _GEN_830 = 4'hf == index ? _ram_0_T_6 : ram_2_15; // @[d_cache.scala 164:{30,30} 21:24]
  wire [31:0] _GEN_831 = 4'h0 == index ? _GEN_5341 : tag_2_0; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_832 = 4'h1 == index ? _GEN_5341 : tag_2_1; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_833 = 4'h2 == index ? _GEN_5341 : tag_2_2; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_834 = 4'h3 == index ? _GEN_5341 : tag_2_3; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_835 = 4'h4 == index ? _GEN_5341 : tag_2_4; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_836 = 4'h5 == index ? _GEN_5341 : tag_2_5; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_837 = 4'h6 == index ? _GEN_5341 : tag_2_6; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_838 = 4'h7 == index ? _GEN_5341 : tag_2_7; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_839 = 4'h8 == index ? _GEN_5341 : tag_2_8; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_840 = 4'h9 == index ? _GEN_5341 : tag_2_9; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_841 = 4'ha == index ? _GEN_5341 : tag_2_10; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_842 = 4'hb == index ? _GEN_5341 : tag_2_11; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_843 = 4'hc == index ? _GEN_5341 : tag_2_12; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_844 = 4'hd == index ? _GEN_5341 : tag_2_13; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_845 = 4'he == index ? _GEN_5341 : tag_2_14; // @[d_cache.scala 165:{30,30} 26:24]
  wire [31:0] _GEN_846 = 4'hf == index ? _GEN_5341 : tag_2_15; // @[d_cache.scala 165:{30,30} 26:24]
  wire  _GEN_847 = _GEN_5351 | valid_2_0; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_848 = _GEN_5356 | valid_2_1; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_849 = _GEN_5357 | valid_2_2; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_850 = _GEN_5361 | valid_2_3; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_851 = _GEN_5365 | valid_2_4; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_852 = _GEN_5367 | valid_2_5; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_853 = _GEN_5369 | valid_2_6; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_854 = _GEN_5370 | valid_2_7; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_855 = _GEN_5374 | valid_2_8; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_856 = _GEN_5375 | valid_2_9; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_857 = _GEN_5380 | valid_2_10; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_858 = _GEN_5381 | valid_2_11; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_859 = _GEN_5384 | valid_2_12; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_860 = _GEN_5388 | valid_2_13; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_861 = _GEN_5390 | valid_2_14; // @[d_cache.scala 166:{32,32} 31:26]
  wire  _GEN_862 = _GEN_5392 | valid_2_15; // @[d_cache.scala 166:{32,32} 31:26]
  wire [10:0] _quene_T_4 = _quene_T | 11'h2; // @[d_cache.scala 167:55]
  wire [7:0] _GEN_863 = 4'h0 == index ? _quene_T_4[7:0] : quene_0; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_864 = 4'h1 == index ? _quene_T_4[7:0] : quene_1; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_865 = 4'h2 == index ? _quene_T_4[7:0] : quene_2; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_866 = 4'h3 == index ? _quene_T_4[7:0] : quene_3; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_867 = 4'h4 == index ? _quene_T_4[7:0] : quene_4; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_868 = 4'h5 == index ? _quene_T_4[7:0] : quene_5; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_869 = 4'h6 == index ? _quene_T_4[7:0] : quene_6; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_870 = 4'h7 == index ? _quene_T_4[7:0] : quene_7; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_871 = 4'h8 == index ? _quene_T_4[7:0] : quene_8; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_872 = 4'h9 == index ? _quene_T_4[7:0] : quene_9; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_873 = 4'ha == index ? _quene_T_4[7:0] : quene_10; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_874 = 4'hb == index ? _quene_T_4[7:0] : quene_11; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_875 = 4'hc == index ? _quene_T_4[7:0] : quene_12; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_876 = 4'hd == index ? _quene_T_4[7:0] : quene_13; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_877 = 4'he == index ? _quene_T_4[7:0] : quene_14; // @[d_cache.scala 167:{30,30} 52:24]
  wire [7:0] _GEN_878 = 4'hf == index ? _quene_T_4[7:0] : quene_15; // @[d_cache.scala 167:{30,30} 52:24]
  wire [511:0] _GEN_879 = 4'h0 == index ? _ram_0_T_6 : ram_3_0; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_880 = 4'h1 == index ? _ram_0_T_6 : ram_3_1; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_881 = 4'h2 == index ? _ram_0_T_6 : ram_3_2; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_882 = 4'h3 == index ? _ram_0_T_6 : ram_3_3; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_883 = 4'h4 == index ? _ram_0_T_6 : ram_3_4; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_884 = 4'h5 == index ? _ram_0_T_6 : ram_3_5; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_885 = 4'h6 == index ? _ram_0_T_6 : ram_3_6; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_886 = 4'h7 == index ? _ram_0_T_6 : ram_3_7; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_887 = 4'h8 == index ? _ram_0_T_6 : ram_3_8; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_888 = 4'h9 == index ? _ram_0_T_6 : ram_3_9; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_889 = 4'ha == index ? _ram_0_T_6 : ram_3_10; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_890 = 4'hb == index ? _ram_0_T_6 : ram_3_11; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_891 = 4'hc == index ? _ram_0_T_6 : ram_3_12; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_892 = 4'hd == index ? _ram_0_T_6 : ram_3_13; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_893 = 4'he == index ? _ram_0_T_6 : ram_3_14; // @[d_cache.scala 170:{30,30} 22:24]
  wire [511:0] _GEN_894 = 4'hf == index ? _ram_0_T_6 : ram_3_15; // @[d_cache.scala 170:{30,30} 22:24]
  wire [31:0] _GEN_895 = 4'h0 == index ? _GEN_5341 : tag_3_0; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_896 = 4'h1 == index ? _GEN_5341 : tag_3_1; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_897 = 4'h2 == index ? _GEN_5341 : tag_3_2; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_898 = 4'h3 == index ? _GEN_5341 : tag_3_3; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_899 = 4'h4 == index ? _GEN_5341 : tag_3_4; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_900 = 4'h5 == index ? _GEN_5341 : tag_3_5; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_901 = 4'h6 == index ? _GEN_5341 : tag_3_6; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_902 = 4'h7 == index ? _GEN_5341 : tag_3_7; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_903 = 4'h8 == index ? _GEN_5341 : tag_3_8; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_904 = 4'h9 == index ? _GEN_5341 : tag_3_9; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_905 = 4'ha == index ? _GEN_5341 : tag_3_10; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_906 = 4'hb == index ? _GEN_5341 : tag_3_11; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_907 = 4'hc == index ? _GEN_5341 : tag_3_12; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_908 = 4'hd == index ? _GEN_5341 : tag_3_13; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_909 = 4'he == index ? _GEN_5341 : tag_3_14; // @[d_cache.scala 171:{30,30} 27:24]
  wire [31:0] _GEN_910 = 4'hf == index ? _GEN_5341 : tag_3_15; // @[d_cache.scala 171:{30,30} 27:24]
  wire  _GEN_911 = _GEN_5351 | valid_3_0; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_912 = _GEN_5356 | valid_3_1; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_913 = _GEN_5357 | valid_3_2; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_914 = _GEN_5361 | valid_3_3; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_915 = _GEN_5365 | valid_3_4; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_916 = _GEN_5367 | valid_3_5; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_917 = _GEN_5369 | valid_3_6; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_918 = _GEN_5370 | valid_3_7; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_919 = _GEN_5374 | valid_3_8; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_920 = _GEN_5375 | valid_3_9; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_921 = _GEN_5380 | valid_3_10; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_922 = _GEN_5381 | valid_3_11; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_923 = _GEN_5384 | valid_3_12; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_924 = _GEN_5388 | valid_3_13; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_925 = _GEN_5390 | valid_3_14; // @[d_cache.scala 172:{32,32} 32:26]
  wire  _GEN_926 = _GEN_5392 | valid_3_15; // @[d_cache.scala 172:{32,32} 32:26]
  wire [10:0] _quene_T_6 = _quene_T | 11'h3; // @[d_cache.scala 173:55]
  wire [7:0] _GEN_927 = 4'h0 == index ? _quene_T_6[7:0] : quene_0; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_928 = 4'h1 == index ? _quene_T_6[7:0] : quene_1; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_929 = 4'h2 == index ? _quene_T_6[7:0] : quene_2; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_930 = 4'h3 == index ? _quene_T_6[7:0] : quene_3; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_931 = 4'h4 == index ? _quene_T_6[7:0] : quene_4; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_932 = 4'h5 == index ? _quene_T_6[7:0] : quene_5; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_933 = 4'h6 == index ? _quene_T_6[7:0] : quene_6; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_934 = 4'h7 == index ? _quene_T_6[7:0] : quene_7; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_935 = 4'h8 == index ? _quene_T_6[7:0] : quene_8; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_936 = 4'h9 == index ? _quene_T_6[7:0] : quene_9; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_937 = 4'ha == index ? _quene_T_6[7:0] : quene_10; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_938 = 4'hb == index ? _quene_T_6[7:0] : quene_11; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_939 = 4'hc == index ? _quene_T_6[7:0] : quene_12; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_940 = 4'hd == index ? _quene_T_6[7:0] : quene_13; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_941 = 4'he == index ? _quene_T_6[7:0] : quene_14; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_942 = 4'hf == index ? _quene_T_6[7:0] : quene_15; // @[d_cache.scala 173:{30,30} 52:24]
  wire  _GEN_944 = 4'h1 == index ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_945 = 4'h2 == index ? dirty_0_2 : _GEN_944; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_946 = 4'h3 == index ? dirty_0_3 : _GEN_945; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_947 = 4'h4 == index ? dirty_0_4 : _GEN_946; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_948 = 4'h5 == index ? dirty_0_5 : _GEN_947; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_949 = 4'h6 == index ? dirty_0_6 : _GEN_948; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_950 = 4'h7 == index ? dirty_0_7 : _GEN_949; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_951 = 4'h8 == index ? dirty_0_8 : _GEN_950; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_952 = 4'h9 == index ? dirty_0_9 : _GEN_951; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_953 = 4'ha == index ? dirty_0_10 : _GEN_952; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_954 = 4'hb == index ? dirty_0_11 : _GEN_953; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_955 = 4'hc == index ? dirty_0_12 : _GEN_954; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_956 = 4'hd == index ? dirty_0_13 : _GEN_955; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_957 = 4'he == index ? dirty_0_14 : _GEN_956; // @[d_cache.scala 176:{40,40}]
  wire  _GEN_958 = 4'hf == index ? dirty_0_15 : _GEN_957; // @[d_cache.scala 176:{40,40}]
  wire [41:0] _write_back_addr_T_1 = {_GEN_15,index,6'h0}; // @[Cat.scala 31:58]
  wire  _GEN_991 = 4'h0 == index ? 1'h0 : dirty_0_0; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_992 = 4'h1 == index ? 1'h0 : dirty_0_1; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_993 = 4'h2 == index ? 1'h0 : dirty_0_2; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_994 = 4'h3 == index ? 1'h0 : dirty_0_3; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_995 = 4'h4 == index ? 1'h0 : dirty_0_4; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_996 = 4'h5 == index ? 1'h0 : dirty_0_5; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_997 = 4'h6 == index ? 1'h0 : dirty_0_6; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_998 = 4'h7 == index ? 1'h0 : dirty_0_7; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_999 = 4'h8 == index ? 1'h0 : dirty_0_8; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_1000 = 4'h9 == index ? 1'h0 : dirty_0_9; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_1001 = 4'ha == index ? 1'h0 : dirty_0_10; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_1002 = 4'hb == index ? 1'h0 : dirty_0_11; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_1003 = 4'hc == index ? 1'h0 : dirty_0_12; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_1004 = 4'hd == index ? 1'h0 : dirty_0_13; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_1005 = 4'he == index ? 1'h0 : dirty_0_14; // @[d_cache.scala 181:{40,40} 34:26]
  wire  _GEN_1006 = 4'hf == index ? 1'h0 : dirty_0_15; // @[d_cache.scala 181:{40,40} 34:26]
  wire [511:0] _GEN_1103 = _GEN_958 ? _GEN_150 : write_back_data; // @[d_cache.scala 176:47 177:41 44:34]
  wire [41:0] _GEN_1104 = _GEN_958 ? _write_back_addr_T_1 : {{10'd0}, write_back_addr}; // @[d_cache.scala 176:47 178:41 45:34]
  wire [511:0] _GEN_1105 = _GEN_958 ? _GEN_671 : _GEN_671; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1106 = _GEN_958 ? _GEN_672 : _GEN_672; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1107 = _GEN_958 ? _GEN_673 : _GEN_673; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1108 = _GEN_958 ? _GEN_674 : _GEN_674; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1109 = _GEN_958 ? _GEN_675 : _GEN_675; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1110 = _GEN_958 ? _GEN_676 : _GEN_676; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1111 = _GEN_958 ? _GEN_677 : _GEN_677; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1112 = _GEN_958 ? _GEN_678 : _GEN_678; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1113 = _GEN_958 ? _GEN_679 : _GEN_679; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1114 = _GEN_958 ? _GEN_680 : _GEN_680; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1115 = _GEN_958 ? _GEN_681 : _GEN_681; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1116 = _GEN_958 ? _GEN_682 : _GEN_682; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1117 = _GEN_958 ? _GEN_683 : _GEN_683; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1118 = _GEN_958 ? _GEN_684 : _GEN_684; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1119 = _GEN_958 ? _GEN_685 : _GEN_685; // @[d_cache.scala 176:47]
  wire [511:0] _GEN_1120 = _GEN_958 ? _GEN_686 : _GEN_686; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1121 = _GEN_958 ? _GEN_687 : _GEN_687; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1122 = _GEN_958 ? _GEN_688 : _GEN_688; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1123 = _GEN_958 ? _GEN_689 : _GEN_689; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1124 = _GEN_958 ? _GEN_690 : _GEN_690; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1125 = _GEN_958 ? _GEN_691 : _GEN_691; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1126 = _GEN_958 ? _GEN_692 : _GEN_692; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1127 = _GEN_958 ? _GEN_693 : _GEN_693; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1128 = _GEN_958 ? _GEN_694 : _GEN_694; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1129 = _GEN_958 ? _GEN_695 : _GEN_695; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1130 = _GEN_958 ? _GEN_696 : _GEN_696; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1131 = _GEN_958 ? _GEN_697 : _GEN_697; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1132 = _GEN_958 ? _GEN_698 : _GEN_698; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1133 = _GEN_958 ? _GEN_699 : _GEN_699; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1134 = _GEN_958 ? _GEN_700 : _GEN_700; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1135 = _GEN_958 ? _GEN_701 : _GEN_701; // @[d_cache.scala 176:47]
  wire [31:0] _GEN_1136 = _GEN_958 ? _GEN_702 : _GEN_702; // @[d_cache.scala 176:47]
  wire  _GEN_1137 = _GEN_958 ? _GEN_991 : dirty_0_0; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1138 = _GEN_958 ? _GEN_992 : dirty_0_1; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1139 = _GEN_958 ? _GEN_993 : dirty_0_2; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1140 = _GEN_958 ? _GEN_994 : dirty_0_3; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1141 = _GEN_958 ? _GEN_995 : dirty_0_4; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1142 = _GEN_958 ? _GEN_996 : dirty_0_5; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1143 = _GEN_958 ? _GEN_997 : dirty_0_6; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1144 = _GEN_958 ? _GEN_998 : dirty_0_7; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1145 = _GEN_958 ? _GEN_999 : dirty_0_8; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1146 = _GEN_958 ? _GEN_1000 : dirty_0_9; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1147 = _GEN_958 ? _GEN_1001 : dirty_0_10; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1148 = _GEN_958 ? _GEN_1002 : dirty_0_11; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1149 = _GEN_958 ? _GEN_1003 : dirty_0_12; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1150 = _GEN_958 ? _GEN_1004 : dirty_0_13; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1151 = _GEN_958 ? _GEN_1005 : dirty_0_14; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1152 = _GEN_958 ? _GEN_1006 : dirty_0_15; // @[d_cache.scala 176:47 34:26]
  wire  _GEN_1153 = _GEN_958 ? _GEN_703 : _GEN_703; // @[d_cache.scala 176:47]
  wire  _GEN_1154 = _GEN_958 ? _GEN_704 : _GEN_704; // @[d_cache.scala 176:47]
  wire  _GEN_1155 = _GEN_958 ? _GEN_705 : _GEN_705; // @[d_cache.scala 176:47]
  wire  _GEN_1156 = _GEN_958 ? _GEN_706 : _GEN_706; // @[d_cache.scala 176:47]
  wire  _GEN_1157 = _GEN_958 ? _GEN_707 : _GEN_707; // @[d_cache.scala 176:47]
  wire  _GEN_1158 = _GEN_958 ? _GEN_708 : _GEN_708; // @[d_cache.scala 176:47]
  wire  _GEN_1159 = _GEN_958 ? _GEN_709 : _GEN_709; // @[d_cache.scala 176:47]
  wire  _GEN_1160 = _GEN_958 ? _GEN_710 : _GEN_710; // @[d_cache.scala 176:47]
  wire  _GEN_1161 = _GEN_958 ? _GEN_711 : _GEN_711; // @[d_cache.scala 176:47]
  wire  _GEN_1162 = _GEN_958 ? _GEN_712 : _GEN_712; // @[d_cache.scala 176:47]
  wire  _GEN_1163 = _GEN_958 ? _GEN_713 : _GEN_713; // @[d_cache.scala 176:47]
  wire  _GEN_1164 = _GEN_958 ? _GEN_714 : _GEN_714; // @[d_cache.scala 176:47]
  wire  _GEN_1165 = _GEN_958 ? _GEN_715 : _GEN_715; // @[d_cache.scala 176:47]
  wire  _GEN_1166 = _GEN_958 ? _GEN_716 : _GEN_716; // @[d_cache.scala 176:47]
  wire  _GEN_1167 = _GEN_958 ? _GEN_717 : _GEN_717; // @[d_cache.scala 176:47]
  wire  _GEN_1168 = _GEN_958 ? _GEN_718 : _GEN_718; // @[d_cache.scala 176:47]
  wire [3:0] _GEN_1169 = _GEN_958 ? 4'h6 : 4'h1; // @[d_cache.scala 176:47 183:31 186:31]
  wire [7:0] _GEN_1170 = _GEN_958 ? _GEN_735 : _GEN_735; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1171 = _GEN_958 ? _GEN_736 : _GEN_736; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1172 = _GEN_958 ? _GEN_737 : _GEN_737; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1173 = _GEN_958 ? _GEN_738 : _GEN_738; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1174 = _GEN_958 ? _GEN_739 : _GEN_739; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1175 = _GEN_958 ? _GEN_740 : _GEN_740; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1176 = _GEN_958 ? _GEN_741 : _GEN_741; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1177 = _GEN_958 ? _GEN_742 : _GEN_742; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1178 = _GEN_958 ? _GEN_743 : _GEN_743; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1179 = _GEN_958 ? _GEN_744 : _GEN_744; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1180 = _GEN_958 ? _GEN_745 : _GEN_745; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1181 = _GEN_958 ? _GEN_746 : _GEN_746; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1182 = _GEN_958 ? _GEN_747 : _GEN_747; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1183 = _GEN_958 ? _GEN_748 : _GEN_748; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1184 = _GEN_958 ? _GEN_749 : _GEN_749; // @[d_cache.scala 176:47]
  wire [7:0] _GEN_1185 = _GEN_958 ? _GEN_750 : _GEN_750; // @[d_cache.scala 176:47]
  wire  _GEN_1187 = 4'h1 == index ? dirty_1_1 : dirty_1_0; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1188 = 4'h2 == index ? dirty_1_2 : _GEN_1187; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1189 = 4'h3 == index ? dirty_1_3 : _GEN_1188; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1190 = 4'h4 == index ? dirty_1_4 : _GEN_1189; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1191 = 4'h5 == index ? dirty_1_5 : _GEN_1190; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1192 = 4'h6 == index ? dirty_1_6 : _GEN_1191; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1193 = 4'h7 == index ? dirty_1_7 : _GEN_1192; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1194 = 4'h8 == index ? dirty_1_8 : _GEN_1193; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1195 = 4'h9 == index ? dirty_1_9 : _GEN_1194; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1196 = 4'ha == index ? dirty_1_10 : _GEN_1195; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1197 = 4'hb == index ? dirty_1_11 : _GEN_1196; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1198 = 4'hc == index ? dirty_1_12 : _GEN_1197; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1199 = 4'hd == index ? dirty_1_13 : _GEN_1198; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1200 = 4'he == index ? dirty_1_14 : _GEN_1199; // @[d_cache.scala 193:{40,40}]
  wire  _GEN_1201 = 4'hf == index ? dirty_1_15 : _GEN_1200; // @[d_cache.scala 193:{40,40}]
  wire [41:0] _write_back_addr_T_3 = {_GEN_47,index,6'h0}; // @[Cat.scala 31:58]
  wire  _GEN_1234 = 4'h0 == index ? 1'h0 : dirty_1_0; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1235 = 4'h1 == index ? 1'h0 : dirty_1_1; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1236 = 4'h2 == index ? 1'h0 : dirty_1_2; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1237 = 4'h3 == index ? 1'h0 : dirty_1_3; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1238 = 4'h4 == index ? 1'h0 : dirty_1_4; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1239 = 4'h5 == index ? 1'h0 : dirty_1_5; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1240 = 4'h6 == index ? 1'h0 : dirty_1_6; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1241 = 4'h7 == index ? 1'h0 : dirty_1_7; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1242 = 4'h8 == index ? 1'h0 : dirty_1_8; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1243 = 4'h9 == index ? 1'h0 : dirty_1_9; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1244 = 4'ha == index ? 1'h0 : dirty_1_10; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1245 = 4'hb == index ? 1'h0 : dirty_1_11; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1246 = 4'hc == index ? 1'h0 : dirty_1_12; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1247 = 4'hd == index ? 1'h0 : dirty_1_13; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1248 = 4'he == index ? 1'h0 : dirty_1_14; // @[d_cache.scala 198:{40,40} 35:26]
  wire  _GEN_1249 = 4'hf == index ? 1'h0 : dirty_1_15; // @[d_cache.scala 198:{40,40} 35:26]
  wire [511:0] _GEN_1346 = _GEN_1201 ? _GEN_198 : write_back_data; // @[d_cache.scala 193:47 194:41 44:34]
  wire [41:0] _GEN_1347 = _GEN_1201 ? _write_back_addr_T_3 : {{10'd0}, write_back_addr}; // @[d_cache.scala 193:47 195:41 45:34]
  wire [511:0] _GEN_1348 = _GEN_1201 ? _GEN_751 : _GEN_751; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1349 = _GEN_1201 ? _GEN_752 : _GEN_752; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1350 = _GEN_1201 ? _GEN_753 : _GEN_753; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1351 = _GEN_1201 ? _GEN_754 : _GEN_754; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1352 = _GEN_1201 ? _GEN_755 : _GEN_755; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1353 = _GEN_1201 ? _GEN_756 : _GEN_756; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1354 = _GEN_1201 ? _GEN_757 : _GEN_757; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1355 = _GEN_1201 ? _GEN_758 : _GEN_758; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1356 = _GEN_1201 ? _GEN_759 : _GEN_759; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1357 = _GEN_1201 ? _GEN_760 : _GEN_760; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1358 = _GEN_1201 ? _GEN_761 : _GEN_761; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1359 = _GEN_1201 ? _GEN_762 : _GEN_762; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1360 = _GEN_1201 ? _GEN_763 : _GEN_763; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1361 = _GEN_1201 ? _GEN_764 : _GEN_764; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1362 = _GEN_1201 ? _GEN_765 : _GEN_765; // @[d_cache.scala 193:47]
  wire [511:0] _GEN_1363 = _GEN_1201 ? _GEN_766 : _GEN_766; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1364 = _GEN_1201 ? _GEN_767 : _GEN_767; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1365 = _GEN_1201 ? _GEN_768 : _GEN_768; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1366 = _GEN_1201 ? _GEN_769 : _GEN_769; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1367 = _GEN_1201 ? _GEN_770 : _GEN_770; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1368 = _GEN_1201 ? _GEN_771 : _GEN_771; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1369 = _GEN_1201 ? _GEN_772 : _GEN_772; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1370 = _GEN_1201 ? _GEN_773 : _GEN_773; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1371 = _GEN_1201 ? _GEN_774 : _GEN_774; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1372 = _GEN_1201 ? _GEN_775 : _GEN_775; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1373 = _GEN_1201 ? _GEN_776 : _GEN_776; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1374 = _GEN_1201 ? _GEN_777 : _GEN_777; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1375 = _GEN_1201 ? _GEN_778 : _GEN_778; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1376 = _GEN_1201 ? _GEN_779 : _GEN_779; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1377 = _GEN_1201 ? _GEN_780 : _GEN_780; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1378 = _GEN_1201 ? _GEN_781 : _GEN_781; // @[d_cache.scala 193:47]
  wire [31:0] _GEN_1379 = _GEN_1201 ? _GEN_782 : _GEN_782; // @[d_cache.scala 193:47]
  wire  _GEN_1380 = _GEN_1201 ? _GEN_1234 : dirty_1_0; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1381 = _GEN_1201 ? _GEN_1235 : dirty_1_1; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1382 = _GEN_1201 ? _GEN_1236 : dirty_1_2; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1383 = _GEN_1201 ? _GEN_1237 : dirty_1_3; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1384 = _GEN_1201 ? _GEN_1238 : dirty_1_4; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1385 = _GEN_1201 ? _GEN_1239 : dirty_1_5; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1386 = _GEN_1201 ? _GEN_1240 : dirty_1_6; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1387 = _GEN_1201 ? _GEN_1241 : dirty_1_7; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1388 = _GEN_1201 ? _GEN_1242 : dirty_1_8; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1389 = _GEN_1201 ? _GEN_1243 : dirty_1_9; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1390 = _GEN_1201 ? _GEN_1244 : dirty_1_10; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1391 = _GEN_1201 ? _GEN_1245 : dirty_1_11; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1392 = _GEN_1201 ? _GEN_1246 : dirty_1_12; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1393 = _GEN_1201 ? _GEN_1247 : dirty_1_13; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1394 = _GEN_1201 ? _GEN_1248 : dirty_1_14; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1395 = _GEN_1201 ? _GEN_1249 : dirty_1_15; // @[d_cache.scala 193:47 35:26]
  wire  _GEN_1396 = _GEN_1201 ? _GEN_783 : _GEN_783; // @[d_cache.scala 193:47]
  wire  _GEN_1397 = _GEN_1201 ? _GEN_784 : _GEN_784; // @[d_cache.scala 193:47]
  wire  _GEN_1398 = _GEN_1201 ? _GEN_785 : _GEN_785; // @[d_cache.scala 193:47]
  wire  _GEN_1399 = _GEN_1201 ? _GEN_786 : _GEN_786; // @[d_cache.scala 193:47]
  wire  _GEN_1400 = _GEN_1201 ? _GEN_787 : _GEN_787; // @[d_cache.scala 193:47]
  wire  _GEN_1401 = _GEN_1201 ? _GEN_788 : _GEN_788; // @[d_cache.scala 193:47]
  wire  _GEN_1402 = _GEN_1201 ? _GEN_789 : _GEN_789; // @[d_cache.scala 193:47]
  wire  _GEN_1403 = _GEN_1201 ? _GEN_790 : _GEN_790; // @[d_cache.scala 193:47]
  wire  _GEN_1404 = _GEN_1201 ? _GEN_791 : _GEN_791; // @[d_cache.scala 193:47]
  wire  _GEN_1405 = _GEN_1201 ? _GEN_792 : _GEN_792; // @[d_cache.scala 193:47]
  wire  _GEN_1406 = _GEN_1201 ? _GEN_793 : _GEN_793; // @[d_cache.scala 193:47]
  wire  _GEN_1407 = _GEN_1201 ? _GEN_794 : _GEN_794; // @[d_cache.scala 193:47]
  wire  _GEN_1408 = _GEN_1201 ? _GEN_795 : _GEN_795; // @[d_cache.scala 193:47]
  wire  _GEN_1409 = _GEN_1201 ? _GEN_796 : _GEN_796; // @[d_cache.scala 193:47]
  wire  _GEN_1410 = _GEN_1201 ? _GEN_797 : _GEN_797; // @[d_cache.scala 193:47]
  wire  _GEN_1411 = _GEN_1201 ? _GEN_798 : _GEN_798; // @[d_cache.scala 193:47]
  wire [3:0] _GEN_1412 = _GEN_1201 ? 4'h6 : 4'h1; // @[d_cache.scala 193:47 200:31 203:31]
  wire [7:0] _GEN_1413 = _GEN_1201 ? _GEN_799 : _GEN_799; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1414 = _GEN_1201 ? _GEN_800 : _GEN_800; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1415 = _GEN_1201 ? _GEN_801 : _GEN_801; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1416 = _GEN_1201 ? _GEN_802 : _GEN_802; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1417 = _GEN_1201 ? _GEN_803 : _GEN_803; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1418 = _GEN_1201 ? _GEN_804 : _GEN_804; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1419 = _GEN_1201 ? _GEN_805 : _GEN_805; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1420 = _GEN_1201 ? _GEN_806 : _GEN_806; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1421 = _GEN_1201 ? _GEN_807 : _GEN_807; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1422 = _GEN_1201 ? _GEN_808 : _GEN_808; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1423 = _GEN_1201 ? _GEN_809 : _GEN_809; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1424 = _GEN_1201 ? _GEN_810 : _GEN_810; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1425 = _GEN_1201 ? _GEN_811 : _GEN_811; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1426 = _GEN_1201 ? _GEN_812 : _GEN_812; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1427 = _GEN_1201 ? _GEN_813 : _GEN_813; // @[d_cache.scala 193:47]
  wire [7:0] _GEN_1428 = _GEN_1201 ? _GEN_814 : _GEN_814; // @[d_cache.scala 193:47]
  wire  _GEN_1430 = 4'h1 == index ? dirty_2_1 : dirty_2_0; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1431 = 4'h2 == index ? dirty_2_2 : _GEN_1430; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1432 = 4'h3 == index ? dirty_2_3 : _GEN_1431; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1433 = 4'h4 == index ? dirty_2_4 : _GEN_1432; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1434 = 4'h5 == index ? dirty_2_5 : _GEN_1433; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1435 = 4'h6 == index ? dirty_2_6 : _GEN_1434; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1436 = 4'h7 == index ? dirty_2_7 : _GEN_1435; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1437 = 4'h8 == index ? dirty_2_8 : _GEN_1436; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1438 = 4'h9 == index ? dirty_2_9 : _GEN_1437; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1439 = 4'ha == index ? dirty_2_10 : _GEN_1438; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1440 = 4'hb == index ? dirty_2_11 : _GEN_1439; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1441 = 4'hc == index ? dirty_2_12 : _GEN_1440; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1442 = 4'hd == index ? dirty_2_13 : _GEN_1441; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1443 = 4'he == index ? dirty_2_14 : _GEN_1442; // @[d_cache.scala 210:{40,40}]
  wire  _GEN_1444 = 4'hf == index ? dirty_2_15 : _GEN_1443; // @[d_cache.scala 210:{40,40}]
  wire [41:0] _write_back_addr_T_5 = {_GEN_79,index,6'h0}; // @[Cat.scala 31:58]
  wire  _GEN_1477 = 4'h0 == index ? 1'h0 : dirty_2_0; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1478 = 4'h1 == index ? 1'h0 : dirty_2_1; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1479 = 4'h2 == index ? 1'h0 : dirty_2_2; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1480 = 4'h3 == index ? 1'h0 : dirty_2_3; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1481 = 4'h4 == index ? 1'h0 : dirty_2_4; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1482 = 4'h5 == index ? 1'h0 : dirty_2_5; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1483 = 4'h6 == index ? 1'h0 : dirty_2_6; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1484 = 4'h7 == index ? 1'h0 : dirty_2_7; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1485 = 4'h8 == index ? 1'h0 : dirty_2_8; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1486 = 4'h9 == index ? 1'h0 : dirty_2_9; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1487 = 4'ha == index ? 1'h0 : dirty_2_10; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1488 = 4'hb == index ? 1'h0 : dirty_2_11; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1489 = 4'hc == index ? 1'h0 : dirty_2_12; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1490 = 4'hd == index ? 1'h0 : dirty_2_13; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1491 = 4'he == index ? 1'h0 : dirty_2_14; // @[d_cache.scala 215:{40,40} 36:26]
  wire  _GEN_1492 = 4'hf == index ? 1'h0 : dirty_2_15; // @[d_cache.scala 215:{40,40} 36:26]
  wire [511:0] _GEN_1589 = _GEN_1444 ? _GEN_246 : write_back_data; // @[d_cache.scala 210:47 211:41 44:34]
  wire [41:0] _GEN_1590 = _GEN_1444 ? _write_back_addr_T_5 : {{10'd0}, write_back_addr}; // @[d_cache.scala 210:47 212:41 45:34]
  wire [511:0] _GEN_1591 = _GEN_1444 ? _GEN_815 : _GEN_815; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1592 = _GEN_1444 ? _GEN_816 : _GEN_816; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1593 = _GEN_1444 ? _GEN_817 : _GEN_817; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1594 = _GEN_1444 ? _GEN_818 : _GEN_818; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1595 = _GEN_1444 ? _GEN_819 : _GEN_819; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1596 = _GEN_1444 ? _GEN_820 : _GEN_820; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1597 = _GEN_1444 ? _GEN_821 : _GEN_821; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1598 = _GEN_1444 ? _GEN_822 : _GEN_822; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1599 = _GEN_1444 ? _GEN_823 : _GEN_823; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1600 = _GEN_1444 ? _GEN_824 : _GEN_824; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1601 = _GEN_1444 ? _GEN_825 : _GEN_825; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1602 = _GEN_1444 ? _GEN_826 : _GEN_826; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1603 = _GEN_1444 ? _GEN_827 : _GEN_827; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1604 = _GEN_1444 ? _GEN_828 : _GEN_828; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1605 = _GEN_1444 ? _GEN_829 : _GEN_829; // @[d_cache.scala 210:47]
  wire [511:0] _GEN_1606 = _GEN_1444 ? _GEN_830 : _GEN_830; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1607 = _GEN_1444 ? _GEN_831 : _GEN_831; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1608 = _GEN_1444 ? _GEN_832 : _GEN_832; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1609 = _GEN_1444 ? _GEN_833 : _GEN_833; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1610 = _GEN_1444 ? _GEN_834 : _GEN_834; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1611 = _GEN_1444 ? _GEN_835 : _GEN_835; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1612 = _GEN_1444 ? _GEN_836 : _GEN_836; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1613 = _GEN_1444 ? _GEN_837 : _GEN_837; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1614 = _GEN_1444 ? _GEN_838 : _GEN_838; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1615 = _GEN_1444 ? _GEN_839 : _GEN_839; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1616 = _GEN_1444 ? _GEN_840 : _GEN_840; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1617 = _GEN_1444 ? _GEN_841 : _GEN_841; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1618 = _GEN_1444 ? _GEN_842 : _GEN_842; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1619 = _GEN_1444 ? _GEN_843 : _GEN_843; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1620 = _GEN_1444 ? _GEN_844 : _GEN_844; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1621 = _GEN_1444 ? _GEN_845 : _GEN_845; // @[d_cache.scala 210:47]
  wire [31:0] _GEN_1622 = _GEN_1444 ? _GEN_846 : _GEN_846; // @[d_cache.scala 210:47]
  wire  _GEN_1623 = _GEN_1444 ? _GEN_1477 : dirty_2_0; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1624 = _GEN_1444 ? _GEN_1478 : dirty_2_1; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1625 = _GEN_1444 ? _GEN_1479 : dirty_2_2; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1626 = _GEN_1444 ? _GEN_1480 : dirty_2_3; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1627 = _GEN_1444 ? _GEN_1481 : dirty_2_4; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1628 = _GEN_1444 ? _GEN_1482 : dirty_2_5; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1629 = _GEN_1444 ? _GEN_1483 : dirty_2_6; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1630 = _GEN_1444 ? _GEN_1484 : dirty_2_7; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1631 = _GEN_1444 ? _GEN_1485 : dirty_2_8; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1632 = _GEN_1444 ? _GEN_1486 : dirty_2_9; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1633 = _GEN_1444 ? _GEN_1487 : dirty_2_10; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1634 = _GEN_1444 ? _GEN_1488 : dirty_2_11; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1635 = _GEN_1444 ? _GEN_1489 : dirty_2_12; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1636 = _GEN_1444 ? _GEN_1490 : dirty_2_13; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1637 = _GEN_1444 ? _GEN_1491 : dirty_2_14; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1638 = _GEN_1444 ? _GEN_1492 : dirty_2_15; // @[d_cache.scala 210:47 36:26]
  wire  _GEN_1639 = _GEN_1444 ? _GEN_847 : _GEN_847; // @[d_cache.scala 210:47]
  wire  _GEN_1640 = _GEN_1444 ? _GEN_848 : _GEN_848; // @[d_cache.scala 210:47]
  wire  _GEN_1641 = _GEN_1444 ? _GEN_849 : _GEN_849; // @[d_cache.scala 210:47]
  wire  _GEN_1642 = _GEN_1444 ? _GEN_850 : _GEN_850; // @[d_cache.scala 210:47]
  wire  _GEN_1643 = _GEN_1444 ? _GEN_851 : _GEN_851; // @[d_cache.scala 210:47]
  wire  _GEN_1644 = _GEN_1444 ? _GEN_852 : _GEN_852; // @[d_cache.scala 210:47]
  wire  _GEN_1645 = _GEN_1444 ? _GEN_853 : _GEN_853; // @[d_cache.scala 210:47]
  wire  _GEN_1646 = _GEN_1444 ? _GEN_854 : _GEN_854; // @[d_cache.scala 210:47]
  wire  _GEN_1647 = _GEN_1444 ? _GEN_855 : _GEN_855; // @[d_cache.scala 210:47]
  wire  _GEN_1648 = _GEN_1444 ? _GEN_856 : _GEN_856; // @[d_cache.scala 210:47]
  wire  _GEN_1649 = _GEN_1444 ? _GEN_857 : _GEN_857; // @[d_cache.scala 210:47]
  wire  _GEN_1650 = _GEN_1444 ? _GEN_858 : _GEN_858; // @[d_cache.scala 210:47]
  wire  _GEN_1651 = _GEN_1444 ? _GEN_859 : _GEN_859; // @[d_cache.scala 210:47]
  wire  _GEN_1652 = _GEN_1444 ? _GEN_860 : _GEN_860; // @[d_cache.scala 210:47]
  wire  _GEN_1653 = _GEN_1444 ? _GEN_861 : _GEN_861; // @[d_cache.scala 210:47]
  wire  _GEN_1654 = _GEN_1444 ? _GEN_862 : _GEN_862; // @[d_cache.scala 210:47]
  wire [3:0] _GEN_1655 = _GEN_1444 ? 4'h6 : 4'h1; // @[d_cache.scala 210:47 217:31 220:31]
  wire [7:0] _GEN_1656 = _GEN_1444 ? _GEN_863 : _GEN_863; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1657 = _GEN_1444 ? _GEN_864 : _GEN_864; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1658 = _GEN_1444 ? _GEN_865 : _GEN_865; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1659 = _GEN_1444 ? _GEN_866 : _GEN_866; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1660 = _GEN_1444 ? _GEN_867 : _GEN_867; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1661 = _GEN_1444 ? _GEN_868 : _GEN_868; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1662 = _GEN_1444 ? _GEN_869 : _GEN_869; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1663 = _GEN_1444 ? _GEN_870 : _GEN_870; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1664 = _GEN_1444 ? _GEN_871 : _GEN_871; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1665 = _GEN_1444 ? _GEN_872 : _GEN_872; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1666 = _GEN_1444 ? _GEN_873 : _GEN_873; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1667 = _GEN_1444 ? _GEN_874 : _GEN_874; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1668 = _GEN_1444 ? _GEN_875 : _GEN_875; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1669 = _GEN_1444 ? _GEN_876 : _GEN_876; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1670 = _GEN_1444 ? _GEN_877 : _GEN_877; // @[d_cache.scala 210:47]
  wire [7:0] _GEN_1671 = _GEN_1444 ? _GEN_878 : _GEN_878; // @[d_cache.scala 210:47]
  wire  _GEN_1673 = 4'h1 == index ? dirty_3_1 : dirty_3_0; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1674 = 4'h2 == index ? dirty_3_2 : _GEN_1673; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1675 = 4'h3 == index ? dirty_3_3 : _GEN_1674; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1676 = 4'h4 == index ? dirty_3_4 : _GEN_1675; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1677 = 4'h5 == index ? dirty_3_5 : _GEN_1676; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1678 = 4'h6 == index ? dirty_3_6 : _GEN_1677; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1679 = 4'h7 == index ? dirty_3_7 : _GEN_1678; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1680 = 4'h8 == index ? dirty_3_8 : _GEN_1679; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1681 = 4'h9 == index ? dirty_3_9 : _GEN_1680; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1682 = 4'ha == index ? dirty_3_10 : _GEN_1681; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1683 = 4'hb == index ? dirty_3_11 : _GEN_1682; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1684 = 4'hc == index ? dirty_3_12 : _GEN_1683; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1685 = 4'hd == index ? dirty_3_13 : _GEN_1684; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1686 = 4'he == index ? dirty_3_14 : _GEN_1685; // @[d_cache.scala 227:{40,40}]
  wire  _GEN_1687 = 4'hf == index ? dirty_3_15 : _GEN_1686; // @[d_cache.scala 227:{40,40}]
  wire [41:0] _write_back_addr_T_7 = {_GEN_111,index,6'h0}; // @[Cat.scala 31:58]
  wire  _GEN_1720 = 4'h0 == index ? 1'h0 : dirty_3_0; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1721 = 4'h1 == index ? 1'h0 : dirty_3_1; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1722 = 4'h2 == index ? 1'h0 : dirty_3_2; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1723 = 4'h3 == index ? 1'h0 : dirty_3_3; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1724 = 4'h4 == index ? 1'h0 : dirty_3_4; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1725 = 4'h5 == index ? 1'h0 : dirty_3_5; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1726 = 4'h6 == index ? 1'h0 : dirty_3_6; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1727 = 4'h7 == index ? 1'h0 : dirty_3_7; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1728 = 4'h8 == index ? 1'h0 : dirty_3_8; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1729 = 4'h9 == index ? 1'h0 : dirty_3_9; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1730 = 4'ha == index ? 1'h0 : dirty_3_10; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1731 = 4'hb == index ? 1'h0 : dirty_3_11; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1732 = 4'hc == index ? 1'h0 : dirty_3_12; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1733 = 4'hd == index ? 1'h0 : dirty_3_13; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1734 = 4'he == index ? 1'h0 : dirty_3_14; // @[d_cache.scala 232:{40,40} 37:26]
  wire  _GEN_1735 = 4'hf == index ? 1'h0 : dirty_3_15; // @[d_cache.scala 232:{40,40} 37:26]
  wire [511:0] _GEN_1832 = _GEN_1687 ? _GEN_294 : write_back_data; // @[d_cache.scala 227:47 228:41 44:34]
  wire [41:0] _GEN_1833 = _GEN_1687 ? _write_back_addr_T_7 : {{10'd0}, write_back_addr}; // @[d_cache.scala 227:47 229:41 45:34]
  wire [511:0] _GEN_1834 = _GEN_1687 ? _GEN_879 : _GEN_879; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1835 = _GEN_1687 ? _GEN_880 : _GEN_880; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1836 = _GEN_1687 ? _GEN_881 : _GEN_881; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1837 = _GEN_1687 ? _GEN_882 : _GEN_882; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1838 = _GEN_1687 ? _GEN_883 : _GEN_883; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1839 = _GEN_1687 ? _GEN_884 : _GEN_884; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1840 = _GEN_1687 ? _GEN_885 : _GEN_885; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1841 = _GEN_1687 ? _GEN_886 : _GEN_886; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1842 = _GEN_1687 ? _GEN_887 : _GEN_887; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1843 = _GEN_1687 ? _GEN_888 : _GEN_888; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1844 = _GEN_1687 ? _GEN_889 : _GEN_889; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1845 = _GEN_1687 ? _GEN_890 : _GEN_890; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1846 = _GEN_1687 ? _GEN_891 : _GEN_891; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1847 = _GEN_1687 ? _GEN_892 : _GEN_892; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1848 = _GEN_1687 ? _GEN_893 : _GEN_893; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1849 = _GEN_1687 ? _GEN_894 : _GEN_894; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1850 = _GEN_1687 ? _GEN_895 : _GEN_895; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1851 = _GEN_1687 ? _GEN_896 : _GEN_896; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1852 = _GEN_1687 ? _GEN_897 : _GEN_897; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1853 = _GEN_1687 ? _GEN_898 : _GEN_898; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1854 = _GEN_1687 ? _GEN_899 : _GEN_899; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1855 = _GEN_1687 ? _GEN_900 : _GEN_900; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1856 = _GEN_1687 ? _GEN_901 : _GEN_901; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1857 = _GEN_1687 ? _GEN_902 : _GEN_902; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1858 = _GEN_1687 ? _GEN_903 : _GEN_903; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1859 = _GEN_1687 ? _GEN_904 : _GEN_904; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1860 = _GEN_1687 ? _GEN_905 : _GEN_905; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1861 = _GEN_1687 ? _GEN_906 : _GEN_906; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1862 = _GEN_1687 ? _GEN_907 : _GEN_907; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1863 = _GEN_1687 ? _GEN_908 : _GEN_908; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1864 = _GEN_1687 ? _GEN_909 : _GEN_909; // @[d_cache.scala 227:47]
  wire [31:0] _GEN_1865 = _GEN_1687 ? _GEN_910 : _GEN_910; // @[d_cache.scala 227:47]
  wire  _GEN_1866 = _GEN_1687 ? _GEN_1720 : dirty_3_0; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1867 = _GEN_1687 ? _GEN_1721 : dirty_3_1; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1868 = _GEN_1687 ? _GEN_1722 : dirty_3_2; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1869 = _GEN_1687 ? _GEN_1723 : dirty_3_3; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1870 = _GEN_1687 ? _GEN_1724 : dirty_3_4; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1871 = _GEN_1687 ? _GEN_1725 : dirty_3_5; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1872 = _GEN_1687 ? _GEN_1726 : dirty_3_6; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1873 = _GEN_1687 ? _GEN_1727 : dirty_3_7; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1874 = _GEN_1687 ? _GEN_1728 : dirty_3_8; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1875 = _GEN_1687 ? _GEN_1729 : dirty_3_9; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1876 = _GEN_1687 ? _GEN_1730 : dirty_3_10; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1877 = _GEN_1687 ? _GEN_1731 : dirty_3_11; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1878 = _GEN_1687 ? _GEN_1732 : dirty_3_12; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1879 = _GEN_1687 ? _GEN_1733 : dirty_3_13; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1880 = _GEN_1687 ? _GEN_1734 : dirty_3_14; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1881 = _GEN_1687 ? _GEN_1735 : dirty_3_15; // @[d_cache.scala 227:47 37:26]
  wire  _GEN_1882 = _GEN_1687 ? _GEN_911 : _GEN_911; // @[d_cache.scala 227:47]
  wire  _GEN_1883 = _GEN_1687 ? _GEN_912 : _GEN_912; // @[d_cache.scala 227:47]
  wire  _GEN_1884 = _GEN_1687 ? _GEN_913 : _GEN_913; // @[d_cache.scala 227:47]
  wire  _GEN_1885 = _GEN_1687 ? _GEN_914 : _GEN_914; // @[d_cache.scala 227:47]
  wire  _GEN_1886 = _GEN_1687 ? _GEN_915 : _GEN_915; // @[d_cache.scala 227:47]
  wire  _GEN_1887 = _GEN_1687 ? _GEN_916 : _GEN_916; // @[d_cache.scala 227:47]
  wire  _GEN_1888 = _GEN_1687 ? _GEN_917 : _GEN_917; // @[d_cache.scala 227:47]
  wire  _GEN_1889 = _GEN_1687 ? _GEN_918 : _GEN_918; // @[d_cache.scala 227:47]
  wire  _GEN_1890 = _GEN_1687 ? _GEN_919 : _GEN_919; // @[d_cache.scala 227:47]
  wire  _GEN_1891 = _GEN_1687 ? _GEN_920 : _GEN_920; // @[d_cache.scala 227:47]
  wire  _GEN_1892 = _GEN_1687 ? _GEN_921 : _GEN_921; // @[d_cache.scala 227:47]
  wire  _GEN_1893 = _GEN_1687 ? _GEN_922 : _GEN_922; // @[d_cache.scala 227:47]
  wire  _GEN_1894 = _GEN_1687 ? _GEN_923 : _GEN_923; // @[d_cache.scala 227:47]
  wire  _GEN_1895 = _GEN_1687 ? _GEN_924 : _GEN_924; // @[d_cache.scala 227:47]
  wire  _GEN_1896 = _GEN_1687 ? _GEN_925 : _GEN_925; // @[d_cache.scala 227:47]
  wire  _GEN_1897 = _GEN_1687 ? _GEN_926 : _GEN_926; // @[d_cache.scala 227:47]
  wire [3:0] _GEN_1898 = _GEN_1687 ? 4'h6 : 4'h1; // @[d_cache.scala 227:47 234:31 237:31]
  wire [7:0] _GEN_1899 = _GEN_1687 ? _GEN_927 : _GEN_927; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1900 = _GEN_1687 ? _GEN_928 : _GEN_928; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1901 = _GEN_1687 ? _GEN_929 : _GEN_929; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1902 = _GEN_1687 ? _GEN_930 : _GEN_930; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1903 = _GEN_1687 ? _GEN_931 : _GEN_931; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1904 = _GEN_1687 ? _GEN_932 : _GEN_932; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1905 = _GEN_1687 ? _GEN_933 : _GEN_933; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1906 = _GEN_1687 ? _GEN_934 : _GEN_934; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1907 = _GEN_1687 ? _GEN_935 : _GEN_935; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1908 = _GEN_1687 ? _GEN_936 : _GEN_936; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1909 = _GEN_1687 ? _GEN_937 : _GEN_937; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1910 = _GEN_1687 ? _GEN_938 : _GEN_938; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1911 = _GEN_1687 ? _GEN_939 : _GEN_939; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1912 = _GEN_1687 ? _GEN_940 : _GEN_940; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1913 = _GEN_1687 ? _GEN_941 : _GEN_941; // @[d_cache.scala 227:47]
  wire [7:0] _GEN_1914 = _GEN_1687 ? _GEN_942 : _GEN_942; // @[d_cache.scala 227:47]
  wire [511:0] _GEN_1915 = _GEN_734[7:6] == 2'h2 ? _GEN_1589 : _GEN_1832; // @[d_cache.scala 209:52]
  wire [41:0] _GEN_1916 = _GEN_734[7:6] == 2'h2 ? _GEN_1590 : _GEN_1833; // @[d_cache.scala 209:52]
  wire [511:0] _GEN_1917 = _GEN_734[7:6] == 2'h2 ? _GEN_1591 : ram_2_0; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1918 = _GEN_734[7:6] == 2'h2 ? _GEN_1592 : ram_2_1; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1919 = _GEN_734[7:6] == 2'h2 ? _GEN_1593 : ram_2_2; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1920 = _GEN_734[7:6] == 2'h2 ? _GEN_1594 : ram_2_3; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1921 = _GEN_734[7:6] == 2'h2 ? _GEN_1595 : ram_2_4; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1922 = _GEN_734[7:6] == 2'h2 ? _GEN_1596 : ram_2_5; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1923 = _GEN_734[7:6] == 2'h2 ? _GEN_1597 : ram_2_6; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1924 = _GEN_734[7:6] == 2'h2 ? _GEN_1598 : ram_2_7; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1925 = _GEN_734[7:6] == 2'h2 ? _GEN_1599 : ram_2_8; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1926 = _GEN_734[7:6] == 2'h2 ? _GEN_1600 : ram_2_9; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1927 = _GEN_734[7:6] == 2'h2 ? _GEN_1601 : ram_2_10; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1928 = _GEN_734[7:6] == 2'h2 ? _GEN_1602 : ram_2_11; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1929 = _GEN_734[7:6] == 2'h2 ? _GEN_1603 : ram_2_12; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1930 = _GEN_734[7:6] == 2'h2 ? _GEN_1604 : ram_2_13; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1931 = _GEN_734[7:6] == 2'h2 ? _GEN_1605 : ram_2_14; // @[d_cache.scala 209:52 21:24]
  wire [511:0] _GEN_1932 = _GEN_734[7:6] == 2'h2 ? _GEN_1606 : ram_2_15; // @[d_cache.scala 209:52 21:24]
  wire [31:0] _GEN_1933 = _GEN_734[7:6] == 2'h2 ? _GEN_1607 : tag_2_0; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1934 = _GEN_734[7:6] == 2'h2 ? _GEN_1608 : tag_2_1; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1935 = _GEN_734[7:6] == 2'h2 ? _GEN_1609 : tag_2_2; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1936 = _GEN_734[7:6] == 2'h2 ? _GEN_1610 : tag_2_3; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1937 = _GEN_734[7:6] == 2'h2 ? _GEN_1611 : tag_2_4; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1938 = _GEN_734[7:6] == 2'h2 ? _GEN_1612 : tag_2_5; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1939 = _GEN_734[7:6] == 2'h2 ? _GEN_1613 : tag_2_6; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1940 = _GEN_734[7:6] == 2'h2 ? _GEN_1614 : tag_2_7; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1941 = _GEN_734[7:6] == 2'h2 ? _GEN_1615 : tag_2_8; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1942 = _GEN_734[7:6] == 2'h2 ? _GEN_1616 : tag_2_9; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1943 = _GEN_734[7:6] == 2'h2 ? _GEN_1617 : tag_2_10; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1944 = _GEN_734[7:6] == 2'h2 ? _GEN_1618 : tag_2_11; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1945 = _GEN_734[7:6] == 2'h2 ? _GEN_1619 : tag_2_12; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1946 = _GEN_734[7:6] == 2'h2 ? _GEN_1620 : tag_2_13; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1947 = _GEN_734[7:6] == 2'h2 ? _GEN_1621 : tag_2_14; // @[d_cache.scala 209:52 26:24]
  wire [31:0] _GEN_1948 = _GEN_734[7:6] == 2'h2 ? _GEN_1622 : tag_2_15; // @[d_cache.scala 209:52 26:24]
  wire  _GEN_1949 = _GEN_734[7:6] == 2'h2 ? _GEN_1623 : dirty_2_0; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1950 = _GEN_734[7:6] == 2'h2 ? _GEN_1624 : dirty_2_1; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1951 = _GEN_734[7:6] == 2'h2 ? _GEN_1625 : dirty_2_2; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1952 = _GEN_734[7:6] == 2'h2 ? _GEN_1626 : dirty_2_3; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1953 = _GEN_734[7:6] == 2'h2 ? _GEN_1627 : dirty_2_4; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1954 = _GEN_734[7:6] == 2'h2 ? _GEN_1628 : dirty_2_5; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1955 = _GEN_734[7:6] == 2'h2 ? _GEN_1629 : dirty_2_6; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1956 = _GEN_734[7:6] == 2'h2 ? _GEN_1630 : dirty_2_7; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1957 = _GEN_734[7:6] == 2'h2 ? _GEN_1631 : dirty_2_8; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1958 = _GEN_734[7:6] == 2'h2 ? _GEN_1632 : dirty_2_9; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1959 = _GEN_734[7:6] == 2'h2 ? _GEN_1633 : dirty_2_10; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1960 = _GEN_734[7:6] == 2'h2 ? _GEN_1634 : dirty_2_11; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1961 = _GEN_734[7:6] == 2'h2 ? _GEN_1635 : dirty_2_12; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1962 = _GEN_734[7:6] == 2'h2 ? _GEN_1636 : dirty_2_13; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1963 = _GEN_734[7:6] == 2'h2 ? _GEN_1637 : dirty_2_14; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1964 = _GEN_734[7:6] == 2'h2 ? _GEN_1638 : dirty_2_15; // @[d_cache.scala 209:52 36:26]
  wire  _GEN_1965 = _GEN_734[7:6] == 2'h2 ? _GEN_1639 : valid_2_0; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1966 = _GEN_734[7:6] == 2'h2 ? _GEN_1640 : valid_2_1; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1967 = _GEN_734[7:6] == 2'h2 ? _GEN_1641 : valid_2_2; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1968 = _GEN_734[7:6] == 2'h2 ? _GEN_1642 : valid_2_3; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1969 = _GEN_734[7:6] == 2'h2 ? _GEN_1643 : valid_2_4; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1970 = _GEN_734[7:6] == 2'h2 ? _GEN_1644 : valid_2_5; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1971 = _GEN_734[7:6] == 2'h2 ? _GEN_1645 : valid_2_6; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1972 = _GEN_734[7:6] == 2'h2 ? _GEN_1646 : valid_2_7; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1973 = _GEN_734[7:6] == 2'h2 ? _GEN_1647 : valid_2_8; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1974 = _GEN_734[7:6] == 2'h2 ? _GEN_1648 : valid_2_9; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1975 = _GEN_734[7:6] == 2'h2 ? _GEN_1649 : valid_2_10; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1976 = _GEN_734[7:6] == 2'h2 ? _GEN_1650 : valid_2_11; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1977 = _GEN_734[7:6] == 2'h2 ? _GEN_1651 : valid_2_12; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1978 = _GEN_734[7:6] == 2'h2 ? _GEN_1652 : valid_2_13; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1979 = _GEN_734[7:6] == 2'h2 ? _GEN_1653 : valid_2_14; // @[d_cache.scala 209:52 31:26]
  wire  _GEN_1980 = _GEN_734[7:6] == 2'h2 ? _GEN_1654 : valid_2_15; // @[d_cache.scala 209:52 31:26]
  wire [3:0] _GEN_1981 = _GEN_734[7:6] == 2'h2 ? _GEN_1655 : _GEN_1898; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1982 = _GEN_734[7:6] == 2'h2 ? _GEN_1656 : _GEN_1899; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1983 = _GEN_734[7:6] == 2'h2 ? _GEN_1657 : _GEN_1900; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1984 = _GEN_734[7:6] == 2'h2 ? _GEN_1658 : _GEN_1901; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1985 = _GEN_734[7:6] == 2'h2 ? _GEN_1659 : _GEN_1902; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1986 = _GEN_734[7:6] == 2'h2 ? _GEN_1660 : _GEN_1903; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1987 = _GEN_734[7:6] == 2'h2 ? _GEN_1661 : _GEN_1904; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1988 = _GEN_734[7:6] == 2'h2 ? _GEN_1662 : _GEN_1905; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1989 = _GEN_734[7:6] == 2'h2 ? _GEN_1663 : _GEN_1906; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1990 = _GEN_734[7:6] == 2'h2 ? _GEN_1664 : _GEN_1907; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1991 = _GEN_734[7:6] == 2'h2 ? _GEN_1665 : _GEN_1908; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1992 = _GEN_734[7:6] == 2'h2 ? _GEN_1666 : _GEN_1909; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1993 = _GEN_734[7:6] == 2'h2 ? _GEN_1667 : _GEN_1910; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1994 = _GEN_734[7:6] == 2'h2 ? _GEN_1668 : _GEN_1911; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1995 = _GEN_734[7:6] == 2'h2 ? _GEN_1669 : _GEN_1912; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1996 = _GEN_734[7:6] == 2'h2 ? _GEN_1670 : _GEN_1913; // @[d_cache.scala 209:52]
  wire [7:0] _GEN_1997 = _GEN_734[7:6] == 2'h2 ? _GEN_1671 : _GEN_1914; // @[d_cache.scala 209:52]
  wire [511:0] _GEN_1998 = _GEN_734[7:6] == 2'h2 ? ram_3_0 : _GEN_1834; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_1999 = _GEN_734[7:6] == 2'h2 ? ram_3_1 : _GEN_1835; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2000 = _GEN_734[7:6] == 2'h2 ? ram_3_2 : _GEN_1836; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2001 = _GEN_734[7:6] == 2'h2 ? ram_3_3 : _GEN_1837; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2002 = _GEN_734[7:6] == 2'h2 ? ram_3_4 : _GEN_1838; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2003 = _GEN_734[7:6] == 2'h2 ? ram_3_5 : _GEN_1839; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2004 = _GEN_734[7:6] == 2'h2 ? ram_3_6 : _GEN_1840; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2005 = _GEN_734[7:6] == 2'h2 ? ram_3_7 : _GEN_1841; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2006 = _GEN_734[7:6] == 2'h2 ? ram_3_8 : _GEN_1842; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2007 = _GEN_734[7:6] == 2'h2 ? ram_3_9 : _GEN_1843; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2008 = _GEN_734[7:6] == 2'h2 ? ram_3_10 : _GEN_1844; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2009 = _GEN_734[7:6] == 2'h2 ? ram_3_11 : _GEN_1845; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2010 = _GEN_734[7:6] == 2'h2 ? ram_3_12 : _GEN_1846; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2011 = _GEN_734[7:6] == 2'h2 ? ram_3_13 : _GEN_1847; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2012 = _GEN_734[7:6] == 2'h2 ? ram_3_14 : _GEN_1848; // @[d_cache.scala 209:52 22:24]
  wire [511:0] _GEN_2013 = _GEN_734[7:6] == 2'h2 ? ram_3_15 : _GEN_1849; // @[d_cache.scala 209:52 22:24]
  wire [31:0] _GEN_2014 = _GEN_734[7:6] == 2'h2 ? tag_3_0 : _GEN_1850; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2015 = _GEN_734[7:6] == 2'h2 ? tag_3_1 : _GEN_1851; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2016 = _GEN_734[7:6] == 2'h2 ? tag_3_2 : _GEN_1852; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2017 = _GEN_734[7:6] == 2'h2 ? tag_3_3 : _GEN_1853; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2018 = _GEN_734[7:6] == 2'h2 ? tag_3_4 : _GEN_1854; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2019 = _GEN_734[7:6] == 2'h2 ? tag_3_5 : _GEN_1855; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2020 = _GEN_734[7:6] == 2'h2 ? tag_3_6 : _GEN_1856; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2021 = _GEN_734[7:6] == 2'h2 ? tag_3_7 : _GEN_1857; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2022 = _GEN_734[7:6] == 2'h2 ? tag_3_8 : _GEN_1858; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2023 = _GEN_734[7:6] == 2'h2 ? tag_3_9 : _GEN_1859; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2024 = _GEN_734[7:6] == 2'h2 ? tag_3_10 : _GEN_1860; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2025 = _GEN_734[7:6] == 2'h2 ? tag_3_11 : _GEN_1861; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2026 = _GEN_734[7:6] == 2'h2 ? tag_3_12 : _GEN_1862; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2027 = _GEN_734[7:6] == 2'h2 ? tag_3_13 : _GEN_1863; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2028 = _GEN_734[7:6] == 2'h2 ? tag_3_14 : _GEN_1864; // @[d_cache.scala 209:52 27:24]
  wire [31:0] _GEN_2029 = _GEN_734[7:6] == 2'h2 ? tag_3_15 : _GEN_1865; // @[d_cache.scala 209:52 27:24]
  wire  _GEN_2030 = _GEN_734[7:6] == 2'h2 ? dirty_3_0 : _GEN_1866; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2031 = _GEN_734[7:6] == 2'h2 ? dirty_3_1 : _GEN_1867; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2032 = _GEN_734[7:6] == 2'h2 ? dirty_3_2 : _GEN_1868; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2033 = _GEN_734[7:6] == 2'h2 ? dirty_3_3 : _GEN_1869; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2034 = _GEN_734[7:6] == 2'h2 ? dirty_3_4 : _GEN_1870; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2035 = _GEN_734[7:6] == 2'h2 ? dirty_3_5 : _GEN_1871; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2036 = _GEN_734[7:6] == 2'h2 ? dirty_3_6 : _GEN_1872; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2037 = _GEN_734[7:6] == 2'h2 ? dirty_3_7 : _GEN_1873; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2038 = _GEN_734[7:6] == 2'h2 ? dirty_3_8 : _GEN_1874; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2039 = _GEN_734[7:6] == 2'h2 ? dirty_3_9 : _GEN_1875; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2040 = _GEN_734[7:6] == 2'h2 ? dirty_3_10 : _GEN_1876; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2041 = _GEN_734[7:6] == 2'h2 ? dirty_3_11 : _GEN_1877; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2042 = _GEN_734[7:6] == 2'h2 ? dirty_3_12 : _GEN_1878; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2043 = _GEN_734[7:6] == 2'h2 ? dirty_3_13 : _GEN_1879; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2044 = _GEN_734[7:6] == 2'h2 ? dirty_3_14 : _GEN_1880; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2045 = _GEN_734[7:6] == 2'h2 ? dirty_3_15 : _GEN_1881; // @[d_cache.scala 209:52 37:26]
  wire  _GEN_2046 = _GEN_734[7:6] == 2'h2 ? valid_3_0 : _GEN_1882; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2047 = _GEN_734[7:6] == 2'h2 ? valid_3_1 : _GEN_1883; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2048 = _GEN_734[7:6] == 2'h2 ? valid_3_2 : _GEN_1884; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2049 = _GEN_734[7:6] == 2'h2 ? valid_3_3 : _GEN_1885; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2050 = _GEN_734[7:6] == 2'h2 ? valid_3_4 : _GEN_1886; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2051 = _GEN_734[7:6] == 2'h2 ? valid_3_5 : _GEN_1887; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2052 = _GEN_734[7:6] == 2'h2 ? valid_3_6 : _GEN_1888; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2053 = _GEN_734[7:6] == 2'h2 ? valid_3_7 : _GEN_1889; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2054 = _GEN_734[7:6] == 2'h2 ? valid_3_8 : _GEN_1890; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2055 = _GEN_734[7:6] == 2'h2 ? valid_3_9 : _GEN_1891; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2056 = _GEN_734[7:6] == 2'h2 ? valid_3_10 : _GEN_1892; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2057 = _GEN_734[7:6] == 2'h2 ? valid_3_11 : _GEN_1893; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2058 = _GEN_734[7:6] == 2'h2 ? valid_3_12 : _GEN_1894; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2059 = _GEN_734[7:6] == 2'h2 ? valid_3_13 : _GEN_1895; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2060 = _GEN_734[7:6] == 2'h2 ? valid_3_14 : _GEN_1896; // @[d_cache.scala 209:52 32:26]
  wire  _GEN_2061 = _GEN_734[7:6] == 2'h2 ? valid_3_15 : _GEN_1897; // @[d_cache.scala 209:52 32:26]
  wire [511:0] _GEN_2062 = _GEN_734[7:6] == 2'h1 ? _GEN_1346 : _GEN_1915; // @[d_cache.scala 192:52]
  wire [41:0] _GEN_2063 = _GEN_734[7:6] == 2'h1 ? _GEN_1347 : _GEN_1916; // @[d_cache.scala 192:52]
  wire [511:0] _GEN_2064 = _GEN_734[7:6] == 2'h1 ? _GEN_1348 : ram_1_0; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2065 = _GEN_734[7:6] == 2'h1 ? _GEN_1349 : ram_1_1; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2066 = _GEN_734[7:6] == 2'h1 ? _GEN_1350 : ram_1_2; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2067 = _GEN_734[7:6] == 2'h1 ? _GEN_1351 : ram_1_3; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2068 = _GEN_734[7:6] == 2'h1 ? _GEN_1352 : ram_1_4; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2069 = _GEN_734[7:6] == 2'h1 ? _GEN_1353 : ram_1_5; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2070 = _GEN_734[7:6] == 2'h1 ? _GEN_1354 : ram_1_6; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2071 = _GEN_734[7:6] == 2'h1 ? _GEN_1355 : ram_1_7; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2072 = _GEN_734[7:6] == 2'h1 ? _GEN_1356 : ram_1_8; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2073 = _GEN_734[7:6] == 2'h1 ? _GEN_1357 : ram_1_9; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2074 = _GEN_734[7:6] == 2'h1 ? _GEN_1358 : ram_1_10; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2075 = _GEN_734[7:6] == 2'h1 ? _GEN_1359 : ram_1_11; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2076 = _GEN_734[7:6] == 2'h1 ? _GEN_1360 : ram_1_12; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2077 = _GEN_734[7:6] == 2'h1 ? _GEN_1361 : ram_1_13; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2078 = _GEN_734[7:6] == 2'h1 ? _GEN_1362 : ram_1_14; // @[d_cache.scala 192:52 20:24]
  wire [511:0] _GEN_2079 = _GEN_734[7:6] == 2'h1 ? _GEN_1363 : ram_1_15; // @[d_cache.scala 192:52 20:24]
  wire [31:0] _GEN_2080 = _GEN_734[7:6] == 2'h1 ? _GEN_1364 : tag_1_0; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2081 = _GEN_734[7:6] == 2'h1 ? _GEN_1365 : tag_1_1; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2082 = _GEN_734[7:6] == 2'h1 ? _GEN_1366 : tag_1_2; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2083 = _GEN_734[7:6] == 2'h1 ? _GEN_1367 : tag_1_3; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2084 = _GEN_734[7:6] == 2'h1 ? _GEN_1368 : tag_1_4; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2085 = _GEN_734[7:6] == 2'h1 ? _GEN_1369 : tag_1_5; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2086 = _GEN_734[7:6] == 2'h1 ? _GEN_1370 : tag_1_6; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2087 = _GEN_734[7:6] == 2'h1 ? _GEN_1371 : tag_1_7; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2088 = _GEN_734[7:6] == 2'h1 ? _GEN_1372 : tag_1_8; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2089 = _GEN_734[7:6] == 2'h1 ? _GEN_1373 : tag_1_9; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2090 = _GEN_734[7:6] == 2'h1 ? _GEN_1374 : tag_1_10; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2091 = _GEN_734[7:6] == 2'h1 ? _GEN_1375 : tag_1_11; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2092 = _GEN_734[7:6] == 2'h1 ? _GEN_1376 : tag_1_12; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2093 = _GEN_734[7:6] == 2'h1 ? _GEN_1377 : tag_1_13; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2094 = _GEN_734[7:6] == 2'h1 ? _GEN_1378 : tag_1_14; // @[d_cache.scala 192:52 25:24]
  wire [31:0] _GEN_2095 = _GEN_734[7:6] == 2'h1 ? _GEN_1379 : tag_1_15; // @[d_cache.scala 192:52 25:24]
  wire  _GEN_2096 = _GEN_734[7:6] == 2'h1 ? _GEN_1380 : dirty_1_0; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2097 = _GEN_734[7:6] == 2'h1 ? _GEN_1381 : dirty_1_1; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2098 = _GEN_734[7:6] == 2'h1 ? _GEN_1382 : dirty_1_2; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2099 = _GEN_734[7:6] == 2'h1 ? _GEN_1383 : dirty_1_3; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2100 = _GEN_734[7:6] == 2'h1 ? _GEN_1384 : dirty_1_4; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2101 = _GEN_734[7:6] == 2'h1 ? _GEN_1385 : dirty_1_5; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2102 = _GEN_734[7:6] == 2'h1 ? _GEN_1386 : dirty_1_6; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2103 = _GEN_734[7:6] == 2'h1 ? _GEN_1387 : dirty_1_7; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2104 = _GEN_734[7:6] == 2'h1 ? _GEN_1388 : dirty_1_8; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2105 = _GEN_734[7:6] == 2'h1 ? _GEN_1389 : dirty_1_9; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2106 = _GEN_734[7:6] == 2'h1 ? _GEN_1390 : dirty_1_10; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2107 = _GEN_734[7:6] == 2'h1 ? _GEN_1391 : dirty_1_11; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2108 = _GEN_734[7:6] == 2'h1 ? _GEN_1392 : dirty_1_12; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2109 = _GEN_734[7:6] == 2'h1 ? _GEN_1393 : dirty_1_13; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2110 = _GEN_734[7:6] == 2'h1 ? _GEN_1394 : dirty_1_14; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2111 = _GEN_734[7:6] == 2'h1 ? _GEN_1395 : dirty_1_15; // @[d_cache.scala 192:52 35:26]
  wire  _GEN_2112 = _GEN_734[7:6] == 2'h1 ? _GEN_1396 : valid_1_0; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2113 = _GEN_734[7:6] == 2'h1 ? _GEN_1397 : valid_1_1; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2114 = _GEN_734[7:6] == 2'h1 ? _GEN_1398 : valid_1_2; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2115 = _GEN_734[7:6] == 2'h1 ? _GEN_1399 : valid_1_3; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2116 = _GEN_734[7:6] == 2'h1 ? _GEN_1400 : valid_1_4; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2117 = _GEN_734[7:6] == 2'h1 ? _GEN_1401 : valid_1_5; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2118 = _GEN_734[7:6] == 2'h1 ? _GEN_1402 : valid_1_6; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2119 = _GEN_734[7:6] == 2'h1 ? _GEN_1403 : valid_1_7; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2120 = _GEN_734[7:6] == 2'h1 ? _GEN_1404 : valid_1_8; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2121 = _GEN_734[7:6] == 2'h1 ? _GEN_1405 : valid_1_9; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2122 = _GEN_734[7:6] == 2'h1 ? _GEN_1406 : valid_1_10; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2123 = _GEN_734[7:6] == 2'h1 ? _GEN_1407 : valid_1_11; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2124 = _GEN_734[7:6] == 2'h1 ? _GEN_1408 : valid_1_12; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2125 = _GEN_734[7:6] == 2'h1 ? _GEN_1409 : valid_1_13; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2126 = _GEN_734[7:6] == 2'h1 ? _GEN_1410 : valid_1_14; // @[d_cache.scala 192:52 30:26]
  wire  _GEN_2127 = _GEN_734[7:6] == 2'h1 ? _GEN_1411 : valid_1_15; // @[d_cache.scala 192:52 30:26]
  wire [3:0] _GEN_2128 = _GEN_734[7:6] == 2'h1 ? _GEN_1412 : _GEN_1981; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2129 = _GEN_734[7:6] == 2'h1 ? _GEN_1413 : _GEN_1982; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2130 = _GEN_734[7:6] == 2'h1 ? _GEN_1414 : _GEN_1983; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2131 = _GEN_734[7:6] == 2'h1 ? _GEN_1415 : _GEN_1984; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2132 = _GEN_734[7:6] == 2'h1 ? _GEN_1416 : _GEN_1985; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2133 = _GEN_734[7:6] == 2'h1 ? _GEN_1417 : _GEN_1986; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2134 = _GEN_734[7:6] == 2'h1 ? _GEN_1418 : _GEN_1987; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2135 = _GEN_734[7:6] == 2'h1 ? _GEN_1419 : _GEN_1988; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2136 = _GEN_734[7:6] == 2'h1 ? _GEN_1420 : _GEN_1989; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2137 = _GEN_734[7:6] == 2'h1 ? _GEN_1421 : _GEN_1990; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2138 = _GEN_734[7:6] == 2'h1 ? _GEN_1422 : _GEN_1991; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2139 = _GEN_734[7:6] == 2'h1 ? _GEN_1423 : _GEN_1992; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2140 = _GEN_734[7:6] == 2'h1 ? _GEN_1424 : _GEN_1993; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2141 = _GEN_734[7:6] == 2'h1 ? _GEN_1425 : _GEN_1994; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2142 = _GEN_734[7:6] == 2'h1 ? _GEN_1426 : _GEN_1995; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2143 = _GEN_734[7:6] == 2'h1 ? _GEN_1427 : _GEN_1996; // @[d_cache.scala 192:52]
  wire [7:0] _GEN_2144 = _GEN_734[7:6] == 2'h1 ? _GEN_1428 : _GEN_1997; // @[d_cache.scala 192:52]
  wire [511:0] _GEN_2145 = _GEN_734[7:6] == 2'h1 ? ram_2_0 : _GEN_1917; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2146 = _GEN_734[7:6] == 2'h1 ? ram_2_1 : _GEN_1918; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2147 = _GEN_734[7:6] == 2'h1 ? ram_2_2 : _GEN_1919; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2148 = _GEN_734[7:6] == 2'h1 ? ram_2_3 : _GEN_1920; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2149 = _GEN_734[7:6] == 2'h1 ? ram_2_4 : _GEN_1921; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2150 = _GEN_734[7:6] == 2'h1 ? ram_2_5 : _GEN_1922; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2151 = _GEN_734[7:6] == 2'h1 ? ram_2_6 : _GEN_1923; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2152 = _GEN_734[7:6] == 2'h1 ? ram_2_7 : _GEN_1924; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2153 = _GEN_734[7:6] == 2'h1 ? ram_2_8 : _GEN_1925; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2154 = _GEN_734[7:6] == 2'h1 ? ram_2_9 : _GEN_1926; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2155 = _GEN_734[7:6] == 2'h1 ? ram_2_10 : _GEN_1927; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2156 = _GEN_734[7:6] == 2'h1 ? ram_2_11 : _GEN_1928; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2157 = _GEN_734[7:6] == 2'h1 ? ram_2_12 : _GEN_1929; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2158 = _GEN_734[7:6] == 2'h1 ? ram_2_13 : _GEN_1930; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2159 = _GEN_734[7:6] == 2'h1 ? ram_2_14 : _GEN_1931; // @[d_cache.scala 192:52 21:24]
  wire [511:0] _GEN_2160 = _GEN_734[7:6] == 2'h1 ? ram_2_15 : _GEN_1932; // @[d_cache.scala 192:52 21:24]
  wire [31:0] _GEN_2161 = _GEN_734[7:6] == 2'h1 ? tag_2_0 : _GEN_1933; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2162 = _GEN_734[7:6] == 2'h1 ? tag_2_1 : _GEN_1934; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2163 = _GEN_734[7:6] == 2'h1 ? tag_2_2 : _GEN_1935; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2164 = _GEN_734[7:6] == 2'h1 ? tag_2_3 : _GEN_1936; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2165 = _GEN_734[7:6] == 2'h1 ? tag_2_4 : _GEN_1937; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2166 = _GEN_734[7:6] == 2'h1 ? tag_2_5 : _GEN_1938; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2167 = _GEN_734[7:6] == 2'h1 ? tag_2_6 : _GEN_1939; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2168 = _GEN_734[7:6] == 2'h1 ? tag_2_7 : _GEN_1940; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2169 = _GEN_734[7:6] == 2'h1 ? tag_2_8 : _GEN_1941; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2170 = _GEN_734[7:6] == 2'h1 ? tag_2_9 : _GEN_1942; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2171 = _GEN_734[7:6] == 2'h1 ? tag_2_10 : _GEN_1943; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2172 = _GEN_734[7:6] == 2'h1 ? tag_2_11 : _GEN_1944; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2173 = _GEN_734[7:6] == 2'h1 ? tag_2_12 : _GEN_1945; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2174 = _GEN_734[7:6] == 2'h1 ? tag_2_13 : _GEN_1946; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2175 = _GEN_734[7:6] == 2'h1 ? tag_2_14 : _GEN_1947; // @[d_cache.scala 192:52 26:24]
  wire [31:0] _GEN_2176 = _GEN_734[7:6] == 2'h1 ? tag_2_15 : _GEN_1948; // @[d_cache.scala 192:52 26:24]
  wire  _GEN_2177 = _GEN_734[7:6] == 2'h1 ? dirty_2_0 : _GEN_1949; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2178 = _GEN_734[7:6] == 2'h1 ? dirty_2_1 : _GEN_1950; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2179 = _GEN_734[7:6] == 2'h1 ? dirty_2_2 : _GEN_1951; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2180 = _GEN_734[7:6] == 2'h1 ? dirty_2_3 : _GEN_1952; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2181 = _GEN_734[7:6] == 2'h1 ? dirty_2_4 : _GEN_1953; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2182 = _GEN_734[7:6] == 2'h1 ? dirty_2_5 : _GEN_1954; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2183 = _GEN_734[7:6] == 2'h1 ? dirty_2_6 : _GEN_1955; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2184 = _GEN_734[7:6] == 2'h1 ? dirty_2_7 : _GEN_1956; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2185 = _GEN_734[7:6] == 2'h1 ? dirty_2_8 : _GEN_1957; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2186 = _GEN_734[7:6] == 2'h1 ? dirty_2_9 : _GEN_1958; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2187 = _GEN_734[7:6] == 2'h1 ? dirty_2_10 : _GEN_1959; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2188 = _GEN_734[7:6] == 2'h1 ? dirty_2_11 : _GEN_1960; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2189 = _GEN_734[7:6] == 2'h1 ? dirty_2_12 : _GEN_1961; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2190 = _GEN_734[7:6] == 2'h1 ? dirty_2_13 : _GEN_1962; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2191 = _GEN_734[7:6] == 2'h1 ? dirty_2_14 : _GEN_1963; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2192 = _GEN_734[7:6] == 2'h1 ? dirty_2_15 : _GEN_1964; // @[d_cache.scala 192:52 36:26]
  wire  _GEN_2193 = _GEN_734[7:6] == 2'h1 ? valid_2_0 : _GEN_1965; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2194 = _GEN_734[7:6] == 2'h1 ? valid_2_1 : _GEN_1966; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2195 = _GEN_734[7:6] == 2'h1 ? valid_2_2 : _GEN_1967; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2196 = _GEN_734[7:6] == 2'h1 ? valid_2_3 : _GEN_1968; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2197 = _GEN_734[7:6] == 2'h1 ? valid_2_4 : _GEN_1969; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2198 = _GEN_734[7:6] == 2'h1 ? valid_2_5 : _GEN_1970; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2199 = _GEN_734[7:6] == 2'h1 ? valid_2_6 : _GEN_1971; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2200 = _GEN_734[7:6] == 2'h1 ? valid_2_7 : _GEN_1972; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2201 = _GEN_734[7:6] == 2'h1 ? valid_2_8 : _GEN_1973; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2202 = _GEN_734[7:6] == 2'h1 ? valid_2_9 : _GEN_1974; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2203 = _GEN_734[7:6] == 2'h1 ? valid_2_10 : _GEN_1975; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2204 = _GEN_734[7:6] == 2'h1 ? valid_2_11 : _GEN_1976; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2205 = _GEN_734[7:6] == 2'h1 ? valid_2_12 : _GEN_1977; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2206 = _GEN_734[7:6] == 2'h1 ? valid_2_13 : _GEN_1978; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2207 = _GEN_734[7:6] == 2'h1 ? valid_2_14 : _GEN_1979; // @[d_cache.scala 192:52 31:26]
  wire  _GEN_2208 = _GEN_734[7:6] == 2'h1 ? valid_2_15 : _GEN_1980; // @[d_cache.scala 192:52 31:26]
  wire [511:0] _GEN_2209 = _GEN_734[7:6] == 2'h1 ? ram_3_0 : _GEN_1998; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2210 = _GEN_734[7:6] == 2'h1 ? ram_3_1 : _GEN_1999; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2211 = _GEN_734[7:6] == 2'h1 ? ram_3_2 : _GEN_2000; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2212 = _GEN_734[7:6] == 2'h1 ? ram_3_3 : _GEN_2001; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2213 = _GEN_734[7:6] == 2'h1 ? ram_3_4 : _GEN_2002; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2214 = _GEN_734[7:6] == 2'h1 ? ram_3_5 : _GEN_2003; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2215 = _GEN_734[7:6] == 2'h1 ? ram_3_6 : _GEN_2004; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2216 = _GEN_734[7:6] == 2'h1 ? ram_3_7 : _GEN_2005; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2217 = _GEN_734[7:6] == 2'h1 ? ram_3_8 : _GEN_2006; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2218 = _GEN_734[7:6] == 2'h1 ? ram_3_9 : _GEN_2007; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2219 = _GEN_734[7:6] == 2'h1 ? ram_3_10 : _GEN_2008; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2220 = _GEN_734[7:6] == 2'h1 ? ram_3_11 : _GEN_2009; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2221 = _GEN_734[7:6] == 2'h1 ? ram_3_12 : _GEN_2010; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2222 = _GEN_734[7:6] == 2'h1 ? ram_3_13 : _GEN_2011; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2223 = _GEN_734[7:6] == 2'h1 ? ram_3_14 : _GEN_2012; // @[d_cache.scala 192:52 22:24]
  wire [511:0] _GEN_2224 = _GEN_734[7:6] == 2'h1 ? ram_3_15 : _GEN_2013; // @[d_cache.scala 192:52 22:24]
  wire [31:0] _GEN_2225 = _GEN_734[7:6] == 2'h1 ? tag_3_0 : _GEN_2014; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2226 = _GEN_734[7:6] == 2'h1 ? tag_3_1 : _GEN_2015; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2227 = _GEN_734[7:6] == 2'h1 ? tag_3_2 : _GEN_2016; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2228 = _GEN_734[7:6] == 2'h1 ? tag_3_3 : _GEN_2017; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2229 = _GEN_734[7:6] == 2'h1 ? tag_3_4 : _GEN_2018; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2230 = _GEN_734[7:6] == 2'h1 ? tag_3_5 : _GEN_2019; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2231 = _GEN_734[7:6] == 2'h1 ? tag_3_6 : _GEN_2020; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2232 = _GEN_734[7:6] == 2'h1 ? tag_3_7 : _GEN_2021; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2233 = _GEN_734[7:6] == 2'h1 ? tag_3_8 : _GEN_2022; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2234 = _GEN_734[7:6] == 2'h1 ? tag_3_9 : _GEN_2023; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2235 = _GEN_734[7:6] == 2'h1 ? tag_3_10 : _GEN_2024; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2236 = _GEN_734[7:6] == 2'h1 ? tag_3_11 : _GEN_2025; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2237 = _GEN_734[7:6] == 2'h1 ? tag_3_12 : _GEN_2026; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2238 = _GEN_734[7:6] == 2'h1 ? tag_3_13 : _GEN_2027; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2239 = _GEN_734[7:6] == 2'h1 ? tag_3_14 : _GEN_2028; // @[d_cache.scala 192:52 27:24]
  wire [31:0] _GEN_2240 = _GEN_734[7:6] == 2'h1 ? tag_3_15 : _GEN_2029; // @[d_cache.scala 192:52 27:24]
  wire  _GEN_2241 = _GEN_734[7:6] == 2'h1 ? dirty_3_0 : _GEN_2030; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2242 = _GEN_734[7:6] == 2'h1 ? dirty_3_1 : _GEN_2031; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2243 = _GEN_734[7:6] == 2'h1 ? dirty_3_2 : _GEN_2032; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2244 = _GEN_734[7:6] == 2'h1 ? dirty_3_3 : _GEN_2033; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2245 = _GEN_734[7:6] == 2'h1 ? dirty_3_4 : _GEN_2034; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2246 = _GEN_734[7:6] == 2'h1 ? dirty_3_5 : _GEN_2035; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2247 = _GEN_734[7:6] == 2'h1 ? dirty_3_6 : _GEN_2036; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2248 = _GEN_734[7:6] == 2'h1 ? dirty_3_7 : _GEN_2037; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2249 = _GEN_734[7:6] == 2'h1 ? dirty_3_8 : _GEN_2038; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2250 = _GEN_734[7:6] == 2'h1 ? dirty_3_9 : _GEN_2039; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2251 = _GEN_734[7:6] == 2'h1 ? dirty_3_10 : _GEN_2040; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2252 = _GEN_734[7:6] == 2'h1 ? dirty_3_11 : _GEN_2041; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2253 = _GEN_734[7:6] == 2'h1 ? dirty_3_12 : _GEN_2042; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2254 = _GEN_734[7:6] == 2'h1 ? dirty_3_13 : _GEN_2043; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2255 = _GEN_734[7:6] == 2'h1 ? dirty_3_14 : _GEN_2044; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2256 = _GEN_734[7:6] == 2'h1 ? dirty_3_15 : _GEN_2045; // @[d_cache.scala 192:52 37:26]
  wire  _GEN_2257 = _GEN_734[7:6] == 2'h1 ? valid_3_0 : _GEN_2046; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2258 = _GEN_734[7:6] == 2'h1 ? valid_3_1 : _GEN_2047; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2259 = _GEN_734[7:6] == 2'h1 ? valid_3_2 : _GEN_2048; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2260 = _GEN_734[7:6] == 2'h1 ? valid_3_3 : _GEN_2049; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2261 = _GEN_734[7:6] == 2'h1 ? valid_3_4 : _GEN_2050; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2262 = _GEN_734[7:6] == 2'h1 ? valid_3_5 : _GEN_2051; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2263 = _GEN_734[7:6] == 2'h1 ? valid_3_6 : _GEN_2052; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2264 = _GEN_734[7:6] == 2'h1 ? valid_3_7 : _GEN_2053; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2265 = _GEN_734[7:6] == 2'h1 ? valid_3_8 : _GEN_2054; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2266 = _GEN_734[7:6] == 2'h1 ? valid_3_9 : _GEN_2055; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2267 = _GEN_734[7:6] == 2'h1 ? valid_3_10 : _GEN_2056; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2268 = _GEN_734[7:6] == 2'h1 ? valid_3_11 : _GEN_2057; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2269 = _GEN_734[7:6] == 2'h1 ? valid_3_12 : _GEN_2058; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2270 = _GEN_734[7:6] == 2'h1 ? valid_3_13 : _GEN_2059; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2271 = _GEN_734[7:6] == 2'h1 ? valid_3_14 : _GEN_2060; // @[d_cache.scala 192:52 32:26]
  wire  _GEN_2272 = _GEN_734[7:6] == 2'h1 ? valid_3_15 : _GEN_2061; // @[d_cache.scala 192:52 32:26]
  wire [511:0] _GEN_2273 = _GEN_734[7:6] == 2'h0 ? _GEN_1103 : _GEN_2062; // @[d_cache.scala 175:46]
  wire [41:0] _GEN_2274 = _GEN_734[7:6] == 2'h0 ? _GEN_1104 : _GEN_2063; // @[d_cache.scala 175:46]
  wire [511:0] _GEN_2275 = _GEN_734[7:6] == 2'h0 ? _GEN_1105 : ram_0_0; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2276 = _GEN_734[7:6] == 2'h0 ? _GEN_1106 : ram_0_1; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2277 = _GEN_734[7:6] == 2'h0 ? _GEN_1107 : ram_0_2; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2278 = _GEN_734[7:6] == 2'h0 ? _GEN_1108 : ram_0_3; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2279 = _GEN_734[7:6] == 2'h0 ? _GEN_1109 : ram_0_4; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2280 = _GEN_734[7:6] == 2'h0 ? _GEN_1110 : ram_0_5; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2281 = _GEN_734[7:6] == 2'h0 ? _GEN_1111 : ram_0_6; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2282 = _GEN_734[7:6] == 2'h0 ? _GEN_1112 : ram_0_7; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2283 = _GEN_734[7:6] == 2'h0 ? _GEN_1113 : ram_0_8; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2284 = _GEN_734[7:6] == 2'h0 ? _GEN_1114 : ram_0_9; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2285 = _GEN_734[7:6] == 2'h0 ? _GEN_1115 : ram_0_10; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2286 = _GEN_734[7:6] == 2'h0 ? _GEN_1116 : ram_0_11; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2287 = _GEN_734[7:6] == 2'h0 ? _GEN_1117 : ram_0_12; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2288 = _GEN_734[7:6] == 2'h0 ? _GEN_1118 : ram_0_13; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2289 = _GEN_734[7:6] == 2'h0 ? _GEN_1119 : ram_0_14; // @[d_cache.scala 175:46 19:24]
  wire [511:0] _GEN_2290 = _GEN_734[7:6] == 2'h0 ? _GEN_1120 : ram_0_15; // @[d_cache.scala 175:46 19:24]
  wire [31:0] _GEN_2291 = _GEN_734[7:6] == 2'h0 ? _GEN_1121 : tag_0_0; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2292 = _GEN_734[7:6] == 2'h0 ? _GEN_1122 : tag_0_1; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2293 = _GEN_734[7:6] == 2'h0 ? _GEN_1123 : tag_0_2; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2294 = _GEN_734[7:6] == 2'h0 ? _GEN_1124 : tag_0_3; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2295 = _GEN_734[7:6] == 2'h0 ? _GEN_1125 : tag_0_4; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2296 = _GEN_734[7:6] == 2'h0 ? _GEN_1126 : tag_0_5; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2297 = _GEN_734[7:6] == 2'h0 ? _GEN_1127 : tag_0_6; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2298 = _GEN_734[7:6] == 2'h0 ? _GEN_1128 : tag_0_7; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2299 = _GEN_734[7:6] == 2'h0 ? _GEN_1129 : tag_0_8; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2300 = _GEN_734[7:6] == 2'h0 ? _GEN_1130 : tag_0_9; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2301 = _GEN_734[7:6] == 2'h0 ? _GEN_1131 : tag_0_10; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2302 = _GEN_734[7:6] == 2'h0 ? _GEN_1132 : tag_0_11; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2303 = _GEN_734[7:6] == 2'h0 ? _GEN_1133 : tag_0_12; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2304 = _GEN_734[7:6] == 2'h0 ? _GEN_1134 : tag_0_13; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2305 = _GEN_734[7:6] == 2'h0 ? _GEN_1135 : tag_0_14; // @[d_cache.scala 175:46 24:24]
  wire [31:0] _GEN_2306 = _GEN_734[7:6] == 2'h0 ? _GEN_1136 : tag_0_15; // @[d_cache.scala 175:46 24:24]
  wire  _GEN_2307 = _GEN_734[7:6] == 2'h0 ? _GEN_1137 : dirty_0_0; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2308 = _GEN_734[7:6] == 2'h0 ? _GEN_1138 : dirty_0_1; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2309 = _GEN_734[7:6] == 2'h0 ? _GEN_1139 : dirty_0_2; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2310 = _GEN_734[7:6] == 2'h0 ? _GEN_1140 : dirty_0_3; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2311 = _GEN_734[7:6] == 2'h0 ? _GEN_1141 : dirty_0_4; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2312 = _GEN_734[7:6] == 2'h0 ? _GEN_1142 : dirty_0_5; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2313 = _GEN_734[7:6] == 2'h0 ? _GEN_1143 : dirty_0_6; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2314 = _GEN_734[7:6] == 2'h0 ? _GEN_1144 : dirty_0_7; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2315 = _GEN_734[7:6] == 2'h0 ? _GEN_1145 : dirty_0_8; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2316 = _GEN_734[7:6] == 2'h0 ? _GEN_1146 : dirty_0_9; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2317 = _GEN_734[7:6] == 2'h0 ? _GEN_1147 : dirty_0_10; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2318 = _GEN_734[7:6] == 2'h0 ? _GEN_1148 : dirty_0_11; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2319 = _GEN_734[7:6] == 2'h0 ? _GEN_1149 : dirty_0_12; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2320 = _GEN_734[7:6] == 2'h0 ? _GEN_1150 : dirty_0_13; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2321 = _GEN_734[7:6] == 2'h0 ? _GEN_1151 : dirty_0_14; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2322 = _GEN_734[7:6] == 2'h0 ? _GEN_1152 : dirty_0_15; // @[d_cache.scala 175:46 34:26]
  wire  _GEN_2323 = _GEN_734[7:6] == 2'h0 ? _GEN_1153 : valid_0_0; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2324 = _GEN_734[7:6] == 2'h0 ? _GEN_1154 : valid_0_1; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2325 = _GEN_734[7:6] == 2'h0 ? _GEN_1155 : valid_0_2; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2326 = _GEN_734[7:6] == 2'h0 ? _GEN_1156 : valid_0_3; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2327 = _GEN_734[7:6] == 2'h0 ? _GEN_1157 : valid_0_4; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2328 = _GEN_734[7:6] == 2'h0 ? _GEN_1158 : valid_0_5; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2329 = _GEN_734[7:6] == 2'h0 ? _GEN_1159 : valid_0_6; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2330 = _GEN_734[7:6] == 2'h0 ? _GEN_1160 : valid_0_7; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2331 = _GEN_734[7:6] == 2'h0 ? _GEN_1161 : valid_0_8; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2332 = _GEN_734[7:6] == 2'h0 ? _GEN_1162 : valid_0_9; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2333 = _GEN_734[7:6] == 2'h0 ? _GEN_1163 : valid_0_10; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2334 = _GEN_734[7:6] == 2'h0 ? _GEN_1164 : valid_0_11; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2335 = _GEN_734[7:6] == 2'h0 ? _GEN_1165 : valid_0_12; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2336 = _GEN_734[7:6] == 2'h0 ? _GEN_1166 : valid_0_13; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2337 = _GEN_734[7:6] == 2'h0 ? _GEN_1167 : valid_0_14; // @[d_cache.scala 175:46 29:26]
  wire  _GEN_2338 = _GEN_734[7:6] == 2'h0 ? _GEN_1168 : valid_0_15; // @[d_cache.scala 175:46 29:26]
  wire [3:0] _GEN_2339 = _GEN_734[7:6] == 2'h0 ? _GEN_1169 : _GEN_2128; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2340 = _GEN_734[7:6] == 2'h0 ? _GEN_1170 : _GEN_2129; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2341 = _GEN_734[7:6] == 2'h0 ? _GEN_1171 : _GEN_2130; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2342 = _GEN_734[7:6] == 2'h0 ? _GEN_1172 : _GEN_2131; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2343 = _GEN_734[7:6] == 2'h0 ? _GEN_1173 : _GEN_2132; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2344 = _GEN_734[7:6] == 2'h0 ? _GEN_1174 : _GEN_2133; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2345 = _GEN_734[7:6] == 2'h0 ? _GEN_1175 : _GEN_2134; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2346 = _GEN_734[7:6] == 2'h0 ? _GEN_1176 : _GEN_2135; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2347 = _GEN_734[7:6] == 2'h0 ? _GEN_1177 : _GEN_2136; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2348 = _GEN_734[7:6] == 2'h0 ? _GEN_1178 : _GEN_2137; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2349 = _GEN_734[7:6] == 2'h0 ? _GEN_1179 : _GEN_2138; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2350 = _GEN_734[7:6] == 2'h0 ? _GEN_1180 : _GEN_2139; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2351 = _GEN_734[7:6] == 2'h0 ? _GEN_1181 : _GEN_2140; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2352 = _GEN_734[7:6] == 2'h0 ? _GEN_1182 : _GEN_2141; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2353 = _GEN_734[7:6] == 2'h0 ? _GEN_1183 : _GEN_2142; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2354 = _GEN_734[7:6] == 2'h0 ? _GEN_1184 : _GEN_2143; // @[d_cache.scala 175:46]
  wire [7:0] _GEN_2355 = _GEN_734[7:6] == 2'h0 ? _GEN_1185 : _GEN_2144; // @[d_cache.scala 175:46]
  wire [511:0] _GEN_2356 = _GEN_734[7:6] == 2'h0 ? ram_1_0 : _GEN_2064; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2357 = _GEN_734[7:6] == 2'h0 ? ram_1_1 : _GEN_2065; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2358 = _GEN_734[7:6] == 2'h0 ? ram_1_2 : _GEN_2066; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2359 = _GEN_734[7:6] == 2'h0 ? ram_1_3 : _GEN_2067; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2360 = _GEN_734[7:6] == 2'h0 ? ram_1_4 : _GEN_2068; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2361 = _GEN_734[7:6] == 2'h0 ? ram_1_5 : _GEN_2069; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2362 = _GEN_734[7:6] == 2'h0 ? ram_1_6 : _GEN_2070; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2363 = _GEN_734[7:6] == 2'h0 ? ram_1_7 : _GEN_2071; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2364 = _GEN_734[7:6] == 2'h0 ? ram_1_8 : _GEN_2072; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2365 = _GEN_734[7:6] == 2'h0 ? ram_1_9 : _GEN_2073; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2366 = _GEN_734[7:6] == 2'h0 ? ram_1_10 : _GEN_2074; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2367 = _GEN_734[7:6] == 2'h0 ? ram_1_11 : _GEN_2075; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2368 = _GEN_734[7:6] == 2'h0 ? ram_1_12 : _GEN_2076; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2369 = _GEN_734[7:6] == 2'h0 ? ram_1_13 : _GEN_2077; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2370 = _GEN_734[7:6] == 2'h0 ? ram_1_14 : _GEN_2078; // @[d_cache.scala 175:46 20:24]
  wire [511:0] _GEN_2371 = _GEN_734[7:6] == 2'h0 ? ram_1_15 : _GEN_2079; // @[d_cache.scala 175:46 20:24]
  wire [31:0] _GEN_2372 = _GEN_734[7:6] == 2'h0 ? tag_1_0 : _GEN_2080; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2373 = _GEN_734[7:6] == 2'h0 ? tag_1_1 : _GEN_2081; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2374 = _GEN_734[7:6] == 2'h0 ? tag_1_2 : _GEN_2082; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2375 = _GEN_734[7:6] == 2'h0 ? tag_1_3 : _GEN_2083; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2376 = _GEN_734[7:6] == 2'h0 ? tag_1_4 : _GEN_2084; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2377 = _GEN_734[7:6] == 2'h0 ? tag_1_5 : _GEN_2085; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2378 = _GEN_734[7:6] == 2'h0 ? tag_1_6 : _GEN_2086; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2379 = _GEN_734[7:6] == 2'h0 ? tag_1_7 : _GEN_2087; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2380 = _GEN_734[7:6] == 2'h0 ? tag_1_8 : _GEN_2088; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2381 = _GEN_734[7:6] == 2'h0 ? tag_1_9 : _GEN_2089; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2382 = _GEN_734[7:6] == 2'h0 ? tag_1_10 : _GEN_2090; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2383 = _GEN_734[7:6] == 2'h0 ? tag_1_11 : _GEN_2091; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2384 = _GEN_734[7:6] == 2'h0 ? tag_1_12 : _GEN_2092; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2385 = _GEN_734[7:6] == 2'h0 ? tag_1_13 : _GEN_2093; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2386 = _GEN_734[7:6] == 2'h0 ? tag_1_14 : _GEN_2094; // @[d_cache.scala 175:46 25:24]
  wire [31:0] _GEN_2387 = _GEN_734[7:6] == 2'h0 ? tag_1_15 : _GEN_2095; // @[d_cache.scala 175:46 25:24]
  wire  _GEN_2388 = _GEN_734[7:6] == 2'h0 ? dirty_1_0 : _GEN_2096; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2389 = _GEN_734[7:6] == 2'h0 ? dirty_1_1 : _GEN_2097; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2390 = _GEN_734[7:6] == 2'h0 ? dirty_1_2 : _GEN_2098; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2391 = _GEN_734[7:6] == 2'h0 ? dirty_1_3 : _GEN_2099; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2392 = _GEN_734[7:6] == 2'h0 ? dirty_1_4 : _GEN_2100; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2393 = _GEN_734[7:6] == 2'h0 ? dirty_1_5 : _GEN_2101; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2394 = _GEN_734[7:6] == 2'h0 ? dirty_1_6 : _GEN_2102; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2395 = _GEN_734[7:6] == 2'h0 ? dirty_1_7 : _GEN_2103; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2396 = _GEN_734[7:6] == 2'h0 ? dirty_1_8 : _GEN_2104; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2397 = _GEN_734[7:6] == 2'h0 ? dirty_1_9 : _GEN_2105; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2398 = _GEN_734[7:6] == 2'h0 ? dirty_1_10 : _GEN_2106; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2399 = _GEN_734[7:6] == 2'h0 ? dirty_1_11 : _GEN_2107; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2400 = _GEN_734[7:6] == 2'h0 ? dirty_1_12 : _GEN_2108; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2401 = _GEN_734[7:6] == 2'h0 ? dirty_1_13 : _GEN_2109; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2402 = _GEN_734[7:6] == 2'h0 ? dirty_1_14 : _GEN_2110; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2403 = _GEN_734[7:6] == 2'h0 ? dirty_1_15 : _GEN_2111; // @[d_cache.scala 175:46 35:26]
  wire  _GEN_2404 = _GEN_734[7:6] == 2'h0 ? valid_1_0 : _GEN_2112; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2405 = _GEN_734[7:6] == 2'h0 ? valid_1_1 : _GEN_2113; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2406 = _GEN_734[7:6] == 2'h0 ? valid_1_2 : _GEN_2114; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2407 = _GEN_734[7:6] == 2'h0 ? valid_1_3 : _GEN_2115; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2408 = _GEN_734[7:6] == 2'h0 ? valid_1_4 : _GEN_2116; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2409 = _GEN_734[7:6] == 2'h0 ? valid_1_5 : _GEN_2117; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2410 = _GEN_734[7:6] == 2'h0 ? valid_1_6 : _GEN_2118; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2411 = _GEN_734[7:6] == 2'h0 ? valid_1_7 : _GEN_2119; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2412 = _GEN_734[7:6] == 2'h0 ? valid_1_8 : _GEN_2120; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2413 = _GEN_734[7:6] == 2'h0 ? valid_1_9 : _GEN_2121; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2414 = _GEN_734[7:6] == 2'h0 ? valid_1_10 : _GEN_2122; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2415 = _GEN_734[7:6] == 2'h0 ? valid_1_11 : _GEN_2123; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2416 = _GEN_734[7:6] == 2'h0 ? valid_1_12 : _GEN_2124; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2417 = _GEN_734[7:6] == 2'h0 ? valid_1_13 : _GEN_2125; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2418 = _GEN_734[7:6] == 2'h0 ? valid_1_14 : _GEN_2126; // @[d_cache.scala 175:46 30:26]
  wire  _GEN_2419 = _GEN_734[7:6] == 2'h0 ? valid_1_15 : _GEN_2127; // @[d_cache.scala 175:46 30:26]
  wire [511:0] _GEN_2420 = _GEN_734[7:6] == 2'h0 ? ram_2_0 : _GEN_2145; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2421 = _GEN_734[7:6] == 2'h0 ? ram_2_1 : _GEN_2146; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2422 = _GEN_734[7:6] == 2'h0 ? ram_2_2 : _GEN_2147; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2423 = _GEN_734[7:6] == 2'h0 ? ram_2_3 : _GEN_2148; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2424 = _GEN_734[7:6] == 2'h0 ? ram_2_4 : _GEN_2149; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2425 = _GEN_734[7:6] == 2'h0 ? ram_2_5 : _GEN_2150; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2426 = _GEN_734[7:6] == 2'h0 ? ram_2_6 : _GEN_2151; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2427 = _GEN_734[7:6] == 2'h0 ? ram_2_7 : _GEN_2152; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2428 = _GEN_734[7:6] == 2'h0 ? ram_2_8 : _GEN_2153; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2429 = _GEN_734[7:6] == 2'h0 ? ram_2_9 : _GEN_2154; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2430 = _GEN_734[7:6] == 2'h0 ? ram_2_10 : _GEN_2155; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2431 = _GEN_734[7:6] == 2'h0 ? ram_2_11 : _GEN_2156; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2432 = _GEN_734[7:6] == 2'h0 ? ram_2_12 : _GEN_2157; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2433 = _GEN_734[7:6] == 2'h0 ? ram_2_13 : _GEN_2158; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2434 = _GEN_734[7:6] == 2'h0 ? ram_2_14 : _GEN_2159; // @[d_cache.scala 175:46 21:24]
  wire [511:0] _GEN_2435 = _GEN_734[7:6] == 2'h0 ? ram_2_15 : _GEN_2160; // @[d_cache.scala 175:46 21:24]
  wire [31:0] _GEN_2436 = _GEN_734[7:6] == 2'h0 ? tag_2_0 : _GEN_2161; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2437 = _GEN_734[7:6] == 2'h0 ? tag_2_1 : _GEN_2162; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2438 = _GEN_734[7:6] == 2'h0 ? tag_2_2 : _GEN_2163; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2439 = _GEN_734[7:6] == 2'h0 ? tag_2_3 : _GEN_2164; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2440 = _GEN_734[7:6] == 2'h0 ? tag_2_4 : _GEN_2165; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2441 = _GEN_734[7:6] == 2'h0 ? tag_2_5 : _GEN_2166; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2442 = _GEN_734[7:6] == 2'h0 ? tag_2_6 : _GEN_2167; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2443 = _GEN_734[7:6] == 2'h0 ? tag_2_7 : _GEN_2168; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2444 = _GEN_734[7:6] == 2'h0 ? tag_2_8 : _GEN_2169; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2445 = _GEN_734[7:6] == 2'h0 ? tag_2_9 : _GEN_2170; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2446 = _GEN_734[7:6] == 2'h0 ? tag_2_10 : _GEN_2171; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2447 = _GEN_734[7:6] == 2'h0 ? tag_2_11 : _GEN_2172; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2448 = _GEN_734[7:6] == 2'h0 ? tag_2_12 : _GEN_2173; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2449 = _GEN_734[7:6] == 2'h0 ? tag_2_13 : _GEN_2174; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2450 = _GEN_734[7:6] == 2'h0 ? tag_2_14 : _GEN_2175; // @[d_cache.scala 175:46 26:24]
  wire [31:0] _GEN_2451 = _GEN_734[7:6] == 2'h0 ? tag_2_15 : _GEN_2176; // @[d_cache.scala 175:46 26:24]
  wire  _GEN_2452 = _GEN_734[7:6] == 2'h0 ? dirty_2_0 : _GEN_2177; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2453 = _GEN_734[7:6] == 2'h0 ? dirty_2_1 : _GEN_2178; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2454 = _GEN_734[7:6] == 2'h0 ? dirty_2_2 : _GEN_2179; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2455 = _GEN_734[7:6] == 2'h0 ? dirty_2_3 : _GEN_2180; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2456 = _GEN_734[7:6] == 2'h0 ? dirty_2_4 : _GEN_2181; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2457 = _GEN_734[7:6] == 2'h0 ? dirty_2_5 : _GEN_2182; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2458 = _GEN_734[7:6] == 2'h0 ? dirty_2_6 : _GEN_2183; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2459 = _GEN_734[7:6] == 2'h0 ? dirty_2_7 : _GEN_2184; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2460 = _GEN_734[7:6] == 2'h0 ? dirty_2_8 : _GEN_2185; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2461 = _GEN_734[7:6] == 2'h0 ? dirty_2_9 : _GEN_2186; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2462 = _GEN_734[7:6] == 2'h0 ? dirty_2_10 : _GEN_2187; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2463 = _GEN_734[7:6] == 2'h0 ? dirty_2_11 : _GEN_2188; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2464 = _GEN_734[7:6] == 2'h0 ? dirty_2_12 : _GEN_2189; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2465 = _GEN_734[7:6] == 2'h0 ? dirty_2_13 : _GEN_2190; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2466 = _GEN_734[7:6] == 2'h0 ? dirty_2_14 : _GEN_2191; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2467 = _GEN_734[7:6] == 2'h0 ? dirty_2_15 : _GEN_2192; // @[d_cache.scala 175:46 36:26]
  wire  _GEN_2468 = _GEN_734[7:6] == 2'h0 ? valid_2_0 : _GEN_2193; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2469 = _GEN_734[7:6] == 2'h0 ? valid_2_1 : _GEN_2194; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2470 = _GEN_734[7:6] == 2'h0 ? valid_2_2 : _GEN_2195; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2471 = _GEN_734[7:6] == 2'h0 ? valid_2_3 : _GEN_2196; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2472 = _GEN_734[7:6] == 2'h0 ? valid_2_4 : _GEN_2197; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2473 = _GEN_734[7:6] == 2'h0 ? valid_2_5 : _GEN_2198; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2474 = _GEN_734[7:6] == 2'h0 ? valid_2_6 : _GEN_2199; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2475 = _GEN_734[7:6] == 2'h0 ? valid_2_7 : _GEN_2200; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2476 = _GEN_734[7:6] == 2'h0 ? valid_2_8 : _GEN_2201; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2477 = _GEN_734[7:6] == 2'h0 ? valid_2_9 : _GEN_2202; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2478 = _GEN_734[7:6] == 2'h0 ? valid_2_10 : _GEN_2203; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2479 = _GEN_734[7:6] == 2'h0 ? valid_2_11 : _GEN_2204; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2480 = _GEN_734[7:6] == 2'h0 ? valid_2_12 : _GEN_2205; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2481 = _GEN_734[7:6] == 2'h0 ? valid_2_13 : _GEN_2206; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2482 = _GEN_734[7:6] == 2'h0 ? valid_2_14 : _GEN_2207; // @[d_cache.scala 175:46 31:26]
  wire  _GEN_2483 = _GEN_734[7:6] == 2'h0 ? valid_2_15 : _GEN_2208; // @[d_cache.scala 175:46 31:26]
  wire [511:0] _GEN_2484 = _GEN_734[7:6] == 2'h0 ? ram_3_0 : _GEN_2209; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2485 = _GEN_734[7:6] == 2'h0 ? ram_3_1 : _GEN_2210; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2486 = _GEN_734[7:6] == 2'h0 ? ram_3_2 : _GEN_2211; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2487 = _GEN_734[7:6] == 2'h0 ? ram_3_3 : _GEN_2212; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2488 = _GEN_734[7:6] == 2'h0 ? ram_3_4 : _GEN_2213; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2489 = _GEN_734[7:6] == 2'h0 ? ram_3_5 : _GEN_2214; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2490 = _GEN_734[7:6] == 2'h0 ? ram_3_6 : _GEN_2215; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2491 = _GEN_734[7:6] == 2'h0 ? ram_3_7 : _GEN_2216; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2492 = _GEN_734[7:6] == 2'h0 ? ram_3_8 : _GEN_2217; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2493 = _GEN_734[7:6] == 2'h0 ? ram_3_9 : _GEN_2218; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2494 = _GEN_734[7:6] == 2'h0 ? ram_3_10 : _GEN_2219; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2495 = _GEN_734[7:6] == 2'h0 ? ram_3_11 : _GEN_2220; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2496 = _GEN_734[7:6] == 2'h0 ? ram_3_12 : _GEN_2221; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2497 = _GEN_734[7:6] == 2'h0 ? ram_3_13 : _GEN_2222; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2498 = _GEN_734[7:6] == 2'h0 ? ram_3_14 : _GEN_2223; // @[d_cache.scala 175:46 22:24]
  wire [511:0] _GEN_2499 = _GEN_734[7:6] == 2'h0 ? ram_3_15 : _GEN_2224; // @[d_cache.scala 175:46 22:24]
  wire [31:0] _GEN_2500 = _GEN_734[7:6] == 2'h0 ? tag_3_0 : _GEN_2225; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2501 = _GEN_734[7:6] == 2'h0 ? tag_3_1 : _GEN_2226; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2502 = _GEN_734[7:6] == 2'h0 ? tag_3_2 : _GEN_2227; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2503 = _GEN_734[7:6] == 2'h0 ? tag_3_3 : _GEN_2228; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2504 = _GEN_734[7:6] == 2'h0 ? tag_3_4 : _GEN_2229; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2505 = _GEN_734[7:6] == 2'h0 ? tag_3_5 : _GEN_2230; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2506 = _GEN_734[7:6] == 2'h0 ? tag_3_6 : _GEN_2231; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2507 = _GEN_734[7:6] == 2'h0 ? tag_3_7 : _GEN_2232; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2508 = _GEN_734[7:6] == 2'h0 ? tag_3_8 : _GEN_2233; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2509 = _GEN_734[7:6] == 2'h0 ? tag_3_9 : _GEN_2234; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2510 = _GEN_734[7:6] == 2'h0 ? tag_3_10 : _GEN_2235; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2511 = _GEN_734[7:6] == 2'h0 ? tag_3_11 : _GEN_2236; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2512 = _GEN_734[7:6] == 2'h0 ? tag_3_12 : _GEN_2237; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2513 = _GEN_734[7:6] == 2'h0 ? tag_3_13 : _GEN_2238; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2514 = _GEN_734[7:6] == 2'h0 ? tag_3_14 : _GEN_2239; // @[d_cache.scala 175:46 27:24]
  wire [31:0] _GEN_2515 = _GEN_734[7:6] == 2'h0 ? tag_3_15 : _GEN_2240; // @[d_cache.scala 175:46 27:24]
  wire  _GEN_2516 = _GEN_734[7:6] == 2'h0 ? dirty_3_0 : _GEN_2241; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2517 = _GEN_734[7:6] == 2'h0 ? dirty_3_1 : _GEN_2242; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2518 = _GEN_734[7:6] == 2'h0 ? dirty_3_2 : _GEN_2243; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2519 = _GEN_734[7:6] == 2'h0 ? dirty_3_3 : _GEN_2244; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2520 = _GEN_734[7:6] == 2'h0 ? dirty_3_4 : _GEN_2245; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2521 = _GEN_734[7:6] == 2'h0 ? dirty_3_5 : _GEN_2246; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2522 = _GEN_734[7:6] == 2'h0 ? dirty_3_6 : _GEN_2247; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2523 = _GEN_734[7:6] == 2'h0 ? dirty_3_7 : _GEN_2248; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2524 = _GEN_734[7:6] == 2'h0 ? dirty_3_8 : _GEN_2249; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2525 = _GEN_734[7:6] == 2'h0 ? dirty_3_9 : _GEN_2250; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2526 = _GEN_734[7:6] == 2'h0 ? dirty_3_10 : _GEN_2251; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2527 = _GEN_734[7:6] == 2'h0 ? dirty_3_11 : _GEN_2252; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2528 = _GEN_734[7:6] == 2'h0 ? dirty_3_12 : _GEN_2253; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2529 = _GEN_734[7:6] == 2'h0 ? dirty_3_13 : _GEN_2254; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2530 = _GEN_734[7:6] == 2'h0 ? dirty_3_14 : _GEN_2255; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2531 = _GEN_734[7:6] == 2'h0 ? dirty_3_15 : _GEN_2256; // @[d_cache.scala 175:46 37:26]
  wire  _GEN_2532 = _GEN_734[7:6] == 2'h0 ? valid_3_0 : _GEN_2257; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2533 = _GEN_734[7:6] == 2'h0 ? valid_3_1 : _GEN_2258; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2534 = _GEN_734[7:6] == 2'h0 ? valid_3_2 : _GEN_2259; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2535 = _GEN_734[7:6] == 2'h0 ? valid_3_3 : _GEN_2260; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2536 = _GEN_734[7:6] == 2'h0 ? valid_3_4 : _GEN_2261; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2537 = _GEN_734[7:6] == 2'h0 ? valid_3_5 : _GEN_2262; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2538 = _GEN_734[7:6] == 2'h0 ? valid_3_6 : _GEN_2263; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2539 = _GEN_734[7:6] == 2'h0 ? valid_3_7 : _GEN_2264; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2540 = _GEN_734[7:6] == 2'h0 ? valid_3_8 : _GEN_2265; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2541 = _GEN_734[7:6] == 2'h0 ? valid_3_9 : _GEN_2266; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2542 = _GEN_734[7:6] == 2'h0 ? valid_3_10 : _GEN_2267; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2543 = _GEN_734[7:6] == 2'h0 ? valid_3_11 : _GEN_2268; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2544 = _GEN_734[7:6] == 2'h0 ? valid_3_12 : _GEN_2269; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2545 = _GEN_734[7:6] == 2'h0 ? valid_3_13 : _GEN_2270; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2546 = _GEN_734[7:6] == 2'h0 ? valid_3_14 : _GEN_2271; // @[d_cache.scala 175:46 32:26]
  wire  _GEN_2547 = _GEN_734[7:6] == 2'h0 ? valid_3_15 : _GEN_2272; // @[d_cache.scala 175:46 32:26]
  wire [3:0] _GEN_2548 = unuse_way == 3'h4 ? 4'h1 : _GEN_2339; // @[d_cache.scala 168:40 169:23]
  wire [511:0] _GEN_2549 = unuse_way == 3'h4 ? _GEN_879 : _GEN_2484; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2550 = unuse_way == 3'h4 ? _GEN_880 : _GEN_2485; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2551 = unuse_way == 3'h4 ? _GEN_881 : _GEN_2486; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2552 = unuse_way == 3'h4 ? _GEN_882 : _GEN_2487; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2553 = unuse_way == 3'h4 ? _GEN_883 : _GEN_2488; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2554 = unuse_way == 3'h4 ? _GEN_884 : _GEN_2489; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2555 = unuse_way == 3'h4 ? _GEN_885 : _GEN_2490; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2556 = unuse_way == 3'h4 ? _GEN_886 : _GEN_2491; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2557 = unuse_way == 3'h4 ? _GEN_887 : _GEN_2492; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2558 = unuse_way == 3'h4 ? _GEN_888 : _GEN_2493; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2559 = unuse_way == 3'h4 ? _GEN_889 : _GEN_2494; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2560 = unuse_way == 3'h4 ? _GEN_890 : _GEN_2495; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2561 = unuse_way == 3'h4 ? _GEN_891 : _GEN_2496; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2562 = unuse_way == 3'h4 ? _GEN_892 : _GEN_2497; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2563 = unuse_way == 3'h4 ? _GEN_893 : _GEN_2498; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2564 = unuse_way == 3'h4 ? _GEN_894 : _GEN_2499; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2565 = unuse_way == 3'h4 ? _GEN_895 : _GEN_2500; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2566 = unuse_way == 3'h4 ? _GEN_896 : _GEN_2501; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2567 = unuse_way == 3'h4 ? _GEN_897 : _GEN_2502; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2568 = unuse_way == 3'h4 ? _GEN_898 : _GEN_2503; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2569 = unuse_way == 3'h4 ? _GEN_899 : _GEN_2504; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2570 = unuse_way == 3'h4 ? _GEN_900 : _GEN_2505; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2571 = unuse_way == 3'h4 ? _GEN_901 : _GEN_2506; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2572 = unuse_way == 3'h4 ? _GEN_902 : _GEN_2507; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2573 = unuse_way == 3'h4 ? _GEN_903 : _GEN_2508; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2574 = unuse_way == 3'h4 ? _GEN_904 : _GEN_2509; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2575 = unuse_way == 3'h4 ? _GEN_905 : _GEN_2510; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2576 = unuse_way == 3'h4 ? _GEN_906 : _GEN_2511; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2577 = unuse_way == 3'h4 ? _GEN_907 : _GEN_2512; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2578 = unuse_way == 3'h4 ? _GEN_908 : _GEN_2513; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2579 = unuse_way == 3'h4 ? _GEN_909 : _GEN_2514; // @[d_cache.scala 168:40]
  wire [31:0] _GEN_2580 = unuse_way == 3'h4 ? _GEN_910 : _GEN_2515; // @[d_cache.scala 168:40]
  wire  _GEN_2581 = unuse_way == 3'h4 ? _GEN_911 : _GEN_2532; // @[d_cache.scala 168:40]
  wire  _GEN_2582 = unuse_way == 3'h4 ? _GEN_912 : _GEN_2533; // @[d_cache.scala 168:40]
  wire  _GEN_2583 = unuse_way == 3'h4 ? _GEN_913 : _GEN_2534; // @[d_cache.scala 168:40]
  wire  _GEN_2584 = unuse_way == 3'h4 ? _GEN_914 : _GEN_2535; // @[d_cache.scala 168:40]
  wire  _GEN_2585 = unuse_way == 3'h4 ? _GEN_915 : _GEN_2536; // @[d_cache.scala 168:40]
  wire  _GEN_2586 = unuse_way == 3'h4 ? _GEN_916 : _GEN_2537; // @[d_cache.scala 168:40]
  wire  _GEN_2587 = unuse_way == 3'h4 ? _GEN_917 : _GEN_2538; // @[d_cache.scala 168:40]
  wire  _GEN_2588 = unuse_way == 3'h4 ? _GEN_918 : _GEN_2539; // @[d_cache.scala 168:40]
  wire  _GEN_2589 = unuse_way == 3'h4 ? _GEN_919 : _GEN_2540; // @[d_cache.scala 168:40]
  wire  _GEN_2590 = unuse_way == 3'h4 ? _GEN_920 : _GEN_2541; // @[d_cache.scala 168:40]
  wire  _GEN_2591 = unuse_way == 3'h4 ? _GEN_921 : _GEN_2542; // @[d_cache.scala 168:40]
  wire  _GEN_2592 = unuse_way == 3'h4 ? _GEN_922 : _GEN_2543; // @[d_cache.scala 168:40]
  wire  _GEN_2593 = unuse_way == 3'h4 ? _GEN_923 : _GEN_2544; // @[d_cache.scala 168:40]
  wire  _GEN_2594 = unuse_way == 3'h4 ? _GEN_924 : _GEN_2545; // @[d_cache.scala 168:40]
  wire  _GEN_2595 = unuse_way == 3'h4 ? _GEN_925 : _GEN_2546; // @[d_cache.scala 168:40]
  wire  _GEN_2596 = unuse_way == 3'h4 ? _GEN_926 : _GEN_2547; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2597 = unuse_way == 3'h4 ? _GEN_927 : _GEN_2340; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2598 = unuse_way == 3'h4 ? _GEN_928 : _GEN_2341; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2599 = unuse_way == 3'h4 ? _GEN_929 : _GEN_2342; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2600 = unuse_way == 3'h4 ? _GEN_930 : _GEN_2343; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2601 = unuse_way == 3'h4 ? _GEN_931 : _GEN_2344; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2602 = unuse_way == 3'h4 ? _GEN_932 : _GEN_2345; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2603 = unuse_way == 3'h4 ? _GEN_933 : _GEN_2346; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2604 = unuse_way == 3'h4 ? _GEN_934 : _GEN_2347; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2605 = unuse_way == 3'h4 ? _GEN_935 : _GEN_2348; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2606 = unuse_way == 3'h4 ? _GEN_936 : _GEN_2349; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2607 = unuse_way == 3'h4 ? _GEN_937 : _GEN_2350; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2608 = unuse_way == 3'h4 ? _GEN_938 : _GEN_2351; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2609 = unuse_way == 3'h4 ? _GEN_939 : _GEN_2352; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2610 = unuse_way == 3'h4 ? _GEN_940 : _GEN_2353; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2611 = unuse_way == 3'h4 ? _GEN_941 : _GEN_2354; // @[d_cache.scala 168:40]
  wire [7:0] _GEN_2612 = unuse_way == 3'h4 ? _GEN_942 : _GEN_2355; // @[d_cache.scala 168:40]
  wire [511:0] _GEN_2613 = unuse_way == 3'h4 ? write_back_data : _GEN_2273; // @[d_cache.scala 168:40 44:34]
  wire [41:0] _GEN_2614 = unuse_way == 3'h4 ? {{10'd0}, write_back_addr} : _GEN_2274; // @[d_cache.scala 168:40 45:34]
  wire [511:0] _GEN_2615 = unuse_way == 3'h4 ? ram_0_0 : _GEN_2275; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2616 = unuse_way == 3'h4 ? ram_0_1 : _GEN_2276; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2617 = unuse_way == 3'h4 ? ram_0_2 : _GEN_2277; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2618 = unuse_way == 3'h4 ? ram_0_3 : _GEN_2278; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2619 = unuse_way == 3'h4 ? ram_0_4 : _GEN_2279; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2620 = unuse_way == 3'h4 ? ram_0_5 : _GEN_2280; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2621 = unuse_way == 3'h4 ? ram_0_6 : _GEN_2281; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2622 = unuse_way == 3'h4 ? ram_0_7 : _GEN_2282; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2623 = unuse_way == 3'h4 ? ram_0_8 : _GEN_2283; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2624 = unuse_way == 3'h4 ? ram_0_9 : _GEN_2284; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2625 = unuse_way == 3'h4 ? ram_0_10 : _GEN_2285; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2626 = unuse_way == 3'h4 ? ram_0_11 : _GEN_2286; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2627 = unuse_way == 3'h4 ? ram_0_12 : _GEN_2287; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2628 = unuse_way == 3'h4 ? ram_0_13 : _GEN_2288; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2629 = unuse_way == 3'h4 ? ram_0_14 : _GEN_2289; // @[d_cache.scala 168:40 19:24]
  wire [511:0] _GEN_2630 = unuse_way == 3'h4 ? ram_0_15 : _GEN_2290; // @[d_cache.scala 168:40 19:24]
  wire [31:0] _GEN_2631 = unuse_way == 3'h4 ? tag_0_0 : _GEN_2291; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2632 = unuse_way == 3'h4 ? tag_0_1 : _GEN_2292; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2633 = unuse_way == 3'h4 ? tag_0_2 : _GEN_2293; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2634 = unuse_way == 3'h4 ? tag_0_3 : _GEN_2294; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2635 = unuse_way == 3'h4 ? tag_0_4 : _GEN_2295; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2636 = unuse_way == 3'h4 ? tag_0_5 : _GEN_2296; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2637 = unuse_way == 3'h4 ? tag_0_6 : _GEN_2297; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2638 = unuse_way == 3'h4 ? tag_0_7 : _GEN_2298; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2639 = unuse_way == 3'h4 ? tag_0_8 : _GEN_2299; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2640 = unuse_way == 3'h4 ? tag_0_9 : _GEN_2300; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2641 = unuse_way == 3'h4 ? tag_0_10 : _GEN_2301; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2642 = unuse_way == 3'h4 ? tag_0_11 : _GEN_2302; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2643 = unuse_way == 3'h4 ? tag_0_12 : _GEN_2303; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2644 = unuse_way == 3'h4 ? tag_0_13 : _GEN_2304; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2645 = unuse_way == 3'h4 ? tag_0_14 : _GEN_2305; // @[d_cache.scala 168:40 24:24]
  wire [31:0] _GEN_2646 = unuse_way == 3'h4 ? tag_0_15 : _GEN_2306; // @[d_cache.scala 168:40 24:24]
  wire  _GEN_2647 = unuse_way == 3'h4 ? dirty_0_0 : _GEN_2307; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2648 = unuse_way == 3'h4 ? dirty_0_1 : _GEN_2308; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2649 = unuse_way == 3'h4 ? dirty_0_2 : _GEN_2309; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2650 = unuse_way == 3'h4 ? dirty_0_3 : _GEN_2310; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2651 = unuse_way == 3'h4 ? dirty_0_4 : _GEN_2311; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2652 = unuse_way == 3'h4 ? dirty_0_5 : _GEN_2312; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2653 = unuse_way == 3'h4 ? dirty_0_6 : _GEN_2313; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2654 = unuse_way == 3'h4 ? dirty_0_7 : _GEN_2314; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2655 = unuse_way == 3'h4 ? dirty_0_8 : _GEN_2315; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2656 = unuse_way == 3'h4 ? dirty_0_9 : _GEN_2316; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2657 = unuse_way == 3'h4 ? dirty_0_10 : _GEN_2317; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2658 = unuse_way == 3'h4 ? dirty_0_11 : _GEN_2318; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2659 = unuse_way == 3'h4 ? dirty_0_12 : _GEN_2319; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2660 = unuse_way == 3'h4 ? dirty_0_13 : _GEN_2320; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2661 = unuse_way == 3'h4 ? dirty_0_14 : _GEN_2321; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2662 = unuse_way == 3'h4 ? dirty_0_15 : _GEN_2322; // @[d_cache.scala 168:40 34:26]
  wire  _GEN_2663 = unuse_way == 3'h4 ? valid_0_0 : _GEN_2323; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2664 = unuse_way == 3'h4 ? valid_0_1 : _GEN_2324; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2665 = unuse_way == 3'h4 ? valid_0_2 : _GEN_2325; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2666 = unuse_way == 3'h4 ? valid_0_3 : _GEN_2326; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2667 = unuse_way == 3'h4 ? valid_0_4 : _GEN_2327; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2668 = unuse_way == 3'h4 ? valid_0_5 : _GEN_2328; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2669 = unuse_way == 3'h4 ? valid_0_6 : _GEN_2329; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2670 = unuse_way == 3'h4 ? valid_0_7 : _GEN_2330; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2671 = unuse_way == 3'h4 ? valid_0_8 : _GEN_2331; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2672 = unuse_way == 3'h4 ? valid_0_9 : _GEN_2332; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2673 = unuse_way == 3'h4 ? valid_0_10 : _GEN_2333; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2674 = unuse_way == 3'h4 ? valid_0_11 : _GEN_2334; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2675 = unuse_way == 3'h4 ? valid_0_12 : _GEN_2335; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2676 = unuse_way == 3'h4 ? valid_0_13 : _GEN_2336; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2677 = unuse_way == 3'h4 ? valid_0_14 : _GEN_2337; // @[d_cache.scala 168:40 29:26]
  wire  _GEN_2678 = unuse_way == 3'h4 ? valid_0_15 : _GEN_2338; // @[d_cache.scala 168:40 29:26]
  wire [511:0] _GEN_2679 = unuse_way == 3'h4 ? ram_1_0 : _GEN_2356; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2680 = unuse_way == 3'h4 ? ram_1_1 : _GEN_2357; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2681 = unuse_way == 3'h4 ? ram_1_2 : _GEN_2358; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2682 = unuse_way == 3'h4 ? ram_1_3 : _GEN_2359; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2683 = unuse_way == 3'h4 ? ram_1_4 : _GEN_2360; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2684 = unuse_way == 3'h4 ? ram_1_5 : _GEN_2361; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2685 = unuse_way == 3'h4 ? ram_1_6 : _GEN_2362; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2686 = unuse_way == 3'h4 ? ram_1_7 : _GEN_2363; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2687 = unuse_way == 3'h4 ? ram_1_8 : _GEN_2364; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2688 = unuse_way == 3'h4 ? ram_1_9 : _GEN_2365; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2689 = unuse_way == 3'h4 ? ram_1_10 : _GEN_2366; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2690 = unuse_way == 3'h4 ? ram_1_11 : _GEN_2367; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2691 = unuse_way == 3'h4 ? ram_1_12 : _GEN_2368; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2692 = unuse_way == 3'h4 ? ram_1_13 : _GEN_2369; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2693 = unuse_way == 3'h4 ? ram_1_14 : _GEN_2370; // @[d_cache.scala 168:40 20:24]
  wire [511:0] _GEN_2694 = unuse_way == 3'h4 ? ram_1_15 : _GEN_2371; // @[d_cache.scala 168:40 20:24]
  wire [31:0] _GEN_2695 = unuse_way == 3'h4 ? tag_1_0 : _GEN_2372; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2696 = unuse_way == 3'h4 ? tag_1_1 : _GEN_2373; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2697 = unuse_way == 3'h4 ? tag_1_2 : _GEN_2374; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2698 = unuse_way == 3'h4 ? tag_1_3 : _GEN_2375; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2699 = unuse_way == 3'h4 ? tag_1_4 : _GEN_2376; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2700 = unuse_way == 3'h4 ? tag_1_5 : _GEN_2377; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2701 = unuse_way == 3'h4 ? tag_1_6 : _GEN_2378; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2702 = unuse_way == 3'h4 ? tag_1_7 : _GEN_2379; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2703 = unuse_way == 3'h4 ? tag_1_8 : _GEN_2380; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2704 = unuse_way == 3'h4 ? tag_1_9 : _GEN_2381; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2705 = unuse_way == 3'h4 ? tag_1_10 : _GEN_2382; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2706 = unuse_way == 3'h4 ? tag_1_11 : _GEN_2383; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2707 = unuse_way == 3'h4 ? tag_1_12 : _GEN_2384; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2708 = unuse_way == 3'h4 ? tag_1_13 : _GEN_2385; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2709 = unuse_way == 3'h4 ? tag_1_14 : _GEN_2386; // @[d_cache.scala 168:40 25:24]
  wire [31:0] _GEN_2710 = unuse_way == 3'h4 ? tag_1_15 : _GEN_2387; // @[d_cache.scala 168:40 25:24]
  wire  _GEN_2711 = unuse_way == 3'h4 ? dirty_1_0 : _GEN_2388; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2712 = unuse_way == 3'h4 ? dirty_1_1 : _GEN_2389; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2713 = unuse_way == 3'h4 ? dirty_1_2 : _GEN_2390; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2714 = unuse_way == 3'h4 ? dirty_1_3 : _GEN_2391; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2715 = unuse_way == 3'h4 ? dirty_1_4 : _GEN_2392; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2716 = unuse_way == 3'h4 ? dirty_1_5 : _GEN_2393; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2717 = unuse_way == 3'h4 ? dirty_1_6 : _GEN_2394; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2718 = unuse_way == 3'h4 ? dirty_1_7 : _GEN_2395; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2719 = unuse_way == 3'h4 ? dirty_1_8 : _GEN_2396; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2720 = unuse_way == 3'h4 ? dirty_1_9 : _GEN_2397; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2721 = unuse_way == 3'h4 ? dirty_1_10 : _GEN_2398; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2722 = unuse_way == 3'h4 ? dirty_1_11 : _GEN_2399; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2723 = unuse_way == 3'h4 ? dirty_1_12 : _GEN_2400; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2724 = unuse_way == 3'h4 ? dirty_1_13 : _GEN_2401; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2725 = unuse_way == 3'h4 ? dirty_1_14 : _GEN_2402; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2726 = unuse_way == 3'h4 ? dirty_1_15 : _GEN_2403; // @[d_cache.scala 168:40 35:26]
  wire  _GEN_2727 = unuse_way == 3'h4 ? valid_1_0 : _GEN_2404; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2728 = unuse_way == 3'h4 ? valid_1_1 : _GEN_2405; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2729 = unuse_way == 3'h4 ? valid_1_2 : _GEN_2406; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2730 = unuse_way == 3'h4 ? valid_1_3 : _GEN_2407; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2731 = unuse_way == 3'h4 ? valid_1_4 : _GEN_2408; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2732 = unuse_way == 3'h4 ? valid_1_5 : _GEN_2409; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2733 = unuse_way == 3'h4 ? valid_1_6 : _GEN_2410; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2734 = unuse_way == 3'h4 ? valid_1_7 : _GEN_2411; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2735 = unuse_way == 3'h4 ? valid_1_8 : _GEN_2412; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2736 = unuse_way == 3'h4 ? valid_1_9 : _GEN_2413; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2737 = unuse_way == 3'h4 ? valid_1_10 : _GEN_2414; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2738 = unuse_way == 3'h4 ? valid_1_11 : _GEN_2415; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2739 = unuse_way == 3'h4 ? valid_1_12 : _GEN_2416; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2740 = unuse_way == 3'h4 ? valid_1_13 : _GEN_2417; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2741 = unuse_way == 3'h4 ? valid_1_14 : _GEN_2418; // @[d_cache.scala 168:40 30:26]
  wire  _GEN_2742 = unuse_way == 3'h4 ? valid_1_15 : _GEN_2419; // @[d_cache.scala 168:40 30:26]
  wire [511:0] _GEN_2743 = unuse_way == 3'h4 ? ram_2_0 : _GEN_2420; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2744 = unuse_way == 3'h4 ? ram_2_1 : _GEN_2421; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2745 = unuse_way == 3'h4 ? ram_2_2 : _GEN_2422; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2746 = unuse_way == 3'h4 ? ram_2_3 : _GEN_2423; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2747 = unuse_way == 3'h4 ? ram_2_4 : _GEN_2424; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2748 = unuse_way == 3'h4 ? ram_2_5 : _GEN_2425; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2749 = unuse_way == 3'h4 ? ram_2_6 : _GEN_2426; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2750 = unuse_way == 3'h4 ? ram_2_7 : _GEN_2427; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2751 = unuse_way == 3'h4 ? ram_2_8 : _GEN_2428; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2752 = unuse_way == 3'h4 ? ram_2_9 : _GEN_2429; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2753 = unuse_way == 3'h4 ? ram_2_10 : _GEN_2430; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2754 = unuse_way == 3'h4 ? ram_2_11 : _GEN_2431; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2755 = unuse_way == 3'h4 ? ram_2_12 : _GEN_2432; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2756 = unuse_way == 3'h4 ? ram_2_13 : _GEN_2433; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2757 = unuse_way == 3'h4 ? ram_2_14 : _GEN_2434; // @[d_cache.scala 168:40 21:24]
  wire [511:0] _GEN_2758 = unuse_way == 3'h4 ? ram_2_15 : _GEN_2435; // @[d_cache.scala 168:40 21:24]
  wire [31:0] _GEN_2759 = unuse_way == 3'h4 ? tag_2_0 : _GEN_2436; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2760 = unuse_way == 3'h4 ? tag_2_1 : _GEN_2437; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2761 = unuse_way == 3'h4 ? tag_2_2 : _GEN_2438; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2762 = unuse_way == 3'h4 ? tag_2_3 : _GEN_2439; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2763 = unuse_way == 3'h4 ? tag_2_4 : _GEN_2440; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2764 = unuse_way == 3'h4 ? tag_2_5 : _GEN_2441; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2765 = unuse_way == 3'h4 ? tag_2_6 : _GEN_2442; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2766 = unuse_way == 3'h4 ? tag_2_7 : _GEN_2443; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2767 = unuse_way == 3'h4 ? tag_2_8 : _GEN_2444; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2768 = unuse_way == 3'h4 ? tag_2_9 : _GEN_2445; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2769 = unuse_way == 3'h4 ? tag_2_10 : _GEN_2446; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2770 = unuse_way == 3'h4 ? tag_2_11 : _GEN_2447; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2771 = unuse_way == 3'h4 ? tag_2_12 : _GEN_2448; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2772 = unuse_way == 3'h4 ? tag_2_13 : _GEN_2449; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2773 = unuse_way == 3'h4 ? tag_2_14 : _GEN_2450; // @[d_cache.scala 168:40 26:24]
  wire [31:0] _GEN_2774 = unuse_way == 3'h4 ? tag_2_15 : _GEN_2451; // @[d_cache.scala 168:40 26:24]
  wire  _GEN_2775 = unuse_way == 3'h4 ? dirty_2_0 : _GEN_2452; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2776 = unuse_way == 3'h4 ? dirty_2_1 : _GEN_2453; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2777 = unuse_way == 3'h4 ? dirty_2_2 : _GEN_2454; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2778 = unuse_way == 3'h4 ? dirty_2_3 : _GEN_2455; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2779 = unuse_way == 3'h4 ? dirty_2_4 : _GEN_2456; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2780 = unuse_way == 3'h4 ? dirty_2_5 : _GEN_2457; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2781 = unuse_way == 3'h4 ? dirty_2_6 : _GEN_2458; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2782 = unuse_way == 3'h4 ? dirty_2_7 : _GEN_2459; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2783 = unuse_way == 3'h4 ? dirty_2_8 : _GEN_2460; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2784 = unuse_way == 3'h4 ? dirty_2_9 : _GEN_2461; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2785 = unuse_way == 3'h4 ? dirty_2_10 : _GEN_2462; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2786 = unuse_way == 3'h4 ? dirty_2_11 : _GEN_2463; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2787 = unuse_way == 3'h4 ? dirty_2_12 : _GEN_2464; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2788 = unuse_way == 3'h4 ? dirty_2_13 : _GEN_2465; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2789 = unuse_way == 3'h4 ? dirty_2_14 : _GEN_2466; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2790 = unuse_way == 3'h4 ? dirty_2_15 : _GEN_2467; // @[d_cache.scala 168:40 36:26]
  wire  _GEN_2791 = unuse_way == 3'h4 ? valid_2_0 : _GEN_2468; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2792 = unuse_way == 3'h4 ? valid_2_1 : _GEN_2469; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2793 = unuse_way == 3'h4 ? valid_2_2 : _GEN_2470; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2794 = unuse_way == 3'h4 ? valid_2_3 : _GEN_2471; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2795 = unuse_way == 3'h4 ? valid_2_4 : _GEN_2472; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2796 = unuse_way == 3'h4 ? valid_2_5 : _GEN_2473; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2797 = unuse_way == 3'h4 ? valid_2_6 : _GEN_2474; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2798 = unuse_way == 3'h4 ? valid_2_7 : _GEN_2475; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2799 = unuse_way == 3'h4 ? valid_2_8 : _GEN_2476; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2800 = unuse_way == 3'h4 ? valid_2_9 : _GEN_2477; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2801 = unuse_way == 3'h4 ? valid_2_10 : _GEN_2478; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2802 = unuse_way == 3'h4 ? valid_2_11 : _GEN_2479; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2803 = unuse_way == 3'h4 ? valid_2_12 : _GEN_2480; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2804 = unuse_way == 3'h4 ? valid_2_13 : _GEN_2481; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2805 = unuse_way == 3'h4 ? valid_2_14 : _GEN_2482; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2806 = unuse_way == 3'h4 ? valid_2_15 : _GEN_2483; // @[d_cache.scala 168:40 31:26]
  wire  _GEN_2807 = unuse_way == 3'h4 ? dirty_3_0 : _GEN_2516; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2808 = unuse_way == 3'h4 ? dirty_3_1 : _GEN_2517; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2809 = unuse_way == 3'h4 ? dirty_3_2 : _GEN_2518; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2810 = unuse_way == 3'h4 ? dirty_3_3 : _GEN_2519; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2811 = unuse_way == 3'h4 ? dirty_3_4 : _GEN_2520; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2812 = unuse_way == 3'h4 ? dirty_3_5 : _GEN_2521; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2813 = unuse_way == 3'h4 ? dirty_3_6 : _GEN_2522; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2814 = unuse_way == 3'h4 ? dirty_3_7 : _GEN_2523; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2815 = unuse_way == 3'h4 ? dirty_3_8 : _GEN_2524; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2816 = unuse_way == 3'h4 ? dirty_3_9 : _GEN_2525; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2817 = unuse_way == 3'h4 ? dirty_3_10 : _GEN_2526; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2818 = unuse_way == 3'h4 ? dirty_3_11 : _GEN_2527; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2819 = unuse_way == 3'h4 ? dirty_3_12 : _GEN_2528; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2820 = unuse_way == 3'h4 ? dirty_3_13 : _GEN_2529; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2821 = unuse_way == 3'h4 ? dirty_3_14 : _GEN_2530; // @[d_cache.scala 168:40 37:26]
  wire  _GEN_2822 = unuse_way == 3'h4 ? dirty_3_15 : _GEN_2531; // @[d_cache.scala 168:40 37:26]
  wire [3:0] _GEN_2823 = unuse_way == 3'h3 ? 4'h1 : _GEN_2548; // @[d_cache.scala 162:40 163:23]
  wire [511:0] _GEN_2824 = unuse_way == 3'h3 ? _GEN_815 : _GEN_2743; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2825 = unuse_way == 3'h3 ? _GEN_816 : _GEN_2744; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2826 = unuse_way == 3'h3 ? _GEN_817 : _GEN_2745; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2827 = unuse_way == 3'h3 ? _GEN_818 : _GEN_2746; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2828 = unuse_way == 3'h3 ? _GEN_819 : _GEN_2747; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2829 = unuse_way == 3'h3 ? _GEN_820 : _GEN_2748; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2830 = unuse_way == 3'h3 ? _GEN_821 : _GEN_2749; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2831 = unuse_way == 3'h3 ? _GEN_822 : _GEN_2750; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2832 = unuse_way == 3'h3 ? _GEN_823 : _GEN_2751; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2833 = unuse_way == 3'h3 ? _GEN_824 : _GEN_2752; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2834 = unuse_way == 3'h3 ? _GEN_825 : _GEN_2753; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2835 = unuse_way == 3'h3 ? _GEN_826 : _GEN_2754; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2836 = unuse_way == 3'h3 ? _GEN_827 : _GEN_2755; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2837 = unuse_way == 3'h3 ? _GEN_828 : _GEN_2756; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2838 = unuse_way == 3'h3 ? _GEN_829 : _GEN_2757; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2839 = unuse_way == 3'h3 ? _GEN_830 : _GEN_2758; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2840 = unuse_way == 3'h3 ? _GEN_831 : _GEN_2759; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2841 = unuse_way == 3'h3 ? _GEN_832 : _GEN_2760; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2842 = unuse_way == 3'h3 ? _GEN_833 : _GEN_2761; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2843 = unuse_way == 3'h3 ? _GEN_834 : _GEN_2762; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2844 = unuse_way == 3'h3 ? _GEN_835 : _GEN_2763; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2845 = unuse_way == 3'h3 ? _GEN_836 : _GEN_2764; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2846 = unuse_way == 3'h3 ? _GEN_837 : _GEN_2765; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2847 = unuse_way == 3'h3 ? _GEN_838 : _GEN_2766; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2848 = unuse_way == 3'h3 ? _GEN_839 : _GEN_2767; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2849 = unuse_way == 3'h3 ? _GEN_840 : _GEN_2768; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2850 = unuse_way == 3'h3 ? _GEN_841 : _GEN_2769; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2851 = unuse_way == 3'h3 ? _GEN_842 : _GEN_2770; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2852 = unuse_way == 3'h3 ? _GEN_843 : _GEN_2771; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2853 = unuse_way == 3'h3 ? _GEN_844 : _GEN_2772; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2854 = unuse_way == 3'h3 ? _GEN_845 : _GEN_2773; // @[d_cache.scala 162:40]
  wire [31:0] _GEN_2855 = unuse_way == 3'h3 ? _GEN_846 : _GEN_2774; // @[d_cache.scala 162:40]
  wire  _GEN_2856 = unuse_way == 3'h3 ? _GEN_847 : _GEN_2791; // @[d_cache.scala 162:40]
  wire  _GEN_2857 = unuse_way == 3'h3 ? _GEN_848 : _GEN_2792; // @[d_cache.scala 162:40]
  wire  _GEN_2858 = unuse_way == 3'h3 ? _GEN_849 : _GEN_2793; // @[d_cache.scala 162:40]
  wire  _GEN_2859 = unuse_way == 3'h3 ? _GEN_850 : _GEN_2794; // @[d_cache.scala 162:40]
  wire  _GEN_2860 = unuse_way == 3'h3 ? _GEN_851 : _GEN_2795; // @[d_cache.scala 162:40]
  wire  _GEN_2861 = unuse_way == 3'h3 ? _GEN_852 : _GEN_2796; // @[d_cache.scala 162:40]
  wire  _GEN_2862 = unuse_way == 3'h3 ? _GEN_853 : _GEN_2797; // @[d_cache.scala 162:40]
  wire  _GEN_2863 = unuse_way == 3'h3 ? _GEN_854 : _GEN_2798; // @[d_cache.scala 162:40]
  wire  _GEN_2864 = unuse_way == 3'h3 ? _GEN_855 : _GEN_2799; // @[d_cache.scala 162:40]
  wire  _GEN_2865 = unuse_way == 3'h3 ? _GEN_856 : _GEN_2800; // @[d_cache.scala 162:40]
  wire  _GEN_2866 = unuse_way == 3'h3 ? _GEN_857 : _GEN_2801; // @[d_cache.scala 162:40]
  wire  _GEN_2867 = unuse_way == 3'h3 ? _GEN_858 : _GEN_2802; // @[d_cache.scala 162:40]
  wire  _GEN_2868 = unuse_way == 3'h3 ? _GEN_859 : _GEN_2803; // @[d_cache.scala 162:40]
  wire  _GEN_2869 = unuse_way == 3'h3 ? _GEN_860 : _GEN_2804; // @[d_cache.scala 162:40]
  wire  _GEN_2870 = unuse_way == 3'h3 ? _GEN_861 : _GEN_2805; // @[d_cache.scala 162:40]
  wire  _GEN_2871 = unuse_way == 3'h3 ? _GEN_862 : _GEN_2806; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2872 = unuse_way == 3'h3 ? _GEN_863 : _GEN_2597; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2873 = unuse_way == 3'h3 ? _GEN_864 : _GEN_2598; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2874 = unuse_way == 3'h3 ? _GEN_865 : _GEN_2599; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2875 = unuse_way == 3'h3 ? _GEN_866 : _GEN_2600; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2876 = unuse_way == 3'h3 ? _GEN_867 : _GEN_2601; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2877 = unuse_way == 3'h3 ? _GEN_868 : _GEN_2602; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2878 = unuse_way == 3'h3 ? _GEN_869 : _GEN_2603; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2879 = unuse_way == 3'h3 ? _GEN_870 : _GEN_2604; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2880 = unuse_way == 3'h3 ? _GEN_871 : _GEN_2605; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2881 = unuse_way == 3'h3 ? _GEN_872 : _GEN_2606; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2882 = unuse_way == 3'h3 ? _GEN_873 : _GEN_2607; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2883 = unuse_way == 3'h3 ? _GEN_874 : _GEN_2608; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2884 = unuse_way == 3'h3 ? _GEN_875 : _GEN_2609; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2885 = unuse_way == 3'h3 ? _GEN_876 : _GEN_2610; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2886 = unuse_way == 3'h3 ? _GEN_877 : _GEN_2611; // @[d_cache.scala 162:40]
  wire [7:0] _GEN_2887 = unuse_way == 3'h3 ? _GEN_878 : _GEN_2612; // @[d_cache.scala 162:40]
  wire [511:0] _GEN_2888 = unuse_way == 3'h3 ? ram_3_0 : _GEN_2549; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2889 = unuse_way == 3'h3 ? ram_3_1 : _GEN_2550; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2890 = unuse_way == 3'h3 ? ram_3_2 : _GEN_2551; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2891 = unuse_way == 3'h3 ? ram_3_3 : _GEN_2552; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2892 = unuse_way == 3'h3 ? ram_3_4 : _GEN_2553; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2893 = unuse_way == 3'h3 ? ram_3_5 : _GEN_2554; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2894 = unuse_way == 3'h3 ? ram_3_6 : _GEN_2555; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2895 = unuse_way == 3'h3 ? ram_3_7 : _GEN_2556; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2896 = unuse_way == 3'h3 ? ram_3_8 : _GEN_2557; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2897 = unuse_way == 3'h3 ? ram_3_9 : _GEN_2558; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2898 = unuse_way == 3'h3 ? ram_3_10 : _GEN_2559; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2899 = unuse_way == 3'h3 ? ram_3_11 : _GEN_2560; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2900 = unuse_way == 3'h3 ? ram_3_12 : _GEN_2561; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2901 = unuse_way == 3'h3 ? ram_3_13 : _GEN_2562; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2902 = unuse_way == 3'h3 ? ram_3_14 : _GEN_2563; // @[d_cache.scala 162:40 22:24]
  wire [511:0] _GEN_2903 = unuse_way == 3'h3 ? ram_3_15 : _GEN_2564; // @[d_cache.scala 162:40 22:24]
  wire [31:0] _GEN_2904 = unuse_way == 3'h3 ? tag_3_0 : _GEN_2565; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2905 = unuse_way == 3'h3 ? tag_3_1 : _GEN_2566; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2906 = unuse_way == 3'h3 ? tag_3_2 : _GEN_2567; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2907 = unuse_way == 3'h3 ? tag_3_3 : _GEN_2568; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2908 = unuse_way == 3'h3 ? tag_3_4 : _GEN_2569; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2909 = unuse_way == 3'h3 ? tag_3_5 : _GEN_2570; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2910 = unuse_way == 3'h3 ? tag_3_6 : _GEN_2571; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2911 = unuse_way == 3'h3 ? tag_3_7 : _GEN_2572; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2912 = unuse_way == 3'h3 ? tag_3_8 : _GEN_2573; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2913 = unuse_way == 3'h3 ? tag_3_9 : _GEN_2574; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2914 = unuse_way == 3'h3 ? tag_3_10 : _GEN_2575; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2915 = unuse_way == 3'h3 ? tag_3_11 : _GEN_2576; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2916 = unuse_way == 3'h3 ? tag_3_12 : _GEN_2577; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2917 = unuse_way == 3'h3 ? tag_3_13 : _GEN_2578; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2918 = unuse_way == 3'h3 ? tag_3_14 : _GEN_2579; // @[d_cache.scala 162:40 27:24]
  wire [31:0] _GEN_2919 = unuse_way == 3'h3 ? tag_3_15 : _GEN_2580; // @[d_cache.scala 162:40 27:24]
  wire  _GEN_2920 = unuse_way == 3'h3 ? valid_3_0 : _GEN_2581; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2921 = unuse_way == 3'h3 ? valid_3_1 : _GEN_2582; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2922 = unuse_way == 3'h3 ? valid_3_2 : _GEN_2583; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2923 = unuse_way == 3'h3 ? valid_3_3 : _GEN_2584; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2924 = unuse_way == 3'h3 ? valid_3_4 : _GEN_2585; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2925 = unuse_way == 3'h3 ? valid_3_5 : _GEN_2586; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2926 = unuse_way == 3'h3 ? valid_3_6 : _GEN_2587; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2927 = unuse_way == 3'h3 ? valid_3_7 : _GEN_2588; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2928 = unuse_way == 3'h3 ? valid_3_8 : _GEN_2589; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2929 = unuse_way == 3'h3 ? valid_3_9 : _GEN_2590; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2930 = unuse_way == 3'h3 ? valid_3_10 : _GEN_2591; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2931 = unuse_way == 3'h3 ? valid_3_11 : _GEN_2592; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2932 = unuse_way == 3'h3 ? valid_3_12 : _GEN_2593; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2933 = unuse_way == 3'h3 ? valid_3_13 : _GEN_2594; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2934 = unuse_way == 3'h3 ? valid_3_14 : _GEN_2595; // @[d_cache.scala 162:40 32:26]
  wire  _GEN_2935 = unuse_way == 3'h3 ? valid_3_15 : _GEN_2596; // @[d_cache.scala 162:40 32:26]
  wire [511:0] _GEN_2936 = unuse_way == 3'h3 ? write_back_data : _GEN_2613; // @[d_cache.scala 162:40 44:34]
  wire [41:0] _GEN_2937 = unuse_way == 3'h3 ? {{10'd0}, write_back_addr} : _GEN_2614; // @[d_cache.scala 162:40 45:34]
  wire [511:0] _GEN_2938 = unuse_way == 3'h3 ? ram_0_0 : _GEN_2615; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2939 = unuse_way == 3'h3 ? ram_0_1 : _GEN_2616; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2940 = unuse_way == 3'h3 ? ram_0_2 : _GEN_2617; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2941 = unuse_way == 3'h3 ? ram_0_3 : _GEN_2618; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2942 = unuse_way == 3'h3 ? ram_0_4 : _GEN_2619; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2943 = unuse_way == 3'h3 ? ram_0_5 : _GEN_2620; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2944 = unuse_way == 3'h3 ? ram_0_6 : _GEN_2621; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2945 = unuse_way == 3'h3 ? ram_0_7 : _GEN_2622; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2946 = unuse_way == 3'h3 ? ram_0_8 : _GEN_2623; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2947 = unuse_way == 3'h3 ? ram_0_9 : _GEN_2624; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2948 = unuse_way == 3'h3 ? ram_0_10 : _GEN_2625; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2949 = unuse_way == 3'h3 ? ram_0_11 : _GEN_2626; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2950 = unuse_way == 3'h3 ? ram_0_12 : _GEN_2627; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2951 = unuse_way == 3'h3 ? ram_0_13 : _GEN_2628; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2952 = unuse_way == 3'h3 ? ram_0_14 : _GEN_2629; // @[d_cache.scala 162:40 19:24]
  wire [511:0] _GEN_2953 = unuse_way == 3'h3 ? ram_0_15 : _GEN_2630; // @[d_cache.scala 162:40 19:24]
  wire [31:0] _GEN_2954 = unuse_way == 3'h3 ? tag_0_0 : _GEN_2631; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2955 = unuse_way == 3'h3 ? tag_0_1 : _GEN_2632; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2956 = unuse_way == 3'h3 ? tag_0_2 : _GEN_2633; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2957 = unuse_way == 3'h3 ? tag_0_3 : _GEN_2634; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2958 = unuse_way == 3'h3 ? tag_0_4 : _GEN_2635; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2959 = unuse_way == 3'h3 ? tag_0_5 : _GEN_2636; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2960 = unuse_way == 3'h3 ? tag_0_6 : _GEN_2637; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2961 = unuse_way == 3'h3 ? tag_0_7 : _GEN_2638; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2962 = unuse_way == 3'h3 ? tag_0_8 : _GEN_2639; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2963 = unuse_way == 3'h3 ? tag_0_9 : _GEN_2640; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2964 = unuse_way == 3'h3 ? tag_0_10 : _GEN_2641; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2965 = unuse_way == 3'h3 ? tag_0_11 : _GEN_2642; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2966 = unuse_way == 3'h3 ? tag_0_12 : _GEN_2643; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2967 = unuse_way == 3'h3 ? tag_0_13 : _GEN_2644; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2968 = unuse_way == 3'h3 ? tag_0_14 : _GEN_2645; // @[d_cache.scala 162:40 24:24]
  wire [31:0] _GEN_2969 = unuse_way == 3'h3 ? tag_0_15 : _GEN_2646; // @[d_cache.scala 162:40 24:24]
  wire  _GEN_2970 = unuse_way == 3'h3 ? dirty_0_0 : _GEN_2647; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2971 = unuse_way == 3'h3 ? dirty_0_1 : _GEN_2648; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2972 = unuse_way == 3'h3 ? dirty_0_2 : _GEN_2649; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2973 = unuse_way == 3'h3 ? dirty_0_3 : _GEN_2650; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2974 = unuse_way == 3'h3 ? dirty_0_4 : _GEN_2651; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2975 = unuse_way == 3'h3 ? dirty_0_5 : _GEN_2652; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2976 = unuse_way == 3'h3 ? dirty_0_6 : _GEN_2653; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2977 = unuse_way == 3'h3 ? dirty_0_7 : _GEN_2654; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2978 = unuse_way == 3'h3 ? dirty_0_8 : _GEN_2655; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2979 = unuse_way == 3'h3 ? dirty_0_9 : _GEN_2656; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2980 = unuse_way == 3'h3 ? dirty_0_10 : _GEN_2657; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2981 = unuse_way == 3'h3 ? dirty_0_11 : _GEN_2658; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2982 = unuse_way == 3'h3 ? dirty_0_12 : _GEN_2659; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2983 = unuse_way == 3'h3 ? dirty_0_13 : _GEN_2660; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2984 = unuse_way == 3'h3 ? dirty_0_14 : _GEN_2661; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2985 = unuse_way == 3'h3 ? dirty_0_15 : _GEN_2662; // @[d_cache.scala 162:40 34:26]
  wire  _GEN_2986 = unuse_way == 3'h3 ? valid_0_0 : _GEN_2663; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2987 = unuse_way == 3'h3 ? valid_0_1 : _GEN_2664; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2988 = unuse_way == 3'h3 ? valid_0_2 : _GEN_2665; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2989 = unuse_way == 3'h3 ? valid_0_3 : _GEN_2666; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2990 = unuse_way == 3'h3 ? valid_0_4 : _GEN_2667; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2991 = unuse_way == 3'h3 ? valid_0_5 : _GEN_2668; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2992 = unuse_way == 3'h3 ? valid_0_6 : _GEN_2669; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2993 = unuse_way == 3'h3 ? valid_0_7 : _GEN_2670; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2994 = unuse_way == 3'h3 ? valid_0_8 : _GEN_2671; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2995 = unuse_way == 3'h3 ? valid_0_9 : _GEN_2672; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2996 = unuse_way == 3'h3 ? valid_0_10 : _GEN_2673; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2997 = unuse_way == 3'h3 ? valid_0_11 : _GEN_2674; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2998 = unuse_way == 3'h3 ? valid_0_12 : _GEN_2675; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_2999 = unuse_way == 3'h3 ? valid_0_13 : _GEN_2676; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_3000 = unuse_way == 3'h3 ? valid_0_14 : _GEN_2677; // @[d_cache.scala 162:40 29:26]
  wire  _GEN_3001 = unuse_way == 3'h3 ? valid_0_15 : _GEN_2678; // @[d_cache.scala 162:40 29:26]
  wire [511:0] _GEN_3002 = unuse_way == 3'h3 ? ram_1_0 : _GEN_2679; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3003 = unuse_way == 3'h3 ? ram_1_1 : _GEN_2680; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3004 = unuse_way == 3'h3 ? ram_1_2 : _GEN_2681; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3005 = unuse_way == 3'h3 ? ram_1_3 : _GEN_2682; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3006 = unuse_way == 3'h3 ? ram_1_4 : _GEN_2683; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3007 = unuse_way == 3'h3 ? ram_1_5 : _GEN_2684; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3008 = unuse_way == 3'h3 ? ram_1_6 : _GEN_2685; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3009 = unuse_way == 3'h3 ? ram_1_7 : _GEN_2686; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3010 = unuse_way == 3'h3 ? ram_1_8 : _GEN_2687; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3011 = unuse_way == 3'h3 ? ram_1_9 : _GEN_2688; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3012 = unuse_way == 3'h3 ? ram_1_10 : _GEN_2689; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3013 = unuse_way == 3'h3 ? ram_1_11 : _GEN_2690; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3014 = unuse_way == 3'h3 ? ram_1_12 : _GEN_2691; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3015 = unuse_way == 3'h3 ? ram_1_13 : _GEN_2692; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3016 = unuse_way == 3'h3 ? ram_1_14 : _GEN_2693; // @[d_cache.scala 162:40 20:24]
  wire [511:0] _GEN_3017 = unuse_way == 3'h3 ? ram_1_15 : _GEN_2694; // @[d_cache.scala 162:40 20:24]
  wire [31:0] _GEN_3018 = unuse_way == 3'h3 ? tag_1_0 : _GEN_2695; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3019 = unuse_way == 3'h3 ? tag_1_1 : _GEN_2696; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3020 = unuse_way == 3'h3 ? tag_1_2 : _GEN_2697; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3021 = unuse_way == 3'h3 ? tag_1_3 : _GEN_2698; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3022 = unuse_way == 3'h3 ? tag_1_4 : _GEN_2699; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3023 = unuse_way == 3'h3 ? tag_1_5 : _GEN_2700; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3024 = unuse_way == 3'h3 ? tag_1_6 : _GEN_2701; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3025 = unuse_way == 3'h3 ? tag_1_7 : _GEN_2702; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3026 = unuse_way == 3'h3 ? tag_1_8 : _GEN_2703; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3027 = unuse_way == 3'h3 ? tag_1_9 : _GEN_2704; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3028 = unuse_way == 3'h3 ? tag_1_10 : _GEN_2705; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3029 = unuse_way == 3'h3 ? tag_1_11 : _GEN_2706; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3030 = unuse_way == 3'h3 ? tag_1_12 : _GEN_2707; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3031 = unuse_way == 3'h3 ? tag_1_13 : _GEN_2708; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3032 = unuse_way == 3'h3 ? tag_1_14 : _GEN_2709; // @[d_cache.scala 162:40 25:24]
  wire [31:0] _GEN_3033 = unuse_way == 3'h3 ? tag_1_15 : _GEN_2710; // @[d_cache.scala 162:40 25:24]
  wire  _GEN_3034 = unuse_way == 3'h3 ? dirty_1_0 : _GEN_2711; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3035 = unuse_way == 3'h3 ? dirty_1_1 : _GEN_2712; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3036 = unuse_way == 3'h3 ? dirty_1_2 : _GEN_2713; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3037 = unuse_way == 3'h3 ? dirty_1_3 : _GEN_2714; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3038 = unuse_way == 3'h3 ? dirty_1_4 : _GEN_2715; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3039 = unuse_way == 3'h3 ? dirty_1_5 : _GEN_2716; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3040 = unuse_way == 3'h3 ? dirty_1_6 : _GEN_2717; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3041 = unuse_way == 3'h3 ? dirty_1_7 : _GEN_2718; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3042 = unuse_way == 3'h3 ? dirty_1_8 : _GEN_2719; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3043 = unuse_way == 3'h3 ? dirty_1_9 : _GEN_2720; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3044 = unuse_way == 3'h3 ? dirty_1_10 : _GEN_2721; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3045 = unuse_way == 3'h3 ? dirty_1_11 : _GEN_2722; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3046 = unuse_way == 3'h3 ? dirty_1_12 : _GEN_2723; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3047 = unuse_way == 3'h3 ? dirty_1_13 : _GEN_2724; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3048 = unuse_way == 3'h3 ? dirty_1_14 : _GEN_2725; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3049 = unuse_way == 3'h3 ? dirty_1_15 : _GEN_2726; // @[d_cache.scala 162:40 35:26]
  wire  _GEN_3050 = unuse_way == 3'h3 ? valid_1_0 : _GEN_2727; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3051 = unuse_way == 3'h3 ? valid_1_1 : _GEN_2728; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3052 = unuse_way == 3'h3 ? valid_1_2 : _GEN_2729; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3053 = unuse_way == 3'h3 ? valid_1_3 : _GEN_2730; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3054 = unuse_way == 3'h3 ? valid_1_4 : _GEN_2731; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3055 = unuse_way == 3'h3 ? valid_1_5 : _GEN_2732; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3056 = unuse_way == 3'h3 ? valid_1_6 : _GEN_2733; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3057 = unuse_way == 3'h3 ? valid_1_7 : _GEN_2734; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3058 = unuse_way == 3'h3 ? valid_1_8 : _GEN_2735; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3059 = unuse_way == 3'h3 ? valid_1_9 : _GEN_2736; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3060 = unuse_way == 3'h3 ? valid_1_10 : _GEN_2737; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3061 = unuse_way == 3'h3 ? valid_1_11 : _GEN_2738; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3062 = unuse_way == 3'h3 ? valid_1_12 : _GEN_2739; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3063 = unuse_way == 3'h3 ? valid_1_13 : _GEN_2740; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3064 = unuse_way == 3'h3 ? valid_1_14 : _GEN_2741; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3065 = unuse_way == 3'h3 ? valid_1_15 : _GEN_2742; // @[d_cache.scala 162:40 30:26]
  wire  _GEN_3066 = unuse_way == 3'h3 ? dirty_2_0 : _GEN_2775; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3067 = unuse_way == 3'h3 ? dirty_2_1 : _GEN_2776; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3068 = unuse_way == 3'h3 ? dirty_2_2 : _GEN_2777; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3069 = unuse_way == 3'h3 ? dirty_2_3 : _GEN_2778; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3070 = unuse_way == 3'h3 ? dirty_2_4 : _GEN_2779; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3071 = unuse_way == 3'h3 ? dirty_2_5 : _GEN_2780; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3072 = unuse_way == 3'h3 ? dirty_2_6 : _GEN_2781; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3073 = unuse_way == 3'h3 ? dirty_2_7 : _GEN_2782; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3074 = unuse_way == 3'h3 ? dirty_2_8 : _GEN_2783; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3075 = unuse_way == 3'h3 ? dirty_2_9 : _GEN_2784; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3076 = unuse_way == 3'h3 ? dirty_2_10 : _GEN_2785; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3077 = unuse_way == 3'h3 ? dirty_2_11 : _GEN_2786; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3078 = unuse_way == 3'h3 ? dirty_2_12 : _GEN_2787; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3079 = unuse_way == 3'h3 ? dirty_2_13 : _GEN_2788; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3080 = unuse_way == 3'h3 ? dirty_2_14 : _GEN_2789; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3081 = unuse_way == 3'h3 ? dirty_2_15 : _GEN_2790; // @[d_cache.scala 162:40 36:26]
  wire  _GEN_3082 = unuse_way == 3'h3 ? dirty_3_0 : _GEN_2807; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3083 = unuse_way == 3'h3 ? dirty_3_1 : _GEN_2808; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3084 = unuse_way == 3'h3 ? dirty_3_2 : _GEN_2809; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3085 = unuse_way == 3'h3 ? dirty_3_3 : _GEN_2810; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3086 = unuse_way == 3'h3 ? dirty_3_4 : _GEN_2811; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3087 = unuse_way == 3'h3 ? dirty_3_5 : _GEN_2812; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3088 = unuse_way == 3'h3 ? dirty_3_6 : _GEN_2813; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3089 = unuse_way == 3'h3 ? dirty_3_7 : _GEN_2814; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3090 = unuse_way == 3'h3 ? dirty_3_8 : _GEN_2815; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3091 = unuse_way == 3'h3 ? dirty_3_9 : _GEN_2816; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3092 = unuse_way == 3'h3 ? dirty_3_10 : _GEN_2817; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3093 = unuse_way == 3'h3 ? dirty_3_11 : _GEN_2818; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3094 = unuse_way == 3'h3 ? dirty_3_12 : _GEN_2819; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3095 = unuse_way == 3'h3 ? dirty_3_13 : _GEN_2820; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3096 = unuse_way == 3'h3 ? dirty_3_14 : _GEN_2821; // @[d_cache.scala 162:40 37:26]
  wire  _GEN_3097 = unuse_way == 3'h3 ? dirty_3_15 : _GEN_2822; // @[d_cache.scala 162:40 37:26]
  wire [3:0] _GEN_3098 = unuse_way == 3'h2 ? 4'h1 : _GEN_2823; // @[d_cache.scala 156:40 157:23]
  wire [511:0] _GEN_3099 = unuse_way == 3'h2 ? _GEN_751 : _GEN_3002; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3100 = unuse_way == 3'h2 ? _GEN_752 : _GEN_3003; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3101 = unuse_way == 3'h2 ? _GEN_753 : _GEN_3004; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3102 = unuse_way == 3'h2 ? _GEN_754 : _GEN_3005; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3103 = unuse_way == 3'h2 ? _GEN_755 : _GEN_3006; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3104 = unuse_way == 3'h2 ? _GEN_756 : _GEN_3007; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3105 = unuse_way == 3'h2 ? _GEN_757 : _GEN_3008; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3106 = unuse_way == 3'h2 ? _GEN_758 : _GEN_3009; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3107 = unuse_way == 3'h2 ? _GEN_759 : _GEN_3010; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3108 = unuse_way == 3'h2 ? _GEN_760 : _GEN_3011; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3109 = unuse_way == 3'h2 ? _GEN_761 : _GEN_3012; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3110 = unuse_way == 3'h2 ? _GEN_762 : _GEN_3013; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3111 = unuse_way == 3'h2 ? _GEN_763 : _GEN_3014; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3112 = unuse_way == 3'h2 ? _GEN_764 : _GEN_3015; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3113 = unuse_way == 3'h2 ? _GEN_765 : _GEN_3016; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3114 = unuse_way == 3'h2 ? _GEN_766 : _GEN_3017; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3115 = unuse_way == 3'h2 ? _GEN_767 : _GEN_3018; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3116 = unuse_way == 3'h2 ? _GEN_768 : _GEN_3019; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3117 = unuse_way == 3'h2 ? _GEN_769 : _GEN_3020; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3118 = unuse_way == 3'h2 ? _GEN_770 : _GEN_3021; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3119 = unuse_way == 3'h2 ? _GEN_771 : _GEN_3022; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3120 = unuse_way == 3'h2 ? _GEN_772 : _GEN_3023; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3121 = unuse_way == 3'h2 ? _GEN_773 : _GEN_3024; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3122 = unuse_way == 3'h2 ? _GEN_774 : _GEN_3025; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3123 = unuse_way == 3'h2 ? _GEN_775 : _GEN_3026; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3124 = unuse_way == 3'h2 ? _GEN_776 : _GEN_3027; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3125 = unuse_way == 3'h2 ? _GEN_777 : _GEN_3028; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3126 = unuse_way == 3'h2 ? _GEN_778 : _GEN_3029; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3127 = unuse_way == 3'h2 ? _GEN_779 : _GEN_3030; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3128 = unuse_way == 3'h2 ? _GEN_780 : _GEN_3031; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3129 = unuse_way == 3'h2 ? _GEN_781 : _GEN_3032; // @[d_cache.scala 156:40]
  wire [31:0] _GEN_3130 = unuse_way == 3'h2 ? _GEN_782 : _GEN_3033; // @[d_cache.scala 156:40]
  wire  _GEN_3131 = unuse_way == 3'h2 ? _GEN_783 : _GEN_3050; // @[d_cache.scala 156:40]
  wire  _GEN_3132 = unuse_way == 3'h2 ? _GEN_784 : _GEN_3051; // @[d_cache.scala 156:40]
  wire  _GEN_3133 = unuse_way == 3'h2 ? _GEN_785 : _GEN_3052; // @[d_cache.scala 156:40]
  wire  _GEN_3134 = unuse_way == 3'h2 ? _GEN_786 : _GEN_3053; // @[d_cache.scala 156:40]
  wire  _GEN_3135 = unuse_way == 3'h2 ? _GEN_787 : _GEN_3054; // @[d_cache.scala 156:40]
  wire  _GEN_3136 = unuse_way == 3'h2 ? _GEN_788 : _GEN_3055; // @[d_cache.scala 156:40]
  wire  _GEN_3137 = unuse_way == 3'h2 ? _GEN_789 : _GEN_3056; // @[d_cache.scala 156:40]
  wire  _GEN_3138 = unuse_way == 3'h2 ? _GEN_790 : _GEN_3057; // @[d_cache.scala 156:40]
  wire  _GEN_3139 = unuse_way == 3'h2 ? _GEN_791 : _GEN_3058; // @[d_cache.scala 156:40]
  wire  _GEN_3140 = unuse_way == 3'h2 ? _GEN_792 : _GEN_3059; // @[d_cache.scala 156:40]
  wire  _GEN_3141 = unuse_way == 3'h2 ? _GEN_793 : _GEN_3060; // @[d_cache.scala 156:40]
  wire  _GEN_3142 = unuse_way == 3'h2 ? _GEN_794 : _GEN_3061; // @[d_cache.scala 156:40]
  wire  _GEN_3143 = unuse_way == 3'h2 ? _GEN_795 : _GEN_3062; // @[d_cache.scala 156:40]
  wire  _GEN_3144 = unuse_way == 3'h2 ? _GEN_796 : _GEN_3063; // @[d_cache.scala 156:40]
  wire  _GEN_3145 = unuse_way == 3'h2 ? _GEN_797 : _GEN_3064; // @[d_cache.scala 156:40]
  wire  _GEN_3146 = unuse_way == 3'h2 ? _GEN_798 : _GEN_3065; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3147 = unuse_way == 3'h2 ? _GEN_799 : _GEN_2872; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3148 = unuse_way == 3'h2 ? _GEN_800 : _GEN_2873; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3149 = unuse_way == 3'h2 ? _GEN_801 : _GEN_2874; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3150 = unuse_way == 3'h2 ? _GEN_802 : _GEN_2875; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3151 = unuse_way == 3'h2 ? _GEN_803 : _GEN_2876; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3152 = unuse_way == 3'h2 ? _GEN_804 : _GEN_2877; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3153 = unuse_way == 3'h2 ? _GEN_805 : _GEN_2878; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3154 = unuse_way == 3'h2 ? _GEN_806 : _GEN_2879; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3155 = unuse_way == 3'h2 ? _GEN_807 : _GEN_2880; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3156 = unuse_way == 3'h2 ? _GEN_808 : _GEN_2881; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3157 = unuse_way == 3'h2 ? _GEN_809 : _GEN_2882; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3158 = unuse_way == 3'h2 ? _GEN_810 : _GEN_2883; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3159 = unuse_way == 3'h2 ? _GEN_811 : _GEN_2884; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3160 = unuse_way == 3'h2 ? _GEN_812 : _GEN_2885; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3161 = unuse_way == 3'h2 ? _GEN_813 : _GEN_2886; // @[d_cache.scala 156:40]
  wire [7:0] _GEN_3162 = unuse_way == 3'h2 ? _GEN_814 : _GEN_2887; // @[d_cache.scala 156:40]
  wire [511:0] _GEN_3163 = unuse_way == 3'h2 ? ram_2_0 : _GEN_2824; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3164 = unuse_way == 3'h2 ? ram_2_1 : _GEN_2825; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3165 = unuse_way == 3'h2 ? ram_2_2 : _GEN_2826; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3166 = unuse_way == 3'h2 ? ram_2_3 : _GEN_2827; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3167 = unuse_way == 3'h2 ? ram_2_4 : _GEN_2828; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3168 = unuse_way == 3'h2 ? ram_2_5 : _GEN_2829; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3169 = unuse_way == 3'h2 ? ram_2_6 : _GEN_2830; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3170 = unuse_way == 3'h2 ? ram_2_7 : _GEN_2831; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3171 = unuse_way == 3'h2 ? ram_2_8 : _GEN_2832; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3172 = unuse_way == 3'h2 ? ram_2_9 : _GEN_2833; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3173 = unuse_way == 3'h2 ? ram_2_10 : _GEN_2834; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3174 = unuse_way == 3'h2 ? ram_2_11 : _GEN_2835; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3175 = unuse_way == 3'h2 ? ram_2_12 : _GEN_2836; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3176 = unuse_way == 3'h2 ? ram_2_13 : _GEN_2837; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3177 = unuse_way == 3'h2 ? ram_2_14 : _GEN_2838; // @[d_cache.scala 156:40 21:24]
  wire [511:0] _GEN_3178 = unuse_way == 3'h2 ? ram_2_15 : _GEN_2839; // @[d_cache.scala 156:40 21:24]
  wire [31:0] _GEN_3179 = unuse_way == 3'h2 ? tag_2_0 : _GEN_2840; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3180 = unuse_way == 3'h2 ? tag_2_1 : _GEN_2841; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3181 = unuse_way == 3'h2 ? tag_2_2 : _GEN_2842; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3182 = unuse_way == 3'h2 ? tag_2_3 : _GEN_2843; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3183 = unuse_way == 3'h2 ? tag_2_4 : _GEN_2844; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3184 = unuse_way == 3'h2 ? tag_2_5 : _GEN_2845; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3185 = unuse_way == 3'h2 ? tag_2_6 : _GEN_2846; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3186 = unuse_way == 3'h2 ? tag_2_7 : _GEN_2847; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3187 = unuse_way == 3'h2 ? tag_2_8 : _GEN_2848; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3188 = unuse_way == 3'h2 ? tag_2_9 : _GEN_2849; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3189 = unuse_way == 3'h2 ? tag_2_10 : _GEN_2850; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3190 = unuse_way == 3'h2 ? tag_2_11 : _GEN_2851; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3191 = unuse_way == 3'h2 ? tag_2_12 : _GEN_2852; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3192 = unuse_way == 3'h2 ? tag_2_13 : _GEN_2853; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3193 = unuse_way == 3'h2 ? tag_2_14 : _GEN_2854; // @[d_cache.scala 156:40 26:24]
  wire [31:0] _GEN_3194 = unuse_way == 3'h2 ? tag_2_15 : _GEN_2855; // @[d_cache.scala 156:40 26:24]
  wire  _GEN_3195 = unuse_way == 3'h2 ? valid_2_0 : _GEN_2856; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3196 = unuse_way == 3'h2 ? valid_2_1 : _GEN_2857; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3197 = unuse_way == 3'h2 ? valid_2_2 : _GEN_2858; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3198 = unuse_way == 3'h2 ? valid_2_3 : _GEN_2859; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3199 = unuse_way == 3'h2 ? valid_2_4 : _GEN_2860; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3200 = unuse_way == 3'h2 ? valid_2_5 : _GEN_2861; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3201 = unuse_way == 3'h2 ? valid_2_6 : _GEN_2862; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3202 = unuse_way == 3'h2 ? valid_2_7 : _GEN_2863; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3203 = unuse_way == 3'h2 ? valid_2_8 : _GEN_2864; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3204 = unuse_way == 3'h2 ? valid_2_9 : _GEN_2865; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3205 = unuse_way == 3'h2 ? valid_2_10 : _GEN_2866; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3206 = unuse_way == 3'h2 ? valid_2_11 : _GEN_2867; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3207 = unuse_way == 3'h2 ? valid_2_12 : _GEN_2868; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3208 = unuse_way == 3'h2 ? valid_2_13 : _GEN_2869; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3209 = unuse_way == 3'h2 ? valid_2_14 : _GEN_2870; // @[d_cache.scala 156:40 31:26]
  wire  _GEN_3210 = unuse_way == 3'h2 ? valid_2_15 : _GEN_2871; // @[d_cache.scala 156:40 31:26]
  wire [511:0] _GEN_3211 = unuse_way == 3'h2 ? ram_3_0 : _GEN_2888; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3212 = unuse_way == 3'h2 ? ram_3_1 : _GEN_2889; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3213 = unuse_way == 3'h2 ? ram_3_2 : _GEN_2890; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3214 = unuse_way == 3'h2 ? ram_3_3 : _GEN_2891; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3215 = unuse_way == 3'h2 ? ram_3_4 : _GEN_2892; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3216 = unuse_way == 3'h2 ? ram_3_5 : _GEN_2893; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3217 = unuse_way == 3'h2 ? ram_3_6 : _GEN_2894; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3218 = unuse_way == 3'h2 ? ram_3_7 : _GEN_2895; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3219 = unuse_way == 3'h2 ? ram_3_8 : _GEN_2896; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3220 = unuse_way == 3'h2 ? ram_3_9 : _GEN_2897; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3221 = unuse_way == 3'h2 ? ram_3_10 : _GEN_2898; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3222 = unuse_way == 3'h2 ? ram_3_11 : _GEN_2899; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3223 = unuse_way == 3'h2 ? ram_3_12 : _GEN_2900; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3224 = unuse_way == 3'h2 ? ram_3_13 : _GEN_2901; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3225 = unuse_way == 3'h2 ? ram_3_14 : _GEN_2902; // @[d_cache.scala 156:40 22:24]
  wire [511:0] _GEN_3226 = unuse_way == 3'h2 ? ram_3_15 : _GEN_2903; // @[d_cache.scala 156:40 22:24]
  wire [31:0] _GEN_3227 = unuse_way == 3'h2 ? tag_3_0 : _GEN_2904; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3228 = unuse_way == 3'h2 ? tag_3_1 : _GEN_2905; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3229 = unuse_way == 3'h2 ? tag_3_2 : _GEN_2906; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3230 = unuse_way == 3'h2 ? tag_3_3 : _GEN_2907; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3231 = unuse_way == 3'h2 ? tag_3_4 : _GEN_2908; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3232 = unuse_way == 3'h2 ? tag_3_5 : _GEN_2909; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3233 = unuse_way == 3'h2 ? tag_3_6 : _GEN_2910; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3234 = unuse_way == 3'h2 ? tag_3_7 : _GEN_2911; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3235 = unuse_way == 3'h2 ? tag_3_8 : _GEN_2912; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3236 = unuse_way == 3'h2 ? tag_3_9 : _GEN_2913; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3237 = unuse_way == 3'h2 ? tag_3_10 : _GEN_2914; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3238 = unuse_way == 3'h2 ? tag_3_11 : _GEN_2915; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3239 = unuse_way == 3'h2 ? tag_3_12 : _GEN_2916; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3240 = unuse_way == 3'h2 ? tag_3_13 : _GEN_2917; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3241 = unuse_way == 3'h2 ? tag_3_14 : _GEN_2918; // @[d_cache.scala 156:40 27:24]
  wire [31:0] _GEN_3242 = unuse_way == 3'h2 ? tag_3_15 : _GEN_2919; // @[d_cache.scala 156:40 27:24]
  wire  _GEN_3243 = unuse_way == 3'h2 ? valid_3_0 : _GEN_2920; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3244 = unuse_way == 3'h2 ? valid_3_1 : _GEN_2921; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3245 = unuse_way == 3'h2 ? valid_3_2 : _GEN_2922; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3246 = unuse_way == 3'h2 ? valid_3_3 : _GEN_2923; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3247 = unuse_way == 3'h2 ? valid_3_4 : _GEN_2924; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3248 = unuse_way == 3'h2 ? valid_3_5 : _GEN_2925; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3249 = unuse_way == 3'h2 ? valid_3_6 : _GEN_2926; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3250 = unuse_way == 3'h2 ? valid_3_7 : _GEN_2927; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3251 = unuse_way == 3'h2 ? valid_3_8 : _GEN_2928; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3252 = unuse_way == 3'h2 ? valid_3_9 : _GEN_2929; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3253 = unuse_way == 3'h2 ? valid_3_10 : _GEN_2930; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3254 = unuse_way == 3'h2 ? valid_3_11 : _GEN_2931; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3255 = unuse_way == 3'h2 ? valid_3_12 : _GEN_2932; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3256 = unuse_way == 3'h2 ? valid_3_13 : _GEN_2933; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3257 = unuse_way == 3'h2 ? valid_3_14 : _GEN_2934; // @[d_cache.scala 156:40 32:26]
  wire  _GEN_3258 = unuse_way == 3'h2 ? valid_3_15 : _GEN_2935; // @[d_cache.scala 156:40 32:26]
  wire [511:0] _GEN_3259 = unuse_way == 3'h2 ? write_back_data : _GEN_2936; // @[d_cache.scala 156:40 44:34]
  wire [41:0] _GEN_3260 = unuse_way == 3'h2 ? {{10'd0}, write_back_addr} : _GEN_2937; // @[d_cache.scala 156:40 45:34]
  wire [511:0] _GEN_3261 = unuse_way == 3'h2 ? ram_0_0 : _GEN_2938; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3262 = unuse_way == 3'h2 ? ram_0_1 : _GEN_2939; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3263 = unuse_way == 3'h2 ? ram_0_2 : _GEN_2940; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3264 = unuse_way == 3'h2 ? ram_0_3 : _GEN_2941; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3265 = unuse_way == 3'h2 ? ram_0_4 : _GEN_2942; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3266 = unuse_way == 3'h2 ? ram_0_5 : _GEN_2943; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3267 = unuse_way == 3'h2 ? ram_0_6 : _GEN_2944; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3268 = unuse_way == 3'h2 ? ram_0_7 : _GEN_2945; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3269 = unuse_way == 3'h2 ? ram_0_8 : _GEN_2946; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3270 = unuse_way == 3'h2 ? ram_0_9 : _GEN_2947; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3271 = unuse_way == 3'h2 ? ram_0_10 : _GEN_2948; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3272 = unuse_way == 3'h2 ? ram_0_11 : _GEN_2949; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3273 = unuse_way == 3'h2 ? ram_0_12 : _GEN_2950; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3274 = unuse_way == 3'h2 ? ram_0_13 : _GEN_2951; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3275 = unuse_way == 3'h2 ? ram_0_14 : _GEN_2952; // @[d_cache.scala 156:40 19:24]
  wire [511:0] _GEN_3276 = unuse_way == 3'h2 ? ram_0_15 : _GEN_2953; // @[d_cache.scala 156:40 19:24]
  wire [31:0] _GEN_3277 = unuse_way == 3'h2 ? tag_0_0 : _GEN_2954; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3278 = unuse_way == 3'h2 ? tag_0_1 : _GEN_2955; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3279 = unuse_way == 3'h2 ? tag_0_2 : _GEN_2956; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3280 = unuse_way == 3'h2 ? tag_0_3 : _GEN_2957; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3281 = unuse_way == 3'h2 ? tag_0_4 : _GEN_2958; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3282 = unuse_way == 3'h2 ? tag_0_5 : _GEN_2959; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3283 = unuse_way == 3'h2 ? tag_0_6 : _GEN_2960; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3284 = unuse_way == 3'h2 ? tag_0_7 : _GEN_2961; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3285 = unuse_way == 3'h2 ? tag_0_8 : _GEN_2962; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3286 = unuse_way == 3'h2 ? tag_0_9 : _GEN_2963; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3287 = unuse_way == 3'h2 ? tag_0_10 : _GEN_2964; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3288 = unuse_way == 3'h2 ? tag_0_11 : _GEN_2965; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3289 = unuse_way == 3'h2 ? tag_0_12 : _GEN_2966; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3290 = unuse_way == 3'h2 ? tag_0_13 : _GEN_2967; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3291 = unuse_way == 3'h2 ? tag_0_14 : _GEN_2968; // @[d_cache.scala 156:40 24:24]
  wire [31:0] _GEN_3292 = unuse_way == 3'h2 ? tag_0_15 : _GEN_2969; // @[d_cache.scala 156:40 24:24]
  wire  _GEN_3293 = unuse_way == 3'h2 ? dirty_0_0 : _GEN_2970; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3294 = unuse_way == 3'h2 ? dirty_0_1 : _GEN_2971; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3295 = unuse_way == 3'h2 ? dirty_0_2 : _GEN_2972; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3296 = unuse_way == 3'h2 ? dirty_0_3 : _GEN_2973; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3297 = unuse_way == 3'h2 ? dirty_0_4 : _GEN_2974; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3298 = unuse_way == 3'h2 ? dirty_0_5 : _GEN_2975; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3299 = unuse_way == 3'h2 ? dirty_0_6 : _GEN_2976; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3300 = unuse_way == 3'h2 ? dirty_0_7 : _GEN_2977; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3301 = unuse_way == 3'h2 ? dirty_0_8 : _GEN_2978; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3302 = unuse_way == 3'h2 ? dirty_0_9 : _GEN_2979; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3303 = unuse_way == 3'h2 ? dirty_0_10 : _GEN_2980; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3304 = unuse_way == 3'h2 ? dirty_0_11 : _GEN_2981; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3305 = unuse_way == 3'h2 ? dirty_0_12 : _GEN_2982; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3306 = unuse_way == 3'h2 ? dirty_0_13 : _GEN_2983; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3307 = unuse_way == 3'h2 ? dirty_0_14 : _GEN_2984; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3308 = unuse_way == 3'h2 ? dirty_0_15 : _GEN_2985; // @[d_cache.scala 156:40 34:26]
  wire  _GEN_3309 = unuse_way == 3'h2 ? valid_0_0 : _GEN_2986; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3310 = unuse_way == 3'h2 ? valid_0_1 : _GEN_2987; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3311 = unuse_way == 3'h2 ? valid_0_2 : _GEN_2988; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3312 = unuse_way == 3'h2 ? valid_0_3 : _GEN_2989; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3313 = unuse_way == 3'h2 ? valid_0_4 : _GEN_2990; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3314 = unuse_way == 3'h2 ? valid_0_5 : _GEN_2991; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3315 = unuse_way == 3'h2 ? valid_0_6 : _GEN_2992; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3316 = unuse_way == 3'h2 ? valid_0_7 : _GEN_2993; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3317 = unuse_way == 3'h2 ? valid_0_8 : _GEN_2994; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3318 = unuse_way == 3'h2 ? valid_0_9 : _GEN_2995; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3319 = unuse_way == 3'h2 ? valid_0_10 : _GEN_2996; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3320 = unuse_way == 3'h2 ? valid_0_11 : _GEN_2997; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3321 = unuse_way == 3'h2 ? valid_0_12 : _GEN_2998; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3322 = unuse_way == 3'h2 ? valid_0_13 : _GEN_2999; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3323 = unuse_way == 3'h2 ? valid_0_14 : _GEN_3000; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3324 = unuse_way == 3'h2 ? valid_0_15 : _GEN_3001; // @[d_cache.scala 156:40 29:26]
  wire  _GEN_3325 = unuse_way == 3'h2 ? dirty_1_0 : _GEN_3034; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3326 = unuse_way == 3'h2 ? dirty_1_1 : _GEN_3035; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3327 = unuse_way == 3'h2 ? dirty_1_2 : _GEN_3036; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3328 = unuse_way == 3'h2 ? dirty_1_3 : _GEN_3037; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3329 = unuse_way == 3'h2 ? dirty_1_4 : _GEN_3038; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3330 = unuse_way == 3'h2 ? dirty_1_5 : _GEN_3039; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3331 = unuse_way == 3'h2 ? dirty_1_6 : _GEN_3040; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3332 = unuse_way == 3'h2 ? dirty_1_7 : _GEN_3041; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3333 = unuse_way == 3'h2 ? dirty_1_8 : _GEN_3042; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3334 = unuse_way == 3'h2 ? dirty_1_9 : _GEN_3043; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3335 = unuse_way == 3'h2 ? dirty_1_10 : _GEN_3044; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3336 = unuse_way == 3'h2 ? dirty_1_11 : _GEN_3045; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3337 = unuse_way == 3'h2 ? dirty_1_12 : _GEN_3046; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3338 = unuse_way == 3'h2 ? dirty_1_13 : _GEN_3047; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3339 = unuse_way == 3'h2 ? dirty_1_14 : _GEN_3048; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3340 = unuse_way == 3'h2 ? dirty_1_15 : _GEN_3049; // @[d_cache.scala 156:40 35:26]
  wire  _GEN_3341 = unuse_way == 3'h2 ? dirty_2_0 : _GEN_3066; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3342 = unuse_way == 3'h2 ? dirty_2_1 : _GEN_3067; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3343 = unuse_way == 3'h2 ? dirty_2_2 : _GEN_3068; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3344 = unuse_way == 3'h2 ? dirty_2_3 : _GEN_3069; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3345 = unuse_way == 3'h2 ? dirty_2_4 : _GEN_3070; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3346 = unuse_way == 3'h2 ? dirty_2_5 : _GEN_3071; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3347 = unuse_way == 3'h2 ? dirty_2_6 : _GEN_3072; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3348 = unuse_way == 3'h2 ? dirty_2_7 : _GEN_3073; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3349 = unuse_way == 3'h2 ? dirty_2_8 : _GEN_3074; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3350 = unuse_way == 3'h2 ? dirty_2_9 : _GEN_3075; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3351 = unuse_way == 3'h2 ? dirty_2_10 : _GEN_3076; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3352 = unuse_way == 3'h2 ? dirty_2_11 : _GEN_3077; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3353 = unuse_way == 3'h2 ? dirty_2_12 : _GEN_3078; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3354 = unuse_way == 3'h2 ? dirty_2_13 : _GEN_3079; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3355 = unuse_way == 3'h2 ? dirty_2_14 : _GEN_3080; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3356 = unuse_way == 3'h2 ? dirty_2_15 : _GEN_3081; // @[d_cache.scala 156:40 36:26]
  wire  _GEN_3357 = unuse_way == 3'h2 ? dirty_3_0 : _GEN_3082; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3358 = unuse_way == 3'h2 ? dirty_3_1 : _GEN_3083; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3359 = unuse_way == 3'h2 ? dirty_3_2 : _GEN_3084; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3360 = unuse_way == 3'h2 ? dirty_3_3 : _GEN_3085; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3361 = unuse_way == 3'h2 ? dirty_3_4 : _GEN_3086; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3362 = unuse_way == 3'h2 ? dirty_3_5 : _GEN_3087; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3363 = unuse_way == 3'h2 ? dirty_3_6 : _GEN_3088; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3364 = unuse_way == 3'h2 ? dirty_3_7 : _GEN_3089; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3365 = unuse_way == 3'h2 ? dirty_3_8 : _GEN_3090; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3366 = unuse_way == 3'h2 ? dirty_3_9 : _GEN_3091; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3367 = unuse_way == 3'h2 ? dirty_3_10 : _GEN_3092; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3368 = unuse_way == 3'h2 ? dirty_3_11 : _GEN_3093; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3369 = unuse_way == 3'h2 ? dirty_3_12 : _GEN_3094; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3370 = unuse_way == 3'h2 ? dirty_3_13 : _GEN_3095; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3371 = unuse_way == 3'h2 ? dirty_3_14 : _GEN_3096; // @[d_cache.scala 156:40 37:26]
  wire  _GEN_3372 = unuse_way == 3'h2 ? dirty_3_15 : _GEN_3097; // @[d_cache.scala 156:40 37:26]
  wire [3:0] _GEN_3373 = unuse_way == 3'h1 ? 4'h1 : _GEN_3098; // @[d_cache.scala 150:34 151:23]
  wire [511:0] _GEN_3374 = unuse_way == 3'h1 ? _GEN_671 : _GEN_3261; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3375 = unuse_way == 3'h1 ? _GEN_672 : _GEN_3262; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3376 = unuse_way == 3'h1 ? _GEN_673 : _GEN_3263; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3377 = unuse_way == 3'h1 ? _GEN_674 : _GEN_3264; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3378 = unuse_way == 3'h1 ? _GEN_675 : _GEN_3265; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3379 = unuse_way == 3'h1 ? _GEN_676 : _GEN_3266; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3380 = unuse_way == 3'h1 ? _GEN_677 : _GEN_3267; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3381 = unuse_way == 3'h1 ? _GEN_678 : _GEN_3268; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3382 = unuse_way == 3'h1 ? _GEN_679 : _GEN_3269; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3383 = unuse_way == 3'h1 ? _GEN_680 : _GEN_3270; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3384 = unuse_way == 3'h1 ? _GEN_681 : _GEN_3271; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3385 = unuse_way == 3'h1 ? _GEN_682 : _GEN_3272; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3386 = unuse_way == 3'h1 ? _GEN_683 : _GEN_3273; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3387 = unuse_way == 3'h1 ? _GEN_684 : _GEN_3274; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3388 = unuse_way == 3'h1 ? _GEN_685 : _GEN_3275; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3389 = unuse_way == 3'h1 ? _GEN_686 : _GEN_3276; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3390 = unuse_way == 3'h1 ? _GEN_687 : _GEN_3277; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3391 = unuse_way == 3'h1 ? _GEN_688 : _GEN_3278; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3392 = unuse_way == 3'h1 ? _GEN_689 : _GEN_3279; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3393 = unuse_way == 3'h1 ? _GEN_690 : _GEN_3280; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3394 = unuse_way == 3'h1 ? _GEN_691 : _GEN_3281; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3395 = unuse_way == 3'h1 ? _GEN_692 : _GEN_3282; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3396 = unuse_way == 3'h1 ? _GEN_693 : _GEN_3283; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3397 = unuse_way == 3'h1 ? _GEN_694 : _GEN_3284; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3398 = unuse_way == 3'h1 ? _GEN_695 : _GEN_3285; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3399 = unuse_way == 3'h1 ? _GEN_696 : _GEN_3286; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3400 = unuse_way == 3'h1 ? _GEN_697 : _GEN_3287; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3401 = unuse_way == 3'h1 ? _GEN_698 : _GEN_3288; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3402 = unuse_way == 3'h1 ? _GEN_699 : _GEN_3289; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3403 = unuse_way == 3'h1 ? _GEN_700 : _GEN_3290; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3404 = unuse_way == 3'h1 ? _GEN_701 : _GEN_3291; // @[d_cache.scala 150:34]
  wire [31:0] _GEN_3405 = unuse_way == 3'h1 ? _GEN_702 : _GEN_3292; // @[d_cache.scala 150:34]
  wire  _GEN_3406 = unuse_way == 3'h1 ? _GEN_703 : _GEN_3309; // @[d_cache.scala 150:34]
  wire  _GEN_3407 = unuse_way == 3'h1 ? _GEN_704 : _GEN_3310; // @[d_cache.scala 150:34]
  wire  _GEN_3408 = unuse_way == 3'h1 ? _GEN_705 : _GEN_3311; // @[d_cache.scala 150:34]
  wire  _GEN_3409 = unuse_way == 3'h1 ? _GEN_706 : _GEN_3312; // @[d_cache.scala 150:34]
  wire  _GEN_3410 = unuse_way == 3'h1 ? _GEN_707 : _GEN_3313; // @[d_cache.scala 150:34]
  wire  _GEN_3411 = unuse_way == 3'h1 ? _GEN_708 : _GEN_3314; // @[d_cache.scala 150:34]
  wire  _GEN_3412 = unuse_way == 3'h1 ? _GEN_709 : _GEN_3315; // @[d_cache.scala 150:34]
  wire  _GEN_3413 = unuse_way == 3'h1 ? _GEN_710 : _GEN_3316; // @[d_cache.scala 150:34]
  wire  _GEN_3414 = unuse_way == 3'h1 ? _GEN_711 : _GEN_3317; // @[d_cache.scala 150:34]
  wire  _GEN_3415 = unuse_way == 3'h1 ? _GEN_712 : _GEN_3318; // @[d_cache.scala 150:34]
  wire  _GEN_3416 = unuse_way == 3'h1 ? _GEN_713 : _GEN_3319; // @[d_cache.scala 150:34]
  wire  _GEN_3417 = unuse_way == 3'h1 ? _GEN_714 : _GEN_3320; // @[d_cache.scala 150:34]
  wire  _GEN_3418 = unuse_way == 3'h1 ? _GEN_715 : _GEN_3321; // @[d_cache.scala 150:34]
  wire  _GEN_3419 = unuse_way == 3'h1 ? _GEN_716 : _GEN_3322; // @[d_cache.scala 150:34]
  wire  _GEN_3420 = unuse_way == 3'h1 ? _GEN_717 : _GEN_3323; // @[d_cache.scala 150:34]
  wire  _GEN_3421 = unuse_way == 3'h1 ? _GEN_718 : _GEN_3324; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3422 = unuse_way == 3'h1 ? _GEN_735 : _GEN_3147; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3423 = unuse_way == 3'h1 ? _GEN_736 : _GEN_3148; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3424 = unuse_way == 3'h1 ? _GEN_737 : _GEN_3149; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3425 = unuse_way == 3'h1 ? _GEN_738 : _GEN_3150; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3426 = unuse_way == 3'h1 ? _GEN_739 : _GEN_3151; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3427 = unuse_way == 3'h1 ? _GEN_740 : _GEN_3152; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3428 = unuse_way == 3'h1 ? _GEN_741 : _GEN_3153; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3429 = unuse_way == 3'h1 ? _GEN_742 : _GEN_3154; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3430 = unuse_way == 3'h1 ? _GEN_743 : _GEN_3155; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3431 = unuse_way == 3'h1 ? _GEN_744 : _GEN_3156; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3432 = unuse_way == 3'h1 ? _GEN_745 : _GEN_3157; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3433 = unuse_way == 3'h1 ? _GEN_746 : _GEN_3158; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3434 = unuse_way == 3'h1 ? _GEN_747 : _GEN_3159; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3435 = unuse_way == 3'h1 ? _GEN_748 : _GEN_3160; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3436 = unuse_way == 3'h1 ? _GEN_749 : _GEN_3161; // @[d_cache.scala 150:34]
  wire [7:0] _GEN_3437 = unuse_way == 3'h1 ? _GEN_750 : _GEN_3162; // @[d_cache.scala 150:34]
  wire [511:0] _GEN_3438 = unuse_way == 3'h1 ? ram_1_0 : _GEN_3099; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3439 = unuse_way == 3'h1 ? ram_1_1 : _GEN_3100; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3440 = unuse_way == 3'h1 ? ram_1_2 : _GEN_3101; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3441 = unuse_way == 3'h1 ? ram_1_3 : _GEN_3102; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3442 = unuse_way == 3'h1 ? ram_1_4 : _GEN_3103; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3443 = unuse_way == 3'h1 ? ram_1_5 : _GEN_3104; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3444 = unuse_way == 3'h1 ? ram_1_6 : _GEN_3105; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3445 = unuse_way == 3'h1 ? ram_1_7 : _GEN_3106; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3446 = unuse_way == 3'h1 ? ram_1_8 : _GEN_3107; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3447 = unuse_way == 3'h1 ? ram_1_9 : _GEN_3108; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3448 = unuse_way == 3'h1 ? ram_1_10 : _GEN_3109; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3449 = unuse_way == 3'h1 ? ram_1_11 : _GEN_3110; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3450 = unuse_way == 3'h1 ? ram_1_12 : _GEN_3111; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3451 = unuse_way == 3'h1 ? ram_1_13 : _GEN_3112; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3452 = unuse_way == 3'h1 ? ram_1_14 : _GEN_3113; // @[d_cache.scala 150:34 20:24]
  wire [511:0] _GEN_3453 = unuse_way == 3'h1 ? ram_1_15 : _GEN_3114; // @[d_cache.scala 150:34 20:24]
  wire [31:0] _GEN_3454 = unuse_way == 3'h1 ? tag_1_0 : _GEN_3115; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3455 = unuse_way == 3'h1 ? tag_1_1 : _GEN_3116; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3456 = unuse_way == 3'h1 ? tag_1_2 : _GEN_3117; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3457 = unuse_way == 3'h1 ? tag_1_3 : _GEN_3118; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3458 = unuse_way == 3'h1 ? tag_1_4 : _GEN_3119; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3459 = unuse_way == 3'h1 ? tag_1_5 : _GEN_3120; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3460 = unuse_way == 3'h1 ? tag_1_6 : _GEN_3121; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3461 = unuse_way == 3'h1 ? tag_1_7 : _GEN_3122; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3462 = unuse_way == 3'h1 ? tag_1_8 : _GEN_3123; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3463 = unuse_way == 3'h1 ? tag_1_9 : _GEN_3124; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3464 = unuse_way == 3'h1 ? tag_1_10 : _GEN_3125; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3465 = unuse_way == 3'h1 ? tag_1_11 : _GEN_3126; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3466 = unuse_way == 3'h1 ? tag_1_12 : _GEN_3127; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3467 = unuse_way == 3'h1 ? tag_1_13 : _GEN_3128; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3468 = unuse_way == 3'h1 ? tag_1_14 : _GEN_3129; // @[d_cache.scala 150:34 25:24]
  wire [31:0] _GEN_3469 = unuse_way == 3'h1 ? tag_1_15 : _GEN_3130; // @[d_cache.scala 150:34 25:24]
  wire  _GEN_3470 = unuse_way == 3'h1 ? valid_1_0 : _GEN_3131; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3471 = unuse_way == 3'h1 ? valid_1_1 : _GEN_3132; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3472 = unuse_way == 3'h1 ? valid_1_2 : _GEN_3133; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3473 = unuse_way == 3'h1 ? valid_1_3 : _GEN_3134; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3474 = unuse_way == 3'h1 ? valid_1_4 : _GEN_3135; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3475 = unuse_way == 3'h1 ? valid_1_5 : _GEN_3136; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3476 = unuse_way == 3'h1 ? valid_1_6 : _GEN_3137; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3477 = unuse_way == 3'h1 ? valid_1_7 : _GEN_3138; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3478 = unuse_way == 3'h1 ? valid_1_8 : _GEN_3139; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3479 = unuse_way == 3'h1 ? valid_1_9 : _GEN_3140; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3480 = unuse_way == 3'h1 ? valid_1_10 : _GEN_3141; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3481 = unuse_way == 3'h1 ? valid_1_11 : _GEN_3142; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3482 = unuse_way == 3'h1 ? valid_1_12 : _GEN_3143; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3483 = unuse_way == 3'h1 ? valid_1_13 : _GEN_3144; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3484 = unuse_way == 3'h1 ? valid_1_14 : _GEN_3145; // @[d_cache.scala 150:34 30:26]
  wire  _GEN_3485 = unuse_way == 3'h1 ? valid_1_15 : _GEN_3146; // @[d_cache.scala 150:34 30:26]
  wire [511:0] _GEN_3486 = unuse_way == 3'h1 ? ram_2_0 : _GEN_3163; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3487 = unuse_way == 3'h1 ? ram_2_1 : _GEN_3164; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3488 = unuse_way == 3'h1 ? ram_2_2 : _GEN_3165; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3489 = unuse_way == 3'h1 ? ram_2_3 : _GEN_3166; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3490 = unuse_way == 3'h1 ? ram_2_4 : _GEN_3167; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3491 = unuse_way == 3'h1 ? ram_2_5 : _GEN_3168; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3492 = unuse_way == 3'h1 ? ram_2_6 : _GEN_3169; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3493 = unuse_way == 3'h1 ? ram_2_7 : _GEN_3170; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3494 = unuse_way == 3'h1 ? ram_2_8 : _GEN_3171; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3495 = unuse_way == 3'h1 ? ram_2_9 : _GEN_3172; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3496 = unuse_way == 3'h1 ? ram_2_10 : _GEN_3173; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3497 = unuse_way == 3'h1 ? ram_2_11 : _GEN_3174; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3498 = unuse_way == 3'h1 ? ram_2_12 : _GEN_3175; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3499 = unuse_way == 3'h1 ? ram_2_13 : _GEN_3176; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3500 = unuse_way == 3'h1 ? ram_2_14 : _GEN_3177; // @[d_cache.scala 150:34 21:24]
  wire [511:0] _GEN_3501 = unuse_way == 3'h1 ? ram_2_15 : _GEN_3178; // @[d_cache.scala 150:34 21:24]
  wire [31:0] _GEN_3502 = unuse_way == 3'h1 ? tag_2_0 : _GEN_3179; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3503 = unuse_way == 3'h1 ? tag_2_1 : _GEN_3180; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3504 = unuse_way == 3'h1 ? tag_2_2 : _GEN_3181; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3505 = unuse_way == 3'h1 ? tag_2_3 : _GEN_3182; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3506 = unuse_way == 3'h1 ? tag_2_4 : _GEN_3183; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3507 = unuse_way == 3'h1 ? tag_2_5 : _GEN_3184; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3508 = unuse_way == 3'h1 ? tag_2_6 : _GEN_3185; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3509 = unuse_way == 3'h1 ? tag_2_7 : _GEN_3186; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3510 = unuse_way == 3'h1 ? tag_2_8 : _GEN_3187; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3511 = unuse_way == 3'h1 ? tag_2_9 : _GEN_3188; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3512 = unuse_way == 3'h1 ? tag_2_10 : _GEN_3189; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3513 = unuse_way == 3'h1 ? tag_2_11 : _GEN_3190; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3514 = unuse_way == 3'h1 ? tag_2_12 : _GEN_3191; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3515 = unuse_way == 3'h1 ? tag_2_13 : _GEN_3192; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3516 = unuse_way == 3'h1 ? tag_2_14 : _GEN_3193; // @[d_cache.scala 150:34 26:24]
  wire [31:0] _GEN_3517 = unuse_way == 3'h1 ? tag_2_15 : _GEN_3194; // @[d_cache.scala 150:34 26:24]
  wire  _GEN_3518 = unuse_way == 3'h1 ? valid_2_0 : _GEN_3195; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3519 = unuse_way == 3'h1 ? valid_2_1 : _GEN_3196; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3520 = unuse_way == 3'h1 ? valid_2_2 : _GEN_3197; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3521 = unuse_way == 3'h1 ? valid_2_3 : _GEN_3198; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3522 = unuse_way == 3'h1 ? valid_2_4 : _GEN_3199; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3523 = unuse_way == 3'h1 ? valid_2_5 : _GEN_3200; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3524 = unuse_way == 3'h1 ? valid_2_6 : _GEN_3201; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3525 = unuse_way == 3'h1 ? valid_2_7 : _GEN_3202; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3526 = unuse_way == 3'h1 ? valid_2_8 : _GEN_3203; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3527 = unuse_way == 3'h1 ? valid_2_9 : _GEN_3204; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3528 = unuse_way == 3'h1 ? valid_2_10 : _GEN_3205; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3529 = unuse_way == 3'h1 ? valid_2_11 : _GEN_3206; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3530 = unuse_way == 3'h1 ? valid_2_12 : _GEN_3207; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3531 = unuse_way == 3'h1 ? valid_2_13 : _GEN_3208; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3532 = unuse_way == 3'h1 ? valid_2_14 : _GEN_3209; // @[d_cache.scala 150:34 31:26]
  wire  _GEN_3533 = unuse_way == 3'h1 ? valid_2_15 : _GEN_3210; // @[d_cache.scala 150:34 31:26]
  wire [511:0] _GEN_3534 = unuse_way == 3'h1 ? ram_3_0 : _GEN_3211; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3535 = unuse_way == 3'h1 ? ram_3_1 : _GEN_3212; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3536 = unuse_way == 3'h1 ? ram_3_2 : _GEN_3213; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3537 = unuse_way == 3'h1 ? ram_3_3 : _GEN_3214; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3538 = unuse_way == 3'h1 ? ram_3_4 : _GEN_3215; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3539 = unuse_way == 3'h1 ? ram_3_5 : _GEN_3216; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3540 = unuse_way == 3'h1 ? ram_3_6 : _GEN_3217; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3541 = unuse_way == 3'h1 ? ram_3_7 : _GEN_3218; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3542 = unuse_way == 3'h1 ? ram_3_8 : _GEN_3219; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3543 = unuse_way == 3'h1 ? ram_3_9 : _GEN_3220; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3544 = unuse_way == 3'h1 ? ram_3_10 : _GEN_3221; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3545 = unuse_way == 3'h1 ? ram_3_11 : _GEN_3222; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3546 = unuse_way == 3'h1 ? ram_3_12 : _GEN_3223; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3547 = unuse_way == 3'h1 ? ram_3_13 : _GEN_3224; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3548 = unuse_way == 3'h1 ? ram_3_14 : _GEN_3225; // @[d_cache.scala 150:34 22:24]
  wire [511:0] _GEN_3549 = unuse_way == 3'h1 ? ram_3_15 : _GEN_3226; // @[d_cache.scala 150:34 22:24]
  wire [31:0] _GEN_3550 = unuse_way == 3'h1 ? tag_3_0 : _GEN_3227; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3551 = unuse_way == 3'h1 ? tag_3_1 : _GEN_3228; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3552 = unuse_way == 3'h1 ? tag_3_2 : _GEN_3229; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3553 = unuse_way == 3'h1 ? tag_3_3 : _GEN_3230; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3554 = unuse_way == 3'h1 ? tag_3_4 : _GEN_3231; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3555 = unuse_way == 3'h1 ? tag_3_5 : _GEN_3232; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3556 = unuse_way == 3'h1 ? tag_3_6 : _GEN_3233; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3557 = unuse_way == 3'h1 ? tag_3_7 : _GEN_3234; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3558 = unuse_way == 3'h1 ? tag_3_8 : _GEN_3235; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3559 = unuse_way == 3'h1 ? tag_3_9 : _GEN_3236; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3560 = unuse_way == 3'h1 ? tag_3_10 : _GEN_3237; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3561 = unuse_way == 3'h1 ? tag_3_11 : _GEN_3238; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3562 = unuse_way == 3'h1 ? tag_3_12 : _GEN_3239; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3563 = unuse_way == 3'h1 ? tag_3_13 : _GEN_3240; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3564 = unuse_way == 3'h1 ? tag_3_14 : _GEN_3241; // @[d_cache.scala 150:34 27:24]
  wire [31:0] _GEN_3565 = unuse_way == 3'h1 ? tag_3_15 : _GEN_3242; // @[d_cache.scala 150:34 27:24]
  wire  _GEN_3566 = unuse_way == 3'h1 ? valid_3_0 : _GEN_3243; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3567 = unuse_way == 3'h1 ? valid_3_1 : _GEN_3244; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3568 = unuse_way == 3'h1 ? valid_3_2 : _GEN_3245; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3569 = unuse_way == 3'h1 ? valid_3_3 : _GEN_3246; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3570 = unuse_way == 3'h1 ? valid_3_4 : _GEN_3247; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3571 = unuse_way == 3'h1 ? valid_3_5 : _GEN_3248; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3572 = unuse_way == 3'h1 ? valid_3_6 : _GEN_3249; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3573 = unuse_way == 3'h1 ? valid_3_7 : _GEN_3250; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3574 = unuse_way == 3'h1 ? valid_3_8 : _GEN_3251; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3575 = unuse_way == 3'h1 ? valid_3_9 : _GEN_3252; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3576 = unuse_way == 3'h1 ? valid_3_10 : _GEN_3253; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3577 = unuse_way == 3'h1 ? valid_3_11 : _GEN_3254; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3578 = unuse_way == 3'h1 ? valid_3_12 : _GEN_3255; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3579 = unuse_way == 3'h1 ? valid_3_13 : _GEN_3256; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3580 = unuse_way == 3'h1 ? valid_3_14 : _GEN_3257; // @[d_cache.scala 150:34 32:26]
  wire  _GEN_3581 = unuse_way == 3'h1 ? valid_3_15 : _GEN_3258; // @[d_cache.scala 150:34 32:26]
  wire [511:0] _GEN_3582 = unuse_way == 3'h1 ? write_back_data : _GEN_3259; // @[d_cache.scala 150:34 44:34]
  wire [41:0] _GEN_3583 = unuse_way == 3'h1 ? {{10'd0}, write_back_addr} : _GEN_3260; // @[d_cache.scala 150:34 45:34]
  wire  _GEN_3584 = unuse_way == 3'h1 ? dirty_0_0 : _GEN_3293; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3585 = unuse_way == 3'h1 ? dirty_0_1 : _GEN_3294; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3586 = unuse_way == 3'h1 ? dirty_0_2 : _GEN_3295; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3587 = unuse_way == 3'h1 ? dirty_0_3 : _GEN_3296; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3588 = unuse_way == 3'h1 ? dirty_0_4 : _GEN_3297; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3589 = unuse_way == 3'h1 ? dirty_0_5 : _GEN_3298; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3590 = unuse_way == 3'h1 ? dirty_0_6 : _GEN_3299; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3591 = unuse_way == 3'h1 ? dirty_0_7 : _GEN_3300; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3592 = unuse_way == 3'h1 ? dirty_0_8 : _GEN_3301; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3593 = unuse_way == 3'h1 ? dirty_0_9 : _GEN_3302; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3594 = unuse_way == 3'h1 ? dirty_0_10 : _GEN_3303; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3595 = unuse_way == 3'h1 ? dirty_0_11 : _GEN_3304; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3596 = unuse_way == 3'h1 ? dirty_0_12 : _GEN_3305; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3597 = unuse_way == 3'h1 ? dirty_0_13 : _GEN_3306; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3598 = unuse_way == 3'h1 ? dirty_0_14 : _GEN_3307; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3599 = unuse_way == 3'h1 ? dirty_0_15 : _GEN_3308; // @[d_cache.scala 150:34 34:26]
  wire  _GEN_3600 = unuse_way == 3'h1 ? dirty_1_0 : _GEN_3325; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3601 = unuse_way == 3'h1 ? dirty_1_1 : _GEN_3326; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3602 = unuse_way == 3'h1 ? dirty_1_2 : _GEN_3327; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3603 = unuse_way == 3'h1 ? dirty_1_3 : _GEN_3328; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3604 = unuse_way == 3'h1 ? dirty_1_4 : _GEN_3329; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3605 = unuse_way == 3'h1 ? dirty_1_5 : _GEN_3330; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3606 = unuse_way == 3'h1 ? dirty_1_6 : _GEN_3331; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3607 = unuse_way == 3'h1 ? dirty_1_7 : _GEN_3332; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3608 = unuse_way == 3'h1 ? dirty_1_8 : _GEN_3333; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3609 = unuse_way == 3'h1 ? dirty_1_9 : _GEN_3334; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3610 = unuse_way == 3'h1 ? dirty_1_10 : _GEN_3335; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3611 = unuse_way == 3'h1 ? dirty_1_11 : _GEN_3336; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3612 = unuse_way == 3'h1 ? dirty_1_12 : _GEN_3337; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3613 = unuse_way == 3'h1 ? dirty_1_13 : _GEN_3338; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3614 = unuse_way == 3'h1 ? dirty_1_14 : _GEN_3339; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3615 = unuse_way == 3'h1 ? dirty_1_15 : _GEN_3340; // @[d_cache.scala 150:34 35:26]
  wire  _GEN_3616 = unuse_way == 3'h1 ? dirty_2_0 : _GEN_3341; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3617 = unuse_way == 3'h1 ? dirty_2_1 : _GEN_3342; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3618 = unuse_way == 3'h1 ? dirty_2_2 : _GEN_3343; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3619 = unuse_way == 3'h1 ? dirty_2_3 : _GEN_3344; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3620 = unuse_way == 3'h1 ? dirty_2_4 : _GEN_3345; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3621 = unuse_way == 3'h1 ? dirty_2_5 : _GEN_3346; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3622 = unuse_way == 3'h1 ? dirty_2_6 : _GEN_3347; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3623 = unuse_way == 3'h1 ? dirty_2_7 : _GEN_3348; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3624 = unuse_way == 3'h1 ? dirty_2_8 : _GEN_3349; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3625 = unuse_way == 3'h1 ? dirty_2_9 : _GEN_3350; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3626 = unuse_way == 3'h1 ? dirty_2_10 : _GEN_3351; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3627 = unuse_way == 3'h1 ? dirty_2_11 : _GEN_3352; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3628 = unuse_way == 3'h1 ? dirty_2_12 : _GEN_3353; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3629 = unuse_way == 3'h1 ? dirty_2_13 : _GEN_3354; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3630 = unuse_way == 3'h1 ? dirty_2_14 : _GEN_3355; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3631 = unuse_way == 3'h1 ? dirty_2_15 : _GEN_3356; // @[d_cache.scala 150:34 36:26]
  wire  _GEN_3632 = unuse_way == 3'h1 ? dirty_3_0 : _GEN_3357; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3633 = unuse_way == 3'h1 ? dirty_3_1 : _GEN_3358; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3634 = unuse_way == 3'h1 ? dirty_3_2 : _GEN_3359; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3635 = unuse_way == 3'h1 ? dirty_3_3 : _GEN_3360; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3636 = unuse_way == 3'h1 ? dirty_3_4 : _GEN_3361; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3637 = unuse_way == 3'h1 ? dirty_3_5 : _GEN_3362; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3638 = unuse_way == 3'h1 ? dirty_3_6 : _GEN_3363; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3639 = unuse_way == 3'h1 ? dirty_3_7 : _GEN_3364; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3640 = unuse_way == 3'h1 ? dirty_3_8 : _GEN_3365; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3641 = unuse_way == 3'h1 ? dirty_3_9 : _GEN_3366; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3642 = unuse_way == 3'h1 ? dirty_3_10 : _GEN_3367; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3643 = unuse_way == 3'h1 ? dirty_3_11 : _GEN_3368; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3644 = unuse_way == 3'h1 ? dirty_3_12 : _GEN_3369; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3645 = unuse_way == 3'h1 ? dirty_3_13 : _GEN_3370; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3646 = unuse_way == 3'h1 ? dirty_3_14 : _GEN_3371; // @[d_cache.scala 150:34 37:26]
  wire  _GEN_3647 = unuse_way == 3'h1 ? dirty_3_15 : _GEN_3372; // @[d_cache.scala 150:34 37:26]
  wire [511:0] _write_back_data_T = {{64'd0}, write_back_data[511:64]}; // @[d_cache.scala 248:52]
  wire [511:0] _GEN_3648 = io_from_axi_wready ? _write_back_data_T : write_back_data; // @[d_cache.scala 247:37 248:33 44:34]
  wire [3:0] _GEN_3649 = io_from_axi_bvalid ? 4'h1 : state; // @[d_cache.scala 250:37 251:23 82:24]
  wire [3:0] _GEN_3650 = io_from_axi_rvalid ? 4'h0 : state; // @[d_cache.scala 255:37 256:23 82:24]
  wire [3:0] _GEN_3651 = 4'h8 == state ? _GEN_670 : state; // @[d_cache.scala 87:18 82:24]
  wire [3:0] _GEN_3652 = 4'h7 == state ? _GEN_3650 : _GEN_3651; // @[d_cache.scala 87:18]
  wire [511:0] _GEN_3653 = 4'h6 == state ? _GEN_3648 : write_back_data; // @[d_cache.scala 87:18 44:34]
  wire [3:0] _GEN_3654 = 4'h6 == state ? _GEN_3649 : _GEN_3652; // @[d_cache.scala 87:18]
  wire [3:0] _GEN_3655 = 4'h5 == state ? _GEN_3373 : _GEN_3654; // @[d_cache.scala 87:18]
  wire [511:0] _GEN_3656 = 4'h5 == state ? _GEN_3374 : ram_0_0; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3657 = 4'h5 == state ? _GEN_3375 : ram_0_1; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3658 = 4'h5 == state ? _GEN_3376 : ram_0_2; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3659 = 4'h5 == state ? _GEN_3377 : ram_0_3; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3660 = 4'h5 == state ? _GEN_3378 : ram_0_4; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3661 = 4'h5 == state ? _GEN_3379 : ram_0_5; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3662 = 4'h5 == state ? _GEN_3380 : ram_0_6; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3663 = 4'h5 == state ? _GEN_3381 : ram_0_7; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3664 = 4'h5 == state ? _GEN_3382 : ram_0_8; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3665 = 4'h5 == state ? _GEN_3383 : ram_0_9; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3666 = 4'h5 == state ? _GEN_3384 : ram_0_10; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3667 = 4'h5 == state ? _GEN_3385 : ram_0_11; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3668 = 4'h5 == state ? _GEN_3386 : ram_0_12; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3669 = 4'h5 == state ? _GEN_3387 : ram_0_13; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3670 = 4'h5 == state ? _GEN_3388 : ram_0_14; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3671 = 4'h5 == state ? _GEN_3389 : ram_0_15; // @[d_cache.scala 87:18 19:24]
  wire [31:0] _GEN_3672 = 4'h5 == state ? _GEN_3390 : tag_0_0; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3673 = 4'h5 == state ? _GEN_3391 : tag_0_1; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3674 = 4'h5 == state ? _GEN_3392 : tag_0_2; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3675 = 4'h5 == state ? _GEN_3393 : tag_0_3; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3676 = 4'h5 == state ? _GEN_3394 : tag_0_4; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3677 = 4'h5 == state ? _GEN_3395 : tag_0_5; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3678 = 4'h5 == state ? _GEN_3396 : tag_0_6; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3679 = 4'h5 == state ? _GEN_3397 : tag_0_7; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3680 = 4'h5 == state ? _GEN_3398 : tag_0_8; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3681 = 4'h5 == state ? _GEN_3399 : tag_0_9; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3682 = 4'h5 == state ? _GEN_3400 : tag_0_10; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3683 = 4'h5 == state ? _GEN_3401 : tag_0_11; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3684 = 4'h5 == state ? _GEN_3402 : tag_0_12; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3685 = 4'h5 == state ? _GEN_3403 : tag_0_13; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3686 = 4'h5 == state ? _GEN_3404 : tag_0_14; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3687 = 4'h5 == state ? _GEN_3405 : tag_0_15; // @[d_cache.scala 87:18 24:24]
  wire  _GEN_3688 = 4'h5 == state ? _GEN_3406 : valid_0_0; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3689 = 4'h5 == state ? _GEN_3407 : valid_0_1; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3690 = 4'h5 == state ? _GEN_3408 : valid_0_2; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3691 = 4'h5 == state ? _GEN_3409 : valid_0_3; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3692 = 4'h5 == state ? _GEN_3410 : valid_0_4; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3693 = 4'h5 == state ? _GEN_3411 : valid_0_5; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3694 = 4'h5 == state ? _GEN_3412 : valid_0_6; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3695 = 4'h5 == state ? _GEN_3413 : valid_0_7; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3696 = 4'h5 == state ? _GEN_3414 : valid_0_8; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3697 = 4'h5 == state ? _GEN_3415 : valid_0_9; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3698 = 4'h5 == state ? _GEN_3416 : valid_0_10; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3699 = 4'h5 == state ? _GEN_3417 : valid_0_11; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3700 = 4'h5 == state ? _GEN_3418 : valid_0_12; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3701 = 4'h5 == state ? _GEN_3419 : valid_0_13; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3702 = 4'h5 == state ? _GEN_3420 : valid_0_14; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3703 = 4'h5 == state ? _GEN_3421 : valid_0_15; // @[d_cache.scala 87:18 29:26]
  wire [7:0] _GEN_3704 = 4'h5 == state ? _GEN_3422 : quene_0; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3705 = 4'h5 == state ? _GEN_3423 : quene_1; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3706 = 4'h5 == state ? _GEN_3424 : quene_2; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3707 = 4'h5 == state ? _GEN_3425 : quene_3; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3708 = 4'h5 == state ? _GEN_3426 : quene_4; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3709 = 4'h5 == state ? _GEN_3427 : quene_5; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3710 = 4'h5 == state ? _GEN_3428 : quene_6; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3711 = 4'h5 == state ? _GEN_3429 : quene_7; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3712 = 4'h5 == state ? _GEN_3430 : quene_8; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3713 = 4'h5 == state ? _GEN_3431 : quene_9; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3714 = 4'h5 == state ? _GEN_3432 : quene_10; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3715 = 4'h5 == state ? _GEN_3433 : quene_11; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3716 = 4'h5 == state ? _GEN_3434 : quene_12; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3717 = 4'h5 == state ? _GEN_3435 : quene_13; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3718 = 4'h5 == state ? _GEN_3436 : quene_14; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3719 = 4'h5 == state ? _GEN_3437 : quene_15; // @[d_cache.scala 87:18 52:24]
  wire [511:0] _GEN_3720 = 4'h5 == state ? _GEN_3438 : ram_1_0; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3721 = 4'h5 == state ? _GEN_3439 : ram_1_1; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3722 = 4'h5 == state ? _GEN_3440 : ram_1_2; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3723 = 4'h5 == state ? _GEN_3441 : ram_1_3; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3724 = 4'h5 == state ? _GEN_3442 : ram_1_4; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3725 = 4'h5 == state ? _GEN_3443 : ram_1_5; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3726 = 4'h5 == state ? _GEN_3444 : ram_1_6; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3727 = 4'h5 == state ? _GEN_3445 : ram_1_7; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3728 = 4'h5 == state ? _GEN_3446 : ram_1_8; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3729 = 4'h5 == state ? _GEN_3447 : ram_1_9; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3730 = 4'h5 == state ? _GEN_3448 : ram_1_10; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3731 = 4'h5 == state ? _GEN_3449 : ram_1_11; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3732 = 4'h5 == state ? _GEN_3450 : ram_1_12; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3733 = 4'h5 == state ? _GEN_3451 : ram_1_13; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3734 = 4'h5 == state ? _GEN_3452 : ram_1_14; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3735 = 4'h5 == state ? _GEN_3453 : ram_1_15; // @[d_cache.scala 87:18 20:24]
  wire [31:0] _GEN_3736 = 4'h5 == state ? _GEN_3454 : tag_1_0; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3737 = 4'h5 == state ? _GEN_3455 : tag_1_1; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3738 = 4'h5 == state ? _GEN_3456 : tag_1_2; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3739 = 4'h5 == state ? _GEN_3457 : tag_1_3; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3740 = 4'h5 == state ? _GEN_3458 : tag_1_4; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3741 = 4'h5 == state ? _GEN_3459 : tag_1_5; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3742 = 4'h5 == state ? _GEN_3460 : tag_1_6; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3743 = 4'h5 == state ? _GEN_3461 : tag_1_7; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3744 = 4'h5 == state ? _GEN_3462 : tag_1_8; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3745 = 4'h5 == state ? _GEN_3463 : tag_1_9; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3746 = 4'h5 == state ? _GEN_3464 : tag_1_10; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3747 = 4'h5 == state ? _GEN_3465 : tag_1_11; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3748 = 4'h5 == state ? _GEN_3466 : tag_1_12; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3749 = 4'h5 == state ? _GEN_3467 : tag_1_13; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3750 = 4'h5 == state ? _GEN_3468 : tag_1_14; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_3751 = 4'h5 == state ? _GEN_3469 : tag_1_15; // @[d_cache.scala 87:18 25:24]
  wire  _GEN_3752 = 4'h5 == state ? _GEN_3470 : valid_1_0; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3753 = 4'h5 == state ? _GEN_3471 : valid_1_1; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3754 = 4'h5 == state ? _GEN_3472 : valid_1_2; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3755 = 4'h5 == state ? _GEN_3473 : valid_1_3; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3756 = 4'h5 == state ? _GEN_3474 : valid_1_4; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3757 = 4'h5 == state ? _GEN_3475 : valid_1_5; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3758 = 4'h5 == state ? _GEN_3476 : valid_1_6; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3759 = 4'h5 == state ? _GEN_3477 : valid_1_7; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3760 = 4'h5 == state ? _GEN_3478 : valid_1_8; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3761 = 4'h5 == state ? _GEN_3479 : valid_1_9; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3762 = 4'h5 == state ? _GEN_3480 : valid_1_10; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3763 = 4'h5 == state ? _GEN_3481 : valid_1_11; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3764 = 4'h5 == state ? _GEN_3482 : valid_1_12; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3765 = 4'h5 == state ? _GEN_3483 : valid_1_13; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3766 = 4'h5 == state ? _GEN_3484 : valid_1_14; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_3767 = 4'h5 == state ? _GEN_3485 : valid_1_15; // @[d_cache.scala 87:18 30:26]
  wire [511:0] _GEN_3768 = 4'h5 == state ? _GEN_3486 : ram_2_0; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3769 = 4'h5 == state ? _GEN_3487 : ram_2_1; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3770 = 4'h5 == state ? _GEN_3488 : ram_2_2; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3771 = 4'h5 == state ? _GEN_3489 : ram_2_3; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3772 = 4'h5 == state ? _GEN_3490 : ram_2_4; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3773 = 4'h5 == state ? _GEN_3491 : ram_2_5; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3774 = 4'h5 == state ? _GEN_3492 : ram_2_6; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3775 = 4'h5 == state ? _GEN_3493 : ram_2_7; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3776 = 4'h5 == state ? _GEN_3494 : ram_2_8; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3777 = 4'h5 == state ? _GEN_3495 : ram_2_9; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3778 = 4'h5 == state ? _GEN_3496 : ram_2_10; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3779 = 4'h5 == state ? _GEN_3497 : ram_2_11; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3780 = 4'h5 == state ? _GEN_3498 : ram_2_12; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3781 = 4'h5 == state ? _GEN_3499 : ram_2_13; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3782 = 4'h5 == state ? _GEN_3500 : ram_2_14; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_3783 = 4'h5 == state ? _GEN_3501 : ram_2_15; // @[d_cache.scala 87:18 21:24]
  wire [31:0] _GEN_3784 = 4'h5 == state ? _GEN_3502 : tag_2_0; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3785 = 4'h5 == state ? _GEN_3503 : tag_2_1; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3786 = 4'h5 == state ? _GEN_3504 : tag_2_2; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3787 = 4'h5 == state ? _GEN_3505 : tag_2_3; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3788 = 4'h5 == state ? _GEN_3506 : tag_2_4; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3789 = 4'h5 == state ? _GEN_3507 : tag_2_5; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3790 = 4'h5 == state ? _GEN_3508 : tag_2_6; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3791 = 4'h5 == state ? _GEN_3509 : tag_2_7; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3792 = 4'h5 == state ? _GEN_3510 : tag_2_8; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3793 = 4'h5 == state ? _GEN_3511 : tag_2_9; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3794 = 4'h5 == state ? _GEN_3512 : tag_2_10; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3795 = 4'h5 == state ? _GEN_3513 : tag_2_11; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3796 = 4'h5 == state ? _GEN_3514 : tag_2_12; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3797 = 4'h5 == state ? _GEN_3515 : tag_2_13; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3798 = 4'h5 == state ? _GEN_3516 : tag_2_14; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_3799 = 4'h5 == state ? _GEN_3517 : tag_2_15; // @[d_cache.scala 87:18 26:24]
  wire  _GEN_3800 = 4'h5 == state ? _GEN_3518 : valid_2_0; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3801 = 4'h5 == state ? _GEN_3519 : valid_2_1; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3802 = 4'h5 == state ? _GEN_3520 : valid_2_2; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3803 = 4'h5 == state ? _GEN_3521 : valid_2_3; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3804 = 4'h5 == state ? _GEN_3522 : valid_2_4; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3805 = 4'h5 == state ? _GEN_3523 : valid_2_5; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3806 = 4'h5 == state ? _GEN_3524 : valid_2_6; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3807 = 4'h5 == state ? _GEN_3525 : valid_2_7; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3808 = 4'h5 == state ? _GEN_3526 : valid_2_8; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3809 = 4'h5 == state ? _GEN_3527 : valid_2_9; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3810 = 4'h5 == state ? _GEN_3528 : valid_2_10; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3811 = 4'h5 == state ? _GEN_3529 : valid_2_11; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3812 = 4'h5 == state ? _GEN_3530 : valid_2_12; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3813 = 4'h5 == state ? _GEN_3531 : valid_2_13; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3814 = 4'h5 == state ? _GEN_3532 : valid_2_14; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_3815 = 4'h5 == state ? _GEN_3533 : valid_2_15; // @[d_cache.scala 87:18 31:26]
  wire [511:0] _GEN_3816 = 4'h5 == state ? _GEN_3534 : ram_3_0; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3817 = 4'h5 == state ? _GEN_3535 : ram_3_1; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3818 = 4'h5 == state ? _GEN_3536 : ram_3_2; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3819 = 4'h5 == state ? _GEN_3537 : ram_3_3; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3820 = 4'h5 == state ? _GEN_3538 : ram_3_4; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3821 = 4'h5 == state ? _GEN_3539 : ram_3_5; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3822 = 4'h5 == state ? _GEN_3540 : ram_3_6; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3823 = 4'h5 == state ? _GEN_3541 : ram_3_7; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3824 = 4'h5 == state ? _GEN_3542 : ram_3_8; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3825 = 4'h5 == state ? _GEN_3543 : ram_3_9; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3826 = 4'h5 == state ? _GEN_3544 : ram_3_10; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3827 = 4'h5 == state ? _GEN_3545 : ram_3_11; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3828 = 4'h5 == state ? _GEN_3546 : ram_3_12; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3829 = 4'h5 == state ? _GEN_3547 : ram_3_13; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3830 = 4'h5 == state ? _GEN_3548 : ram_3_14; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_3831 = 4'h5 == state ? _GEN_3549 : ram_3_15; // @[d_cache.scala 87:18 22:24]
  wire [31:0] _GEN_3832 = 4'h5 == state ? _GEN_3550 : tag_3_0; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3833 = 4'h5 == state ? _GEN_3551 : tag_3_1; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3834 = 4'h5 == state ? _GEN_3552 : tag_3_2; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3835 = 4'h5 == state ? _GEN_3553 : tag_3_3; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3836 = 4'h5 == state ? _GEN_3554 : tag_3_4; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3837 = 4'h5 == state ? _GEN_3555 : tag_3_5; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3838 = 4'h5 == state ? _GEN_3556 : tag_3_6; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3839 = 4'h5 == state ? _GEN_3557 : tag_3_7; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3840 = 4'h5 == state ? _GEN_3558 : tag_3_8; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3841 = 4'h5 == state ? _GEN_3559 : tag_3_9; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3842 = 4'h5 == state ? _GEN_3560 : tag_3_10; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3843 = 4'h5 == state ? _GEN_3561 : tag_3_11; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3844 = 4'h5 == state ? _GEN_3562 : tag_3_12; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3845 = 4'h5 == state ? _GEN_3563 : tag_3_13; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3846 = 4'h5 == state ? _GEN_3564 : tag_3_14; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_3847 = 4'h5 == state ? _GEN_3565 : tag_3_15; // @[d_cache.scala 87:18 27:24]
  wire  _GEN_3848 = 4'h5 == state ? _GEN_3566 : valid_3_0; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3849 = 4'h5 == state ? _GEN_3567 : valid_3_1; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3850 = 4'h5 == state ? _GEN_3568 : valid_3_2; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3851 = 4'h5 == state ? _GEN_3569 : valid_3_3; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3852 = 4'h5 == state ? _GEN_3570 : valid_3_4; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3853 = 4'h5 == state ? _GEN_3571 : valid_3_5; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3854 = 4'h5 == state ? _GEN_3572 : valid_3_6; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3855 = 4'h5 == state ? _GEN_3573 : valid_3_7; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3856 = 4'h5 == state ? _GEN_3574 : valid_3_8; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3857 = 4'h5 == state ? _GEN_3575 : valid_3_9; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3858 = 4'h5 == state ? _GEN_3576 : valid_3_10; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3859 = 4'h5 == state ? _GEN_3577 : valid_3_11; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3860 = 4'h5 == state ? _GEN_3578 : valid_3_12; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3861 = 4'h5 == state ? _GEN_3579 : valid_3_13; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3862 = 4'h5 == state ? _GEN_3580 : valid_3_14; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_3863 = 4'h5 == state ? _GEN_3581 : valid_3_15; // @[d_cache.scala 87:18 32:26]
  wire [511:0] _GEN_3864 = 4'h5 == state ? _GEN_3582 : _GEN_3653; // @[d_cache.scala 87:18]
  wire [41:0] _GEN_3865 = 4'h5 == state ? _GEN_3583 : {{10'd0}, write_back_addr}; // @[d_cache.scala 87:18 45:34]
  wire  _GEN_3866 = 4'h5 == state ? _GEN_3584 : dirty_0_0; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3867 = 4'h5 == state ? _GEN_3585 : dirty_0_1; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3868 = 4'h5 == state ? _GEN_3586 : dirty_0_2; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3869 = 4'h5 == state ? _GEN_3587 : dirty_0_3; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3870 = 4'h5 == state ? _GEN_3588 : dirty_0_4; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3871 = 4'h5 == state ? _GEN_3589 : dirty_0_5; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3872 = 4'h5 == state ? _GEN_3590 : dirty_0_6; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3873 = 4'h5 == state ? _GEN_3591 : dirty_0_7; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3874 = 4'h5 == state ? _GEN_3592 : dirty_0_8; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3875 = 4'h5 == state ? _GEN_3593 : dirty_0_9; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3876 = 4'h5 == state ? _GEN_3594 : dirty_0_10; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3877 = 4'h5 == state ? _GEN_3595 : dirty_0_11; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3878 = 4'h5 == state ? _GEN_3596 : dirty_0_12; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3879 = 4'h5 == state ? _GEN_3597 : dirty_0_13; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3880 = 4'h5 == state ? _GEN_3598 : dirty_0_14; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3881 = 4'h5 == state ? _GEN_3599 : dirty_0_15; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_3882 = 4'h5 == state ? _GEN_3600 : dirty_1_0; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3883 = 4'h5 == state ? _GEN_3601 : dirty_1_1; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3884 = 4'h5 == state ? _GEN_3602 : dirty_1_2; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3885 = 4'h5 == state ? _GEN_3603 : dirty_1_3; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3886 = 4'h5 == state ? _GEN_3604 : dirty_1_4; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3887 = 4'h5 == state ? _GEN_3605 : dirty_1_5; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3888 = 4'h5 == state ? _GEN_3606 : dirty_1_6; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3889 = 4'h5 == state ? _GEN_3607 : dirty_1_7; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3890 = 4'h5 == state ? _GEN_3608 : dirty_1_8; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3891 = 4'h5 == state ? _GEN_3609 : dirty_1_9; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3892 = 4'h5 == state ? _GEN_3610 : dirty_1_10; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3893 = 4'h5 == state ? _GEN_3611 : dirty_1_11; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3894 = 4'h5 == state ? _GEN_3612 : dirty_1_12; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3895 = 4'h5 == state ? _GEN_3613 : dirty_1_13; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3896 = 4'h5 == state ? _GEN_3614 : dirty_1_14; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3897 = 4'h5 == state ? _GEN_3615 : dirty_1_15; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_3898 = 4'h5 == state ? _GEN_3616 : dirty_2_0; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3899 = 4'h5 == state ? _GEN_3617 : dirty_2_1; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3900 = 4'h5 == state ? _GEN_3618 : dirty_2_2; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3901 = 4'h5 == state ? _GEN_3619 : dirty_2_3; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3902 = 4'h5 == state ? _GEN_3620 : dirty_2_4; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3903 = 4'h5 == state ? _GEN_3621 : dirty_2_5; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3904 = 4'h5 == state ? _GEN_3622 : dirty_2_6; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3905 = 4'h5 == state ? _GEN_3623 : dirty_2_7; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3906 = 4'h5 == state ? _GEN_3624 : dirty_2_8; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3907 = 4'h5 == state ? _GEN_3625 : dirty_2_9; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3908 = 4'h5 == state ? _GEN_3626 : dirty_2_10; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3909 = 4'h5 == state ? _GEN_3627 : dirty_2_11; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3910 = 4'h5 == state ? _GEN_3628 : dirty_2_12; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3911 = 4'h5 == state ? _GEN_3629 : dirty_2_13; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3912 = 4'h5 == state ? _GEN_3630 : dirty_2_14; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3913 = 4'h5 == state ? _GEN_3631 : dirty_2_15; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_3914 = 4'h5 == state ? _GEN_3632 : dirty_3_0; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3915 = 4'h5 == state ? _GEN_3633 : dirty_3_1; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3916 = 4'h5 == state ? _GEN_3634 : dirty_3_2; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3917 = 4'h5 == state ? _GEN_3635 : dirty_3_3; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3918 = 4'h5 == state ? _GEN_3636 : dirty_3_4; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3919 = 4'h5 == state ? _GEN_3637 : dirty_3_5; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3920 = 4'h5 == state ? _GEN_3638 : dirty_3_6; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3921 = 4'h5 == state ? _GEN_3639 : dirty_3_7; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3922 = 4'h5 == state ? _GEN_3640 : dirty_3_8; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3923 = 4'h5 == state ? _GEN_3641 : dirty_3_9; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3924 = 4'h5 == state ? _GEN_3642 : dirty_3_10; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3925 = 4'h5 == state ? _GEN_3643 : dirty_3_11; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3926 = 4'h5 == state ? _GEN_3644 : dirty_3_12; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3927 = 4'h5 == state ? _GEN_3645 : dirty_3_13; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3928 = 4'h5 == state ? _GEN_3646 : dirty_3_14; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_3929 = 4'h5 == state ? _GEN_3647 : dirty_3_15; // @[d_cache.scala 87:18 37:26]
  wire [3:0] _GEN_3930 = 4'h4 == state ? _GEN_670 : _GEN_3655; // @[d_cache.scala 87:18]
  wire [511:0] _GEN_3931 = 4'h4 == state ? ram_0_0 : _GEN_3656; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3932 = 4'h4 == state ? ram_0_1 : _GEN_3657; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3933 = 4'h4 == state ? ram_0_2 : _GEN_3658; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3934 = 4'h4 == state ? ram_0_3 : _GEN_3659; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3935 = 4'h4 == state ? ram_0_4 : _GEN_3660; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3936 = 4'h4 == state ? ram_0_5 : _GEN_3661; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3937 = 4'h4 == state ? ram_0_6 : _GEN_3662; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3938 = 4'h4 == state ? ram_0_7 : _GEN_3663; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3939 = 4'h4 == state ? ram_0_8 : _GEN_3664; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3940 = 4'h4 == state ? ram_0_9 : _GEN_3665; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3941 = 4'h4 == state ? ram_0_10 : _GEN_3666; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3942 = 4'h4 == state ? ram_0_11 : _GEN_3667; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3943 = 4'h4 == state ? ram_0_12 : _GEN_3668; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3944 = 4'h4 == state ? ram_0_13 : _GEN_3669; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3945 = 4'h4 == state ? ram_0_14 : _GEN_3670; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_3946 = 4'h4 == state ? ram_0_15 : _GEN_3671; // @[d_cache.scala 87:18 19:24]
  wire [31:0] _GEN_3947 = 4'h4 == state ? tag_0_0 : _GEN_3672; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3948 = 4'h4 == state ? tag_0_1 : _GEN_3673; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3949 = 4'h4 == state ? tag_0_2 : _GEN_3674; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3950 = 4'h4 == state ? tag_0_3 : _GEN_3675; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3951 = 4'h4 == state ? tag_0_4 : _GEN_3676; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3952 = 4'h4 == state ? tag_0_5 : _GEN_3677; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3953 = 4'h4 == state ? tag_0_6 : _GEN_3678; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3954 = 4'h4 == state ? tag_0_7 : _GEN_3679; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3955 = 4'h4 == state ? tag_0_8 : _GEN_3680; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3956 = 4'h4 == state ? tag_0_9 : _GEN_3681; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3957 = 4'h4 == state ? tag_0_10 : _GEN_3682; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3958 = 4'h4 == state ? tag_0_11 : _GEN_3683; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3959 = 4'h4 == state ? tag_0_12 : _GEN_3684; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3960 = 4'h4 == state ? tag_0_13 : _GEN_3685; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3961 = 4'h4 == state ? tag_0_14 : _GEN_3686; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_3962 = 4'h4 == state ? tag_0_15 : _GEN_3687; // @[d_cache.scala 87:18 24:24]
  wire  _GEN_3963 = 4'h4 == state ? valid_0_0 : _GEN_3688; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3964 = 4'h4 == state ? valid_0_1 : _GEN_3689; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3965 = 4'h4 == state ? valid_0_2 : _GEN_3690; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3966 = 4'h4 == state ? valid_0_3 : _GEN_3691; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3967 = 4'h4 == state ? valid_0_4 : _GEN_3692; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3968 = 4'h4 == state ? valid_0_5 : _GEN_3693; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3969 = 4'h4 == state ? valid_0_6 : _GEN_3694; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3970 = 4'h4 == state ? valid_0_7 : _GEN_3695; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3971 = 4'h4 == state ? valid_0_8 : _GEN_3696; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3972 = 4'h4 == state ? valid_0_9 : _GEN_3697; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3973 = 4'h4 == state ? valid_0_10 : _GEN_3698; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3974 = 4'h4 == state ? valid_0_11 : _GEN_3699; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3975 = 4'h4 == state ? valid_0_12 : _GEN_3700; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3976 = 4'h4 == state ? valid_0_13 : _GEN_3701; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3977 = 4'h4 == state ? valid_0_14 : _GEN_3702; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_3978 = 4'h4 == state ? valid_0_15 : _GEN_3703; // @[d_cache.scala 87:18 29:26]
  wire [7:0] _GEN_3979 = 4'h4 == state ? quene_0 : _GEN_3704; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3980 = 4'h4 == state ? quene_1 : _GEN_3705; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3981 = 4'h4 == state ? quene_2 : _GEN_3706; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3982 = 4'h4 == state ? quene_3 : _GEN_3707; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3983 = 4'h4 == state ? quene_4 : _GEN_3708; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3984 = 4'h4 == state ? quene_5 : _GEN_3709; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3985 = 4'h4 == state ? quene_6 : _GEN_3710; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3986 = 4'h4 == state ? quene_7 : _GEN_3711; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3987 = 4'h4 == state ? quene_8 : _GEN_3712; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3988 = 4'h4 == state ? quene_9 : _GEN_3713; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3989 = 4'h4 == state ? quene_10 : _GEN_3714; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3990 = 4'h4 == state ? quene_11 : _GEN_3715; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3991 = 4'h4 == state ? quene_12 : _GEN_3716; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3992 = 4'h4 == state ? quene_13 : _GEN_3717; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3993 = 4'h4 == state ? quene_14 : _GEN_3718; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_3994 = 4'h4 == state ? quene_15 : _GEN_3719; // @[d_cache.scala 87:18 52:24]
  wire [511:0] _GEN_3995 = 4'h4 == state ? ram_1_0 : _GEN_3720; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3996 = 4'h4 == state ? ram_1_1 : _GEN_3721; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3997 = 4'h4 == state ? ram_1_2 : _GEN_3722; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3998 = 4'h4 == state ? ram_1_3 : _GEN_3723; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_3999 = 4'h4 == state ? ram_1_4 : _GEN_3724; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4000 = 4'h4 == state ? ram_1_5 : _GEN_3725; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4001 = 4'h4 == state ? ram_1_6 : _GEN_3726; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4002 = 4'h4 == state ? ram_1_7 : _GEN_3727; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4003 = 4'h4 == state ? ram_1_8 : _GEN_3728; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4004 = 4'h4 == state ? ram_1_9 : _GEN_3729; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4005 = 4'h4 == state ? ram_1_10 : _GEN_3730; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4006 = 4'h4 == state ? ram_1_11 : _GEN_3731; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4007 = 4'h4 == state ? ram_1_12 : _GEN_3732; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4008 = 4'h4 == state ? ram_1_13 : _GEN_3733; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4009 = 4'h4 == state ? ram_1_14 : _GEN_3734; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4010 = 4'h4 == state ? ram_1_15 : _GEN_3735; // @[d_cache.scala 87:18 20:24]
  wire [31:0] _GEN_4011 = 4'h4 == state ? tag_1_0 : _GEN_3736; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4012 = 4'h4 == state ? tag_1_1 : _GEN_3737; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4013 = 4'h4 == state ? tag_1_2 : _GEN_3738; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4014 = 4'h4 == state ? tag_1_3 : _GEN_3739; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4015 = 4'h4 == state ? tag_1_4 : _GEN_3740; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4016 = 4'h4 == state ? tag_1_5 : _GEN_3741; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4017 = 4'h4 == state ? tag_1_6 : _GEN_3742; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4018 = 4'h4 == state ? tag_1_7 : _GEN_3743; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4019 = 4'h4 == state ? tag_1_8 : _GEN_3744; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4020 = 4'h4 == state ? tag_1_9 : _GEN_3745; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4021 = 4'h4 == state ? tag_1_10 : _GEN_3746; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4022 = 4'h4 == state ? tag_1_11 : _GEN_3747; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4023 = 4'h4 == state ? tag_1_12 : _GEN_3748; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4024 = 4'h4 == state ? tag_1_13 : _GEN_3749; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4025 = 4'h4 == state ? tag_1_14 : _GEN_3750; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4026 = 4'h4 == state ? tag_1_15 : _GEN_3751; // @[d_cache.scala 87:18 25:24]
  wire  _GEN_4027 = 4'h4 == state ? valid_1_0 : _GEN_3752; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4028 = 4'h4 == state ? valid_1_1 : _GEN_3753; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4029 = 4'h4 == state ? valid_1_2 : _GEN_3754; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4030 = 4'h4 == state ? valid_1_3 : _GEN_3755; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4031 = 4'h4 == state ? valid_1_4 : _GEN_3756; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4032 = 4'h4 == state ? valid_1_5 : _GEN_3757; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4033 = 4'h4 == state ? valid_1_6 : _GEN_3758; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4034 = 4'h4 == state ? valid_1_7 : _GEN_3759; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4035 = 4'h4 == state ? valid_1_8 : _GEN_3760; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4036 = 4'h4 == state ? valid_1_9 : _GEN_3761; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4037 = 4'h4 == state ? valid_1_10 : _GEN_3762; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4038 = 4'h4 == state ? valid_1_11 : _GEN_3763; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4039 = 4'h4 == state ? valid_1_12 : _GEN_3764; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4040 = 4'h4 == state ? valid_1_13 : _GEN_3765; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4041 = 4'h4 == state ? valid_1_14 : _GEN_3766; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4042 = 4'h4 == state ? valid_1_15 : _GEN_3767; // @[d_cache.scala 87:18 30:26]
  wire [511:0] _GEN_4043 = 4'h4 == state ? ram_2_0 : _GEN_3768; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4044 = 4'h4 == state ? ram_2_1 : _GEN_3769; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4045 = 4'h4 == state ? ram_2_2 : _GEN_3770; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4046 = 4'h4 == state ? ram_2_3 : _GEN_3771; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4047 = 4'h4 == state ? ram_2_4 : _GEN_3772; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4048 = 4'h4 == state ? ram_2_5 : _GEN_3773; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4049 = 4'h4 == state ? ram_2_6 : _GEN_3774; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4050 = 4'h4 == state ? ram_2_7 : _GEN_3775; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4051 = 4'h4 == state ? ram_2_8 : _GEN_3776; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4052 = 4'h4 == state ? ram_2_9 : _GEN_3777; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4053 = 4'h4 == state ? ram_2_10 : _GEN_3778; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4054 = 4'h4 == state ? ram_2_11 : _GEN_3779; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4055 = 4'h4 == state ? ram_2_12 : _GEN_3780; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4056 = 4'h4 == state ? ram_2_13 : _GEN_3781; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4057 = 4'h4 == state ? ram_2_14 : _GEN_3782; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4058 = 4'h4 == state ? ram_2_15 : _GEN_3783; // @[d_cache.scala 87:18 21:24]
  wire [31:0] _GEN_4059 = 4'h4 == state ? tag_2_0 : _GEN_3784; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4060 = 4'h4 == state ? tag_2_1 : _GEN_3785; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4061 = 4'h4 == state ? tag_2_2 : _GEN_3786; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4062 = 4'h4 == state ? tag_2_3 : _GEN_3787; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4063 = 4'h4 == state ? tag_2_4 : _GEN_3788; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4064 = 4'h4 == state ? tag_2_5 : _GEN_3789; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4065 = 4'h4 == state ? tag_2_6 : _GEN_3790; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4066 = 4'h4 == state ? tag_2_7 : _GEN_3791; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4067 = 4'h4 == state ? tag_2_8 : _GEN_3792; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4068 = 4'h4 == state ? tag_2_9 : _GEN_3793; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4069 = 4'h4 == state ? tag_2_10 : _GEN_3794; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4070 = 4'h4 == state ? tag_2_11 : _GEN_3795; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4071 = 4'h4 == state ? tag_2_12 : _GEN_3796; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4072 = 4'h4 == state ? tag_2_13 : _GEN_3797; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4073 = 4'h4 == state ? tag_2_14 : _GEN_3798; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4074 = 4'h4 == state ? tag_2_15 : _GEN_3799; // @[d_cache.scala 87:18 26:24]
  wire  _GEN_4075 = 4'h4 == state ? valid_2_0 : _GEN_3800; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4076 = 4'h4 == state ? valid_2_1 : _GEN_3801; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4077 = 4'h4 == state ? valid_2_2 : _GEN_3802; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4078 = 4'h4 == state ? valid_2_3 : _GEN_3803; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4079 = 4'h4 == state ? valid_2_4 : _GEN_3804; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4080 = 4'h4 == state ? valid_2_5 : _GEN_3805; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4081 = 4'h4 == state ? valid_2_6 : _GEN_3806; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4082 = 4'h4 == state ? valid_2_7 : _GEN_3807; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4083 = 4'h4 == state ? valid_2_8 : _GEN_3808; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4084 = 4'h4 == state ? valid_2_9 : _GEN_3809; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4085 = 4'h4 == state ? valid_2_10 : _GEN_3810; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4086 = 4'h4 == state ? valid_2_11 : _GEN_3811; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4087 = 4'h4 == state ? valid_2_12 : _GEN_3812; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4088 = 4'h4 == state ? valid_2_13 : _GEN_3813; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4089 = 4'h4 == state ? valid_2_14 : _GEN_3814; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4090 = 4'h4 == state ? valid_2_15 : _GEN_3815; // @[d_cache.scala 87:18 31:26]
  wire [511:0] _GEN_4091 = 4'h4 == state ? ram_3_0 : _GEN_3816; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4092 = 4'h4 == state ? ram_3_1 : _GEN_3817; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4093 = 4'h4 == state ? ram_3_2 : _GEN_3818; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4094 = 4'h4 == state ? ram_3_3 : _GEN_3819; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4095 = 4'h4 == state ? ram_3_4 : _GEN_3820; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4096 = 4'h4 == state ? ram_3_5 : _GEN_3821; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4097 = 4'h4 == state ? ram_3_6 : _GEN_3822; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4098 = 4'h4 == state ? ram_3_7 : _GEN_3823; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4099 = 4'h4 == state ? ram_3_8 : _GEN_3824; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4100 = 4'h4 == state ? ram_3_9 : _GEN_3825; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4101 = 4'h4 == state ? ram_3_10 : _GEN_3826; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4102 = 4'h4 == state ? ram_3_11 : _GEN_3827; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4103 = 4'h4 == state ? ram_3_12 : _GEN_3828; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4104 = 4'h4 == state ? ram_3_13 : _GEN_3829; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4105 = 4'h4 == state ? ram_3_14 : _GEN_3830; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4106 = 4'h4 == state ? ram_3_15 : _GEN_3831; // @[d_cache.scala 87:18 22:24]
  wire [31:0] _GEN_4107 = 4'h4 == state ? tag_3_0 : _GEN_3832; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4108 = 4'h4 == state ? tag_3_1 : _GEN_3833; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4109 = 4'h4 == state ? tag_3_2 : _GEN_3834; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4110 = 4'h4 == state ? tag_3_3 : _GEN_3835; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4111 = 4'h4 == state ? tag_3_4 : _GEN_3836; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4112 = 4'h4 == state ? tag_3_5 : _GEN_3837; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4113 = 4'h4 == state ? tag_3_6 : _GEN_3838; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4114 = 4'h4 == state ? tag_3_7 : _GEN_3839; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4115 = 4'h4 == state ? tag_3_8 : _GEN_3840; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4116 = 4'h4 == state ? tag_3_9 : _GEN_3841; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4117 = 4'h4 == state ? tag_3_10 : _GEN_3842; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4118 = 4'h4 == state ? tag_3_11 : _GEN_3843; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4119 = 4'h4 == state ? tag_3_12 : _GEN_3844; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4120 = 4'h4 == state ? tag_3_13 : _GEN_3845; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4121 = 4'h4 == state ? tag_3_14 : _GEN_3846; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4122 = 4'h4 == state ? tag_3_15 : _GEN_3847; // @[d_cache.scala 87:18 27:24]
  wire  _GEN_4123 = 4'h4 == state ? valid_3_0 : _GEN_3848; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4124 = 4'h4 == state ? valid_3_1 : _GEN_3849; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4125 = 4'h4 == state ? valid_3_2 : _GEN_3850; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4126 = 4'h4 == state ? valid_3_3 : _GEN_3851; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4127 = 4'h4 == state ? valid_3_4 : _GEN_3852; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4128 = 4'h4 == state ? valid_3_5 : _GEN_3853; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4129 = 4'h4 == state ? valid_3_6 : _GEN_3854; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4130 = 4'h4 == state ? valid_3_7 : _GEN_3855; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4131 = 4'h4 == state ? valid_3_8 : _GEN_3856; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4132 = 4'h4 == state ? valid_3_9 : _GEN_3857; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4133 = 4'h4 == state ? valid_3_10 : _GEN_3858; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4134 = 4'h4 == state ? valid_3_11 : _GEN_3859; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4135 = 4'h4 == state ? valid_3_12 : _GEN_3860; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4136 = 4'h4 == state ? valid_3_13 : _GEN_3861; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4137 = 4'h4 == state ? valid_3_14 : _GEN_3862; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4138 = 4'h4 == state ? valid_3_15 : _GEN_3863; // @[d_cache.scala 87:18 32:26]
  wire [511:0] _GEN_4139 = 4'h4 == state ? write_back_data : _GEN_3864; // @[d_cache.scala 87:18 44:34]
  wire [41:0] _GEN_4140 = 4'h4 == state ? {{10'd0}, write_back_addr} : _GEN_3865; // @[d_cache.scala 87:18 45:34]
  wire  _GEN_4141 = 4'h4 == state ? dirty_0_0 : _GEN_3866; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4142 = 4'h4 == state ? dirty_0_1 : _GEN_3867; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4143 = 4'h4 == state ? dirty_0_2 : _GEN_3868; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4144 = 4'h4 == state ? dirty_0_3 : _GEN_3869; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4145 = 4'h4 == state ? dirty_0_4 : _GEN_3870; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4146 = 4'h4 == state ? dirty_0_5 : _GEN_3871; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4147 = 4'h4 == state ? dirty_0_6 : _GEN_3872; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4148 = 4'h4 == state ? dirty_0_7 : _GEN_3873; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4149 = 4'h4 == state ? dirty_0_8 : _GEN_3874; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4150 = 4'h4 == state ? dirty_0_9 : _GEN_3875; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4151 = 4'h4 == state ? dirty_0_10 : _GEN_3876; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4152 = 4'h4 == state ? dirty_0_11 : _GEN_3877; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4153 = 4'h4 == state ? dirty_0_12 : _GEN_3878; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4154 = 4'h4 == state ? dirty_0_13 : _GEN_3879; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4155 = 4'h4 == state ? dirty_0_14 : _GEN_3880; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4156 = 4'h4 == state ? dirty_0_15 : _GEN_3881; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4157 = 4'h4 == state ? dirty_1_0 : _GEN_3882; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4158 = 4'h4 == state ? dirty_1_1 : _GEN_3883; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4159 = 4'h4 == state ? dirty_1_2 : _GEN_3884; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4160 = 4'h4 == state ? dirty_1_3 : _GEN_3885; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4161 = 4'h4 == state ? dirty_1_4 : _GEN_3886; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4162 = 4'h4 == state ? dirty_1_5 : _GEN_3887; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4163 = 4'h4 == state ? dirty_1_6 : _GEN_3888; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4164 = 4'h4 == state ? dirty_1_7 : _GEN_3889; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4165 = 4'h4 == state ? dirty_1_8 : _GEN_3890; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4166 = 4'h4 == state ? dirty_1_9 : _GEN_3891; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4167 = 4'h4 == state ? dirty_1_10 : _GEN_3892; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4168 = 4'h4 == state ? dirty_1_11 : _GEN_3893; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4169 = 4'h4 == state ? dirty_1_12 : _GEN_3894; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4170 = 4'h4 == state ? dirty_1_13 : _GEN_3895; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4171 = 4'h4 == state ? dirty_1_14 : _GEN_3896; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4172 = 4'h4 == state ? dirty_1_15 : _GEN_3897; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4173 = 4'h4 == state ? dirty_2_0 : _GEN_3898; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4174 = 4'h4 == state ? dirty_2_1 : _GEN_3899; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4175 = 4'h4 == state ? dirty_2_2 : _GEN_3900; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4176 = 4'h4 == state ? dirty_2_3 : _GEN_3901; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4177 = 4'h4 == state ? dirty_2_4 : _GEN_3902; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4178 = 4'h4 == state ? dirty_2_5 : _GEN_3903; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4179 = 4'h4 == state ? dirty_2_6 : _GEN_3904; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4180 = 4'h4 == state ? dirty_2_7 : _GEN_3905; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4181 = 4'h4 == state ? dirty_2_8 : _GEN_3906; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4182 = 4'h4 == state ? dirty_2_9 : _GEN_3907; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4183 = 4'h4 == state ? dirty_2_10 : _GEN_3908; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4184 = 4'h4 == state ? dirty_2_11 : _GEN_3909; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4185 = 4'h4 == state ? dirty_2_12 : _GEN_3910; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4186 = 4'h4 == state ? dirty_2_13 : _GEN_3911; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4187 = 4'h4 == state ? dirty_2_14 : _GEN_3912; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4188 = 4'h4 == state ? dirty_2_15 : _GEN_3913; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4189 = 4'h4 == state ? dirty_3_0 : _GEN_3914; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4190 = 4'h4 == state ? dirty_3_1 : _GEN_3915; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4191 = 4'h4 == state ? dirty_3_2 : _GEN_3916; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4192 = 4'h4 == state ? dirty_3_3 : _GEN_3917; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4193 = 4'h4 == state ? dirty_3_4 : _GEN_3918; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4194 = 4'h4 == state ? dirty_3_5 : _GEN_3919; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4195 = 4'h4 == state ? dirty_3_6 : _GEN_3920; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4196 = 4'h4 == state ? dirty_3_7 : _GEN_3921; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4197 = 4'h4 == state ? dirty_3_8 : _GEN_3922; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4198 = 4'h4 == state ? dirty_3_9 : _GEN_3923; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4199 = 4'h4 == state ? dirty_3_10 : _GEN_3924; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4200 = 4'h4 == state ? dirty_3_11 : _GEN_3925; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4201 = 4'h4 == state ? dirty_3_12 : _GEN_3926; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4202 = 4'h4 == state ? dirty_3_13 : _GEN_3927; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4203 = 4'h4 == state ? dirty_3_14 : _GEN_3928; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4204 = 4'h4 == state ? dirty_3_15 : _GEN_3929; // @[d_cache.scala 87:18 37:26]
  wire [63:0] _GEN_4205 = 4'h3 == state ? _GEN_660 : receive_data_0; // @[d_cache.scala 87:18 50:31]
  wire [63:0] _GEN_4206 = 4'h3 == state ? _GEN_661 : receive_data_1; // @[d_cache.scala 87:18 50:31]
  wire [63:0] _GEN_4207 = 4'h3 == state ? _GEN_662 : receive_data_2; // @[d_cache.scala 87:18 50:31]
  wire [63:0] _GEN_4208 = 4'h3 == state ? _GEN_663 : receive_data_3; // @[d_cache.scala 87:18 50:31]
  wire [63:0] _GEN_4209 = 4'h3 == state ? _GEN_664 : receive_data_4; // @[d_cache.scala 87:18 50:31]
  wire [63:0] _GEN_4210 = 4'h3 == state ? _GEN_665 : receive_data_5; // @[d_cache.scala 87:18 50:31]
  wire [63:0] _GEN_4211 = 4'h3 == state ? _GEN_666 : receive_data_6; // @[d_cache.scala 87:18 50:31]
  wire [63:0] _GEN_4212 = 4'h3 == state ? _GEN_667 : receive_data_7; // @[d_cache.scala 87:18 50:31]
  wire [2:0] _GEN_4213 = 4'h3 == state ? _GEN_668 : receive_num; // @[d_cache.scala 87:18 51:30]
  wire [3:0] _GEN_4214 = 4'h3 == state ? _GEN_669 : _GEN_3930; // @[d_cache.scala 87:18]
  wire [511:0] _GEN_4215 = 4'h3 == state ? ram_0_0 : _GEN_3931; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4216 = 4'h3 == state ? ram_0_1 : _GEN_3932; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4217 = 4'h3 == state ? ram_0_2 : _GEN_3933; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4218 = 4'h3 == state ? ram_0_3 : _GEN_3934; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4219 = 4'h3 == state ? ram_0_4 : _GEN_3935; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4220 = 4'h3 == state ? ram_0_5 : _GEN_3936; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4221 = 4'h3 == state ? ram_0_6 : _GEN_3937; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4222 = 4'h3 == state ? ram_0_7 : _GEN_3938; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4223 = 4'h3 == state ? ram_0_8 : _GEN_3939; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4224 = 4'h3 == state ? ram_0_9 : _GEN_3940; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4225 = 4'h3 == state ? ram_0_10 : _GEN_3941; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4226 = 4'h3 == state ? ram_0_11 : _GEN_3942; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4227 = 4'h3 == state ? ram_0_12 : _GEN_3943; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4228 = 4'h3 == state ? ram_0_13 : _GEN_3944; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4229 = 4'h3 == state ? ram_0_14 : _GEN_3945; // @[d_cache.scala 87:18 19:24]
  wire [511:0] _GEN_4230 = 4'h3 == state ? ram_0_15 : _GEN_3946; // @[d_cache.scala 87:18 19:24]
  wire [31:0] _GEN_4231 = 4'h3 == state ? tag_0_0 : _GEN_3947; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4232 = 4'h3 == state ? tag_0_1 : _GEN_3948; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4233 = 4'h3 == state ? tag_0_2 : _GEN_3949; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4234 = 4'h3 == state ? tag_0_3 : _GEN_3950; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4235 = 4'h3 == state ? tag_0_4 : _GEN_3951; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4236 = 4'h3 == state ? tag_0_5 : _GEN_3952; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4237 = 4'h3 == state ? tag_0_6 : _GEN_3953; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4238 = 4'h3 == state ? tag_0_7 : _GEN_3954; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4239 = 4'h3 == state ? tag_0_8 : _GEN_3955; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4240 = 4'h3 == state ? tag_0_9 : _GEN_3956; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4241 = 4'h3 == state ? tag_0_10 : _GEN_3957; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4242 = 4'h3 == state ? tag_0_11 : _GEN_3958; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4243 = 4'h3 == state ? tag_0_12 : _GEN_3959; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4244 = 4'h3 == state ? tag_0_13 : _GEN_3960; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4245 = 4'h3 == state ? tag_0_14 : _GEN_3961; // @[d_cache.scala 87:18 24:24]
  wire [31:0] _GEN_4246 = 4'h3 == state ? tag_0_15 : _GEN_3962; // @[d_cache.scala 87:18 24:24]
  wire  _GEN_4247 = 4'h3 == state ? valid_0_0 : _GEN_3963; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4248 = 4'h3 == state ? valid_0_1 : _GEN_3964; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4249 = 4'h3 == state ? valid_0_2 : _GEN_3965; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4250 = 4'h3 == state ? valid_0_3 : _GEN_3966; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4251 = 4'h3 == state ? valid_0_4 : _GEN_3967; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4252 = 4'h3 == state ? valid_0_5 : _GEN_3968; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4253 = 4'h3 == state ? valid_0_6 : _GEN_3969; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4254 = 4'h3 == state ? valid_0_7 : _GEN_3970; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4255 = 4'h3 == state ? valid_0_8 : _GEN_3971; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4256 = 4'h3 == state ? valid_0_9 : _GEN_3972; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4257 = 4'h3 == state ? valid_0_10 : _GEN_3973; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4258 = 4'h3 == state ? valid_0_11 : _GEN_3974; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4259 = 4'h3 == state ? valid_0_12 : _GEN_3975; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4260 = 4'h3 == state ? valid_0_13 : _GEN_3976; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4261 = 4'h3 == state ? valid_0_14 : _GEN_3977; // @[d_cache.scala 87:18 29:26]
  wire  _GEN_4262 = 4'h3 == state ? valid_0_15 : _GEN_3978; // @[d_cache.scala 87:18 29:26]
  wire [7:0] _GEN_4263 = 4'h3 == state ? quene_0 : _GEN_3979; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4264 = 4'h3 == state ? quene_1 : _GEN_3980; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4265 = 4'h3 == state ? quene_2 : _GEN_3981; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4266 = 4'h3 == state ? quene_3 : _GEN_3982; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4267 = 4'h3 == state ? quene_4 : _GEN_3983; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4268 = 4'h3 == state ? quene_5 : _GEN_3984; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4269 = 4'h3 == state ? quene_6 : _GEN_3985; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4270 = 4'h3 == state ? quene_7 : _GEN_3986; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4271 = 4'h3 == state ? quene_8 : _GEN_3987; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4272 = 4'h3 == state ? quene_9 : _GEN_3988; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4273 = 4'h3 == state ? quene_10 : _GEN_3989; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4274 = 4'h3 == state ? quene_11 : _GEN_3990; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4275 = 4'h3 == state ? quene_12 : _GEN_3991; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4276 = 4'h3 == state ? quene_13 : _GEN_3992; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4277 = 4'h3 == state ? quene_14 : _GEN_3993; // @[d_cache.scala 87:18 52:24]
  wire [7:0] _GEN_4278 = 4'h3 == state ? quene_15 : _GEN_3994; // @[d_cache.scala 87:18 52:24]
  wire [511:0] _GEN_4279 = 4'h3 == state ? ram_1_0 : _GEN_3995; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4280 = 4'h3 == state ? ram_1_1 : _GEN_3996; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4281 = 4'h3 == state ? ram_1_2 : _GEN_3997; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4282 = 4'h3 == state ? ram_1_3 : _GEN_3998; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4283 = 4'h3 == state ? ram_1_4 : _GEN_3999; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4284 = 4'h3 == state ? ram_1_5 : _GEN_4000; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4285 = 4'h3 == state ? ram_1_6 : _GEN_4001; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4286 = 4'h3 == state ? ram_1_7 : _GEN_4002; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4287 = 4'h3 == state ? ram_1_8 : _GEN_4003; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4288 = 4'h3 == state ? ram_1_9 : _GEN_4004; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4289 = 4'h3 == state ? ram_1_10 : _GEN_4005; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4290 = 4'h3 == state ? ram_1_11 : _GEN_4006; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4291 = 4'h3 == state ? ram_1_12 : _GEN_4007; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4292 = 4'h3 == state ? ram_1_13 : _GEN_4008; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4293 = 4'h3 == state ? ram_1_14 : _GEN_4009; // @[d_cache.scala 87:18 20:24]
  wire [511:0] _GEN_4294 = 4'h3 == state ? ram_1_15 : _GEN_4010; // @[d_cache.scala 87:18 20:24]
  wire [31:0] _GEN_4295 = 4'h3 == state ? tag_1_0 : _GEN_4011; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4296 = 4'h3 == state ? tag_1_1 : _GEN_4012; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4297 = 4'h3 == state ? tag_1_2 : _GEN_4013; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4298 = 4'h3 == state ? tag_1_3 : _GEN_4014; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4299 = 4'h3 == state ? tag_1_4 : _GEN_4015; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4300 = 4'h3 == state ? tag_1_5 : _GEN_4016; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4301 = 4'h3 == state ? tag_1_6 : _GEN_4017; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4302 = 4'h3 == state ? tag_1_7 : _GEN_4018; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4303 = 4'h3 == state ? tag_1_8 : _GEN_4019; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4304 = 4'h3 == state ? tag_1_9 : _GEN_4020; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4305 = 4'h3 == state ? tag_1_10 : _GEN_4021; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4306 = 4'h3 == state ? tag_1_11 : _GEN_4022; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4307 = 4'h3 == state ? tag_1_12 : _GEN_4023; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4308 = 4'h3 == state ? tag_1_13 : _GEN_4024; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4309 = 4'h3 == state ? tag_1_14 : _GEN_4025; // @[d_cache.scala 87:18 25:24]
  wire [31:0] _GEN_4310 = 4'h3 == state ? tag_1_15 : _GEN_4026; // @[d_cache.scala 87:18 25:24]
  wire  _GEN_4311 = 4'h3 == state ? valid_1_0 : _GEN_4027; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4312 = 4'h3 == state ? valid_1_1 : _GEN_4028; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4313 = 4'h3 == state ? valid_1_2 : _GEN_4029; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4314 = 4'h3 == state ? valid_1_3 : _GEN_4030; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4315 = 4'h3 == state ? valid_1_4 : _GEN_4031; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4316 = 4'h3 == state ? valid_1_5 : _GEN_4032; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4317 = 4'h3 == state ? valid_1_6 : _GEN_4033; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4318 = 4'h3 == state ? valid_1_7 : _GEN_4034; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4319 = 4'h3 == state ? valid_1_8 : _GEN_4035; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4320 = 4'h3 == state ? valid_1_9 : _GEN_4036; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4321 = 4'h3 == state ? valid_1_10 : _GEN_4037; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4322 = 4'h3 == state ? valid_1_11 : _GEN_4038; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4323 = 4'h3 == state ? valid_1_12 : _GEN_4039; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4324 = 4'h3 == state ? valid_1_13 : _GEN_4040; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4325 = 4'h3 == state ? valid_1_14 : _GEN_4041; // @[d_cache.scala 87:18 30:26]
  wire  _GEN_4326 = 4'h3 == state ? valid_1_15 : _GEN_4042; // @[d_cache.scala 87:18 30:26]
  wire [511:0] _GEN_4327 = 4'h3 == state ? ram_2_0 : _GEN_4043; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4328 = 4'h3 == state ? ram_2_1 : _GEN_4044; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4329 = 4'h3 == state ? ram_2_2 : _GEN_4045; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4330 = 4'h3 == state ? ram_2_3 : _GEN_4046; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4331 = 4'h3 == state ? ram_2_4 : _GEN_4047; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4332 = 4'h3 == state ? ram_2_5 : _GEN_4048; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4333 = 4'h3 == state ? ram_2_6 : _GEN_4049; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4334 = 4'h3 == state ? ram_2_7 : _GEN_4050; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4335 = 4'h3 == state ? ram_2_8 : _GEN_4051; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4336 = 4'h3 == state ? ram_2_9 : _GEN_4052; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4337 = 4'h3 == state ? ram_2_10 : _GEN_4053; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4338 = 4'h3 == state ? ram_2_11 : _GEN_4054; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4339 = 4'h3 == state ? ram_2_12 : _GEN_4055; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4340 = 4'h3 == state ? ram_2_13 : _GEN_4056; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4341 = 4'h3 == state ? ram_2_14 : _GEN_4057; // @[d_cache.scala 87:18 21:24]
  wire [511:0] _GEN_4342 = 4'h3 == state ? ram_2_15 : _GEN_4058; // @[d_cache.scala 87:18 21:24]
  wire [31:0] _GEN_4343 = 4'h3 == state ? tag_2_0 : _GEN_4059; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4344 = 4'h3 == state ? tag_2_1 : _GEN_4060; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4345 = 4'h3 == state ? tag_2_2 : _GEN_4061; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4346 = 4'h3 == state ? tag_2_3 : _GEN_4062; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4347 = 4'h3 == state ? tag_2_4 : _GEN_4063; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4348 = 4'h3 == state ? tag_2_5 : _GEN_4064; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4349 = 4'h3 == state ? tag_2_6 : _GEN_4065; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4350 = 4'h3 == state ? tag_2_7 : _GEN_4066; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4351 = 4'h3 == state ? tag_2_8 : _GEN_4067; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4352 = 4'h3 == state ? tag_2_9 : _GEN_4068; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4353 = 4'h3 == state ? tag_2_10 : _GEN_4069; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4354 = 4'h3 == state ? tag_2_11 : _GEN_4070; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4355 = 4'h3 == state ? tag_2_12 : _GEN_4071; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4356 = 4'h3 == state ? tag_2_13 : _GEN_4072; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4357 = 4'h3 == state ? tag_2_14 : _GEN_4073; // @[d_cache.scala 87:18 26:24]
  wire [31:0] _GEN_4358 = 4'h3 == state ? tag_2_15 : _GEN_4074; // @[d_cache.scala 87:18 26:24]
  wire  _GEN_4359 = 4'h3 == state ? valid_2_0 : _GEN_4075; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4360 = 4'h3 == state ? valid_2_1 : _GEN_4076; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4361 = 4'h3 == state ? valid_2_2 : _GEN_4077; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4362 = 4'h3 == state ? valid_2_3 : _GEN_4078; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4363 = 4'h3 == state ? valid_2_4 : _GEN_4079; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4364 = 4'h3 == state ? valid_2_5 : _GEN_4080; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4365 = 4'h3 == state ? valid_2_6 : _GEN_4081; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4366 = 4'h3 == state ? valid_2_7 : _GEN_4082; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4367 = 4'h3 == state ? valid_2_8 : _GEN_4083; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4368 = 4'h3 == state ? valid_2_9 : _GEN_4084; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4369 = 4'h3 == state ? valid_2_10 : _GEN_4085; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4370 = 4'h3 == state ? valid_2_11 : _GEN_4086; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4371 = 4'h3 == state ? valid_2_12 : _GEN_4087; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4372 = 4'h3 == state ? valid_2_13 : _GEN_4088; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4373 = 4'h3 == state ? valid_2_14 : _GEN_4089; // @[d_cache.scala 87:18 31:26]
  wire  _GEN_4374 = 4'h3 == state ? valid_2_15 : _GEN_4090; // @[d_cache.scala 87:18 31:26]
  wire [511:0] _GEN_4375 = 4'h3 == state ? ram_3_0 : _GEN_4091; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4376 = 4'h3 == state ? ram_3_1 : _GEN_4092; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4377 = 4'h3 == state ? ram_3_2 : _GEN_4093; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4378 = 4'h3 == state ? ram_3_3 : _GEN_4094; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4379 = 4'h3 == state ? ram_3_4 : _GEN_4095; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4380 = 4'h3 == state ? ram_3_5 : _GEN_4096; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4381 = 4'h3 == state ? ram_3_6 : _GEN_4097; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4382 = 4'h3 == state ? ram_3_7 : _GEN_4098; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4383 = 4'h3 == state ? ram_3_8 : _GEN_4099; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4384 = 4'h3 == state ? ram_3_9 : _GEN_4100; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4385 = 4'h3 == state ? ram_3_10 : _GEN_4101; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4386 = 4'h3 == state ? ram_3_11 : _GEN_4102; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4387 = 4'h3 == state ? ram_3_12 : _GEN_4103; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4388 = 4'h3 == state ? ram_3_13 : _GEN_4104; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4389 = 4'h3 == state ? ram_3_14 : _GEN_4105; // @[d_cache.scala 87:18 22:24]
  wire [511:0] _GEN_4390 = 4'h3 == state ? ram_3_15 : _GEN_4106; // @[d_cache.scala 87:18 22:24]
  wire [31:0] _GEN_4391 = 4'h3 == state ? tag_3_0 : _GEN_4107; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4392 = 4'h3 == state ? tag_3_1 : _GEN_4108; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4393 = 4'h3 == state ? tag_3_2 : _GEN_4109; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4394 = 4'h3 == state ? tag_3_3 : _GEN_4110; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4395 = 4'h3 == state ? tag_3_4 : _GEN_4111; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4396 = 4'h3 == state ? tag_3_5 : _GEN_4112; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4397 = 4'h3 == state ? tag_3_6 : _GEN_4113; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4398 = 4'h3 == state ? tag_3_7 : _GEN_4114; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4399 = 4'h3 == state ? tag_3_8 : _GEN_4115; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4400 = 4'h3 == state ? tag_3_9 : _GEN_4116; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4401 = 4'h3 == state ? tag_3_10 : _GEN_4117; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4402 = 4'h3 == state ? tag_3_11 : _GEN_4118; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4403 = 4'h3 == state ? tag_3_12 : _GEN_4119; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4404 = 4'h3 == state ? tag_3_13 : _GEN_4120; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4405 = 4'h3 == state ? tag_3_14 : _GEN_4121; // @[d_cache.scala 87:18 27:24]
  wire [31:0] _GEN_4406 = 4'h3 == state ? tag_3_15 : _GEN_4122; // @[d_cache.scala 87:18 27:24]
  wire  _GEN_4407 = 4'h3 == state ? valid_3_0 : _GEN_4123; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4408 = 4'h3 == state ? valid_3_1 : _GEN_4124; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4409 = 4'h3 == state ? valid_3_2 : _GEN_4125; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4410 = 4'h3 == state ? valid_3_3 : _GEN_4126; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4411 = 4'h3 == state ? valid_3_4 : _GEN_4127; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4412 = 4'h3 == state ? valid_3_5 : _GEN_4128; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4413 = 4'h3 == state ? valid_3_6 : _GEN_4129; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4414 = 4'h3 == state ? valid_3_7 : _GEN_4130; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4415 = 4'h3 == state ? valid_3_8 : _GEN_4131; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4416 = 4'h3 == state ? valid_3_9 : _GEN_4132; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4417 = 4'h3 == state ? valid_3_10 : _GEN_4133; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4418 = 4'h3 == state ? valid_3_11 : _GEN_4134; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4419 = 4'h3 == state ? valid_3_12 : _GEN_4135; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4420 = 4'h3 == state ? valid_3_13 : _GEN_4136; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4421 = 4'h3 == state ? valid_3_14 : _GEN_4137; // @[d_cache.scala 87:18 32:26]
  wire  _GEN_4422 = 4'h3 == state ? valid_3_15 : _GEN_4138; // @[d_cache.scala 87:18 32:26]
  wire [511:0] _GEN_4423 = 4'h3 == state ? write_back_data : _GEN_4139; // @[d_cache.scala 87:18 44:34]
  wire [41:0] _GEN_4424 = 4'h3 == state ? {{10'd0}, write_back_addr} : _GEN_4140; // @[d_cache.scala 87:18 45:34]
  wire  _GEN_4425 = 4'h3 == state ? dirty_0_0 : _GEN_4141; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4426 = 4'h3 == state ? dirty_0_1 : _GEN_4142; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4427 = 4'h3 == state ? dirty_0_2 : _GEN_4143; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4428 = 4'h3 == state ? dirty_0_3 : _GEN_4144; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4429 = 4'h3 == state ? dirty_0_4 : _GEN_4145; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4430 = 4'h3 == state ? dirty_0_5 : _GEN_4146; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4431 = 4'h3 == state ? dirty_0_6 : _GEN_4147; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4432 = 4'h3 == state ? dirty_0_7 : _GEN_4148; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4433 = 4'h3 == state ? dirty_0_8 : _GEN_4149; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4434 = 4'h3 == state ? dirty_0_9 : _GEN_4150; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4435 = 4'h3 == state ? dirty_0_10 : _GEN_4151; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4436 = 4'h3 == state ? dirty_0_11 : _GEN_4152; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4437 = 4'h3 == state ? dirty_0_12 : _GEN_4153; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4438 = 4'h3 == state ? dirty_0_13 : _GEN_4154; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4439 = 4'h3 == state ? dirty_0_14 : _GEN_4155; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4440 = 4'h3 == state ? dirty_0_15 : _GEN_4156; // @[d_cache.scala 87:18 34:26]
  wire  _GEN_4441 = 4'h3 == state ? dirty_1_0 : _GEN_4157; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4442 = 4'h3 == state ? dirty_1_1 : _GEN_4158; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4443 = 4'h3 == state ? dirty_1_2 : _GEN_4159; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4444 = 4'h3 == state ? dirty_1_3 : _GEN_4160; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4445 = 4'h3 == state ? dirty_1_4 : _GEN_4161; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4446 = 4'h3 == state ? dirty_1_5 : _GEN_4162; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4447 = 4'h3 == state ? dirty_1_6 : _GEN_4163; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4448 = 4'h3 == state ? dirty_1_7 : _GEN_4164; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4449 = 4'h3 == state ? dirty_1_8 : _GEN_4165; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4450 = 4'h3 == state ? dirty_1_9 : _GEN_4166; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4451 = 4'h3 == state ? dirty_1_10 : _GEN_4167; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4452 = 4'h3 == state ? dirty_1_11 : _GEN_4168; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4453 = 4'h3 == state ? dirty_1_12 : _GEN_4169; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4454 = 4'h3 == state ? dirty_1_13 : _GEN_4170; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4455 = 4'h3 == state ? dirty_1_14 : _GEN_4171; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4456 = 4'h3 == state ? dirty_1_15 : _GEN_4172; // @[d_cache.scala 87:18 35:26]
  wire  _GEN_4457 = 4'h3 == state ? dirty_2_0 : _GEN_4173; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4458 = 4'h3 == state ? dirty_2_1 : _GEN_4174; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4459 = 4'h3 == state ? dirty_2_2 : _GEN_4175; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4460 = 4'h3 == state ? dirty_2_3 : _GEN_4176; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4461 = 4'h3 == state ? dirty_2_4 : _GEN_4177; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4462 = 4'h3 == state ? dirty_2_5 : _GEN_4178; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4463 = 4'h3 == state ? dirty_2_6 : _GEN_4179; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4464 = 4'h3 == state ? dirty_2_7 : _GEN_4180; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4465 = 4'h3 == state ? dirty_2_8 : _GEN_4181; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4466 = 4'h3 == state ? dirty_2_9 : _GEN_4182; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4467 = 4'h3 == state ? dirty_2_10 : _GEN_4183; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4468 = 4'h3 == state ? dirty_2_11 : _GEN_4184; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4469 = 4'h3 == state ? dirty_2_12 : _GEN_4185; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4470 = 4'h3 == state ? dirty_2_13 : _GEN_4186; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4471 = 4'h3 == state ? dirty_2_14 : _GEN_4187; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4472 = 4'h3 == state ? dirty_2_15 : _GEN_4188; // @[d_cache.scala 87:18 36:26]
  wire  _GEN_4473 = 4'h3 == state ? dirty_3_0 : _GEN_4189; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4474 = 4'h3 == state ? dirty_3_1 : _GEN_4190; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4475 = 4'h3 == state ? dirty_3_2 : _GEN_4191; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4476 = 4'h3 == state ? dirty_3_3 : _GEN_4192; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4477 = 4'h3 == state ? dirty_3_4 : _GEN_4193; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4478 = 4'h3 == state ? dirty_3_5 : _GEN_4194; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4479 = 4'h3 == state ? dirty_3_6 : _GEN_4195; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4480 = 4'h3 == state ? dirty_3_7 : _GEN_4196; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4481 = 4'h3 == state ? dirty_3_8 : _GEN_4197; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4482 = 4'h3 == state ? dirty_3_9 : _GEN_4198; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4483 = 4'h3 == state ? dirty_3_10 : _GEN_4199; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4484 = 4'h3 == state ? dirty_3_11 : _GEN_4200; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4485 = 4'h3 == state ? dirty_3_12 : _GEN_4201; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4486 = 4'h3 == state ? dirty_3_13 : _GEN_4202; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4487 = 4'h3 == state ? dirty_3_14 : _GEN_4203; // @[d_cache.scala 87:18 37:26]
  wire  _GEN_4488 = 4'h3 == state ? dirty_3_15 : _GEN_4204; // @[d_cache.scala 87:18 37:26]
  wire [41:0] _GEN_4772 = 4'h2 == state ? {{10'd0}, write_back_addr} : _GEN_4424; // @[d_cache.scala 87:18 45:34]
  wire [41:0] _GEN_5056 = 4'h1 == state ? {{10'd0}, write_back_addr} : _GEN_4772; // @[d_cache.scala 87:18 45:34]
  wire [41:0] _GEN_5340 = 4'h0 == state ? {{10'd0}, write_back_addr} : _GEN_5056; // @[d_cache.scala 87:18 45:34]
  wire [511:0] _io_to_lsu_rdata_T = _GEN_150 >> shift_bit; // @[d_cache.scala 298:56]
  wire [511:0] _io_to_lsu_rdata_T_1 = _GEN_198 >> shift_bit; // @[d_cache.scala 298:98]
  wire [511:0] _io_to_lsu_rdata_T_2 = _GEN_246 >> shift_bit; // @[d_cache.scala 298:140]
  wire [511:0] _io_to_lsu_rdata_T_3 = _GEN_294 >> shift_bit; // @[d_cache.scala 298:169]
  wire [511:0] _io_to_lsu_rdata_T_4 = way2_hit ? _io_to_lsu_rdata_T_2 : _io_to_lsu_rdata_T_3; // @[d_cache.scala 298:116]
  wire [511:0] _io_to_lsu_rdata_T_5 = way1_hit ? _io_to_lsu_rdata_T_1 : _io_to_lsu_rdata_T_4; // @[d_cache.scala 298:74]
  wire [511:0] _io_to_lsu_rdata_T_6 = way0_hit ? _io_to_lsu_rdata_T : _io_to_lsu_rdata_T_5; // @[d_cache.scala 298:32]
  wire [63:0] _GEN_5702 = {{32'd0}, io_from_lsu_araddr}; // @[d_cache.scala 340:49]
  wire [63:0] _io_to_axi_araddr_T = _GEN_5702 & 64'hffffffffffffffc0; // @[d_cache.scala 340:49]
  wire  _T_35 = state == 4'h7; // @[d_cache.scala 420:21]
  wire [63:0] _GEN_5342 = state == 4'h7 ? io_from_axi_rdata : 64'h0; // @[d_cache.scala 420:30 421:19 424:25]
  wire  _GEN_5344 = state == 4'h7 & io_from_axi_rvalid; // @[d_cache.scala 420:30 421:19 426:26]
  wire  _GEN_5346 = state == 4'h7 & io_from_axi_wready; // @[d_cache.scala 420:30 421:19 428:26]
  wire  _GEN_5352 = state == 4'h7 & io_from_lsu_arvalid; // @[d_cache.scala 420:30 422:19 431:27]
  wire [31:0] _GEN_5354 = state == 4'h7 ? io_from_lsu_awaddr : 32'h0; // @[d_cache.scala 420:30 422:19 437:26]
  wire  _GEN_5358 = state == 4'h7 & io_from_lsu_awvalid; // @[d_cache.scala 420:30 422:19 438:27]
  wire [63:0] _GEN_5359 = state == 4'h7 ? io_from_lsu_wdata : 64'h0; // @[d_cache.scala 420:30 422:19 442:25]
  wire [7:0] _GEN_5360 = state == 4'h7 ? io_from_lsu_wstrb : 8'h0; // @[d_cache.scala 420:30 422:19 443:25]
  wire  _GEN_5362 = state == 4'h7 & io_from_lsu_wvalid; // @[d_cache.scala 420:30 422:19 445:26]
  wire [63:0] _GEN_5364 = state == 4'h6 ? 64'h0 : _GEN_5342; // @[d_cache.scala 396:35 397:25]
  wire  _GEN_5366 = state == 4'h6 ? 1'h0 : _GEN_5344; // @[d_cache.scala 396:35 399:26]
  wire  _GEN_5368 = state == 4'h6 ? 1'h0 : _GEN_5346; // @[d_cache.scala 396:35 401:26]
  wire  _GEN_5371 = state == 4'h6 ? 1'h0 : _GEN_5352; // @[d_cache.scala 396:35 404:27]
  wire [31:0] _GEN_5372 = state == 4'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 396:35 405:26]
  wire [7:0] _GEN_5373 = state == 4'h6 ? 8'h7 : 8'h0; // @[d_cache.scala 396:35 406:25]
  wire  _GEN_5376 = state == 4'h6 ? 1'h0 : 1'h1; // @[d_cache.scala 396:35 409:26]
  wire [31:0] _GEN_5377 = state == 4'h6 ? write_back_addr : _GEN_5354; // @[d_cache.scala 396:35 410:26]
  wire  _GEN_5378 = state == 4'h6 | _GEN_5358; // @[d_cache.scala 396:35 411:27]
  wire [63:0] _GEN_5382 = state == 4'h6 ? write_back_data[63:0] : _GEN_5359; // @[d_cache.scala 396:35 415:25]
  wire [7:0] _GEN_5383 = state == 4'h6 ? 8'hff : _GEN_5360; // @[d_cache.scala 396:35 416:25]
  wire  _GEN_5385 = state == 4'h6 | _GEN_5362; // @[d_cache.scala 396:35 418:26]
  wire  _GEN_5386 = state == 4'h6 | _T_35; // @[d_cache.scala 396:35 419:26]
  wire [63:0] _GEN_5387 = state == 4'h4 | state == 4'h8 ? 64'h0 : _GEN_5364; // @[d_cache.scala 355:50 356:25]
  wire  _GEN_5389 = state == 4'h4 | state == 4'h8 ? 1'h0 : _GEN_5366; // @[d_cache.scala 355:50 358:26]
  wire  _GEN_5391 = state == 4'h4 | state == 4'h8 ? io_from_axi_wready : _GEN_5368; // @[d_cache.scala 355:50 360:26]
  wire  _GEN_5394 = state == 4'h4 | state == 4'h8 ? 1'h0 : _GEN_5371; // @[d_cache.scala 355:50 363:27]
  wire [31:0] _GEN_5395 = state == 4'h4 | state == 4'h8 ? 32'h0 : _GEN_5372; // @[d_cache.scala 355:50 364:26]
  wire [7:0] _GEN_5396 = state == 4'h4 | state == 4'h8 ? 8'h0 : _GEN_5373; // @[d_cache.scala 355:50 365:25]
  wire  _GEN_5399 = state == 4'h4 | state == 4'h8 | _GEN_5376; // @[d_cache.scala 355:50 368:26]
  wire [31:0] _GEN_5400 = state == 4'h4 | state == 4'h8 ? io_from_lsu_awaddr : _GEN_5377; // @[d_cache.scala 355:50 369:26]
  wire  _GEN_5401 = state == 4'h4 | state == 4'h8 ? io_from_lsu_awvalid : _GEN_5378; // @[d_cache.scala 355:50 370:27]
  wire [63:0] _GEN_5405 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wdata : _GEN_5382; // @[d_cache.scala 355:50 374:25]
  wire [7:0] _GEN_5406 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wstrb : _GEN_5383; // @[d_cache.scala 355:50 375:25]
  wire  _GEN_5408 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wvalid : _GEN_5385; // @[d_cache.scala 355:50 377:26]
  wire  _GEN_5409 = state == 4'h4 | state == 4'h8 | _GEN_5386; // @[d_cache.scala 355:50 378:26]
  wire [63:0] _GEN_5410 = state == 4'h3 ? 64'h0 : _GEN_5387; // @[d_cache.scala 331:31 332:25]
  wire  _GEN_5412 = state == 4'h3 ? 1'h0 : _GEN_5389; // @[d_cache.scala 331:31 334:26]
  wire  _GEN_5414 = state == 4'h3 ? 1'h0 : _GEN_5391; // @[d_cache.scala 331:31 336:26]
  wire  _GEN_5417 = state == 4'h3 | _GEN_5394; // @[d_cache.scala 331:31 339:27]
  wire [63:0] _GEN_5418 = state == 4'h3 ? _io_to_axi_araddr_T : {{32'd0}, _GEN_5395}; // @[d_cache.scala 331:31 340:26]
  wire [7:0] _GEN_5419 = state == 4'h3 ? 8'h7 : _GEN_5396; // @[d_cache.scala 331:31 341:25]
  wire  _GEN_5422 = state == 4'h3 | _GEN_5399; // @[d_cache.scala 331:31 344:26]
  wire [31:0] _GEN_5423 = state == 4'h3 ? 32'h0 : _GEN_5400; // @[d_cache.scala 331:31 345:26]
  wire  _GEN_5424 = state == 4'h3 ? 1'h0 : _GEN_5401; // @[d_cache.scala 331:31 346:27]
  wire [7:0] _GEN_5425 = state == 4'h3 ? 8'h0 : _GEN_5396; // @[d_cache.scala 331:31 347:25]
  wire [63:0] _GEN_5428 = state == 4'h3 ? 64'h0 : _GEN_5405; // @[d_cache.scala 331:31 350:25]
  wire [7:0] _GEN_5429 = state == 4'h3 ? 8'h0 : _GEN_5406; // @[d_cache.scala 331:31 351:25]
  wire  _GEN_5431 = state == 4'h3 ? 1'h0 : _GEN_5408; // @[d_cache.scala 331:31 353:26]
  wire  _GEN_5432 = state == 4'h3 ? 1'h0 : _GEN_5409; // @[d_cache.scala 331:31 354:26]
  wire  _GEN_5433 = state == 4'h2 ? 1'h0 : _GEN_5417; // @[d_cache.scala 305:33 306:27]
  wire [63:0] _GEN_5434 = state == 4'h2 ? {{32'd0}, io_from_lsu_araddr} : _GEN_5418; // @[d_cache.scala 305:33 307:26]
  wire [7:0] _GEN_5435 = state == 4'h2 ? 8'h0 : _GEN_5419; // @[d_cache.scala 305:33 308:25]
  wire  _GEN_5438 = state == 4'h2 ? 1'h0 : _GEN_5422; // @[d_cache.scala 305:33 311:26]
  wire [31:0] _GEN_5439 = state == 4'h2 ? 32'h0 : _GEN_5423; // @[d_cache.scala 305:33 312:26]
  wire  _GEN_5440 = state == 4'h2 ? 1'h0 : _GEN_5424; // @[d_cache.scala 305:33 313:27]
  wire [7:0] _GEN_5441 = state == 4'h2 ? 8'h0 : _GEN_5425; // @[d_cache.scala 305:33 314:25]
  wire [63:0] _GEN_5444 = state == 4'h2 ? 64'h0 : _GEN_5428; // @[d_cache.scala 305:33 317:25]
  wire [7:0] _GEN_5445 = state == 4'h2 ? 8'h0 : _GEN_5429; // @[d_cache.scala 305:33 318:25]
  wire  _GEN_5447 = state == 4'h2 ? 1'h0 : _GEN_5431; // @[d_cache.scala 305:33 320:26]
  wire  _GEN_5448 = state == 4'h2 ? 1'h0 : _GEN_5432; // @[d_cache.scala 305:33 321:26]
  wire [63:0] _GEN_5449 = state == 4'h2 ? 64'h0 : _GEN_5410; // @[d_cache.scala 305:33 323:25]
  wire  _GEN_5451 = state == 4'h2 ? 1'h0 : _GEN_5412; // @[d_cache.scala 305:33 325:26]
  wire  _GEN_5453 = state == 4'h2 ? _T_6 : _GEN_5414; // @[d_cache.scala 305:33 327:26]
  wire [63:0] _GEN_5457 = state == 4'h1 ? {{32'd0}, io_from_lsu_araddr} : _GEN_5434; // @[d_cache.scala 281:27 283:26]
  wire [511:0] _GEN_5472 = state == 4'h1 ? _io_to_lsu_rdata_T_6 : {{448'd0}, _GEN_5449}; // @[d_cache.scala 281:27 298:25]
  wire [41:0] _GEN_5703 = reset ? 42'h0 : _GEN_5340; // @[d_cache.scala 45:{34,34}]
  assign io_to_lsu_rdata = _GEN_5472[63:0];
  assign io_to_lsu_rvalid = state == 4'h1 ? _T_6 : _GEN_5451; // @[d_cache.scala 281:27 300:26]
  assign io_to_lsu_wready = state == 4'h1 ? 1'h0 : _GEN_5453; // @[d_cache.scala 281:27 302:26]
  assign io_to_axi_araddr = _GEN_5457[31:0];
  assign io_to_axi_arlen = state == 4'h1 ? 8'h0 : _GEN_5435; // @[d_cache.scala 281:27 284:25]
  assign io_to_axi_arvalid = state == 4'h1 ? 1'h0 : _GEN_5433; // @[d_cache.scala 281:27 282:27]
  assign io_to_axi_rready = state == 4'h1 ? 1'h0 : _GEN_5438; // @[d_cache.scala 281:27 287:26]
  assign io_to_axi_awaddr = state == 4'h1 ? 32'h0 : _GEN_5439; // @[d_cache.scala 281:27 288:26]
  assign io_to_axi_awlen = state == 4'h1 ? 8'h0 : _GEN_5441; // @[d_cache.scala 281:27 290:25]
  assign io_to_axi_awvalid = state == 4'h1 ? 1'h0 : _GEN_5440; // @[d_cache.scala 281:27 289:27]
  assign io_to_axi_wdata = state == 4'h1 ? 64'h0 : _GEN_5444; // @[d_cache.scala 281:27 293:25]
  assign io_to_axi_wstrb = state == 4'h1 ? 8'h0 : _GEN_5445; // @[d_cache.scala 281:27 294:25]
  assign io_to_axi_wvalid = state == 4'h1 ? 1'h0 : _GEN_5447; // @[d_cache.scala 281:27 296:26]
  assign io_to_axi_bready = state == 4'h1 ? 1'h0 : _GEN_5448; // @[d_cache.scala 281:27 297:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_0 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_0 <= _GEN_523;
        end else begin
          ram_0_0 <= _GEN_4215;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_1 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_1 <= _GEN_524;
        end else begin
          ram_0_1 <= _GEN_4216;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_2 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_2 <= _GEN_525;
        end else begin
          ram_0_2 <= _GEN_4217;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_3 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_3 <= _GEN_526;
        end else begin
          ram_0_3 <= _GEN_4218;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_4 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_4 <= _GEN_527;
        end else begin
          ram_0_4 <= _GEN_4219;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_5 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_5 <= _GEN_528;
        end else begin
          ram_0_5 <= _GEN_4220;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_6 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_6 <= _GEN_529;
        end else begin
          ram_0_6 <= _GEN_4221;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_7 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_7 <= _GEN_530;
        end else begin
          ram_0_7 <= _GEN_4222;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_8 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_8 <= _GEN_531;
        end else begin
          ram_0_8 <= _GEN_4223;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_9 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_9 <= _GEN_532;
        end else begin
          ram_0_9 <= _GEN_4224;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_10 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_10 <= _GEN_533;
        end else begin
          ram_0_10 <= _GEN_4225;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_11 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_11 <= _GEN_534;
        end else begin
          ram_0_11 <= _GEN_4226;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_12 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_12 <= _GEN_535;
        end else begin
          ram_0_12 <= _GEN_4227;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_13 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_13 <= _GEN_536;
        end else begin
          ram_0_13 <= _GEN_4228;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_14 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_14 <= _GEN_537;
        end else begin
          ram_0_14 <= _GEN_4229;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_15 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_0_15 <= _GEN_538;
        end else begin
          ram_0_15 <= _GEN_4230;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_0 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_0 <= _GEN_555;
        end else begin
          ram_1_0 <= _GEN_4279;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_1 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_1 <= _GEN_556;
        end else begin
          ram_1_1 <= _GEN_4280;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_2 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_2 <= _GEN_557;
        end else begin
          ram_1_2 <= _GEN_4281;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_3 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_3 <= _GEN_558;
        end else begin
          ram_1_3 <= _GEN_4282;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_4 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_4 <= _GEN_559;
        end else begin
          ram_1_4 <= _GEN_4283;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_5 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_5 <= _GEN_560;
        end else begin
          ram_1_5 <= _GEN_4284;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_6 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_6 <= _GEN_561;
        end else begin
          ram_1_6 <= _GEN_4285;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_7 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_7 <= _GEN_562;
        end else begin
          ram_1_7 <= _GEN_4286;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_8 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_8 <= _GEN_563;
        end else begin
          ram_1_8 <= _GEN_4287;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_9 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_9 <= _GEN_564;
        end else begin
          ram_1_9 <= _GEN_4288;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_10 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_10 <= _GEN_565;
        end else begin
          ram_1_10 <= _GEN_4289;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_11 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_11 <= _GEN_566;
        end else begin
          ram_1_11 <= _GEN_4290;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_12 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_12 <= _GEN_567;
        end else begin
          ram_1_12 <= _GEN_4291;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_13 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_13 <= _GEN_568;
        end else begin
          ram_1_13 <= _GEN_4292;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_14 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_14 <= _GEN_569;
        end else begin
          ram_1_14 <= _GEN_4293;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_15 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_1_15 <= _GEN_570;
        end else begin
          ram_1_15 <= _GEN_4294;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_0 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_0 <= _GEN_587;
        end else begin
          ram_2_0 <= _GEN_4327;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_1 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_1 <= _GEN_588;
        end else begin
          ram_2_1 <= _GEN_4328;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_2 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_2 <= _GEN_589;
        end else begin
          ram_2_2 <= _GEN_4329;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_3 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_3 <= _GEN_590;
        end else begin
          ram_2_3 <= _GEN_4330;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_4 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_4 <= _GEN_591;
        end else begin
          ram_2_4 <= _GEN_4331;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_5 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_5 <= _GEN_592;
        end else begin
          ram_2_5 <= _GEN_4332;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_6 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_6 <= _GEN_593;
        end else begin
          ram_2_6 <= _GEN_4333;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_7 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_7 <= _GEN_594;
        end else begin
          ram_2_7 <= _GEN_4334;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_8 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_8 <= _GEN_595;
        end else begin
          ram_2_8 <= _GEN_4335;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_9 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_9 <= _GEN_596;
        end else begin
          ram_2_9 <= _GEN_4336;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_10 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_10 <= _GEN_597;
        end else begin
          ram_2_10 <= _GEN_4337;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_11 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_11 <= _GEN_598;
        end else begin
          ram_2_11 <= _GEN_4338;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_12 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_12 <= _GEN_599;
        end else begin
          ram_2_12 <= _GEN_4339;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_13 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_13 <= _GEN_600;
        end else begin
          ram_2_13 <= _GEN_4340;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_14 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_14 <= _GEN_601;
        end else begin
          ram_2_14 <= _GEN_4341;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_15 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_2_15 <= _GEN_602;
        end else begin
          ram_2_15 <= _GEN_4342;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_0 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_0 <= _GEN_619;
        end else begin
          ram_3_0 <= _GEN_4375;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_1 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_1 <= _GEN_620;
        end else begin
          ram_3_1 <= _GEN_4376;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_2 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_2 <= _GEN_621;
        end else begin
          ram_3_2 <= _GEN_4377;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_3 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_3 <= _GEN_622;
        end else begin
          ram_3_3 <= _GEN_4378;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_4 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_4 <= _GEN_623;
        end else begin
          ram_3_4 <= _GEN_4379;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_5 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_5 <= _GEN_624;
        end else begin
          ram_3_5 <= _GEN_4380;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_6 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_6 <= _GEN_625;
        end else begin
          ram_3_6 <= _GEN_4381;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_7 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_7 <= _GEN_626;
        end else begin
          ram_3_7 <= _GEN_4382;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_8 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_8 <= _GEN_627;
        end else begin
          ram_3_8 <= _GEN_4383;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_9 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_9 <= _GEN_628;
        end else begin
          ram_3_9 <= _GEN_4384;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_10 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_10 <= _GEN_629;
        end else begin
          ram_3_10 <= _GEN_4385;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_11 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_11 <= _GEN_630;
        end else begin
          ram_3_11 <= _GEN_4386;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_12 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_12 <= _GEN_631;
        end else begin
          ram_3_12 <= _GEN_4387;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_13 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_13 <= _GEN_632;
        end else begin
          ram_3_13 <= _GEN_4388;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_14 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_14 <= _GEN_633;
        end else begin
          ram_3_14 <= _GEN_4389;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_15 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          ram_3_15 <= _GEN_634;
        end else begin
          ram_3_15 <= _GEN_4390;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_0 <= _GEN_4231;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_1 <= _GEN_4232;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_2 <= _GEN_4233;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_3 <= _GEN_4234;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_4 <= _GEN_4235;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_5 <= _GEN_4236;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_6 <= _GEN_4237;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_7 <= _GEN_4238;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_8 <= _GEN_4239;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_9 <= _GEN_4240;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_10 <= _GEN_4241;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_11 <= _GEN_4242;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_12 <= _GEN_4243;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_13 <= _GEN_4244;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_14 <= _GEN_4245;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_0_15 <= _GEN_4246;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_0 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_0 <= _GEN_4295;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_1 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_1 <= _GEN_4296;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_2 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_2 <= _GEN_4297;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_3 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_3 <= _GEN_4298;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_4 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_4 <= _GEN_4299;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_5 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_5 <= _GEN_4300;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_6 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_6 <= _GEN_4301;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_7 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_7 <= _GEN_4302;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_8 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_8 <= _GEN_4303;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_9 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_9 <= _GEN_4304;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_10 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_10 <= _GEN_4305;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_11 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_11 <= _GEN_4306;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_12 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_12 <= _GEN_4307;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_13 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_13 <= _GEN_4308;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_14 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_14 <= _GEN_4309;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_15 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_1_15 <= _GEN_4310;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_0 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_0 <= _GEN_4343;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_1 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_1 <= _GEN_4344;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_2 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_2 <= _GEN_4345;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_3 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_3 <= _GEN_4346;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_4 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_4 <= _GEN_4347;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_5 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_5 <= _GEN_4348;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_6 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_6 <= _GEN_4349;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_7 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_7 <= _GEN_4350;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_8 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_8 <= _GEN_4351;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_9 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_9 <= _GEN_4352;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_10 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_10 <= _GEN_4353;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_11 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_11 <= _GEN_4354;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_12 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_12 <= _GEN_4355;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_13 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_13 <= _GEN_4356;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_14 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_14 <= _GEN_4357;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_15 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_2_15 <= _GEN_4358;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_0 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_0 <= _GEN_4391;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_1 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_1 <= _GEN_4392;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_2 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_2 <= _GEN_4393;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_3 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_3 <= _GEN_4394;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_4 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_4 <= _GEN_4395;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_5 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_5 <= _GEN_4396;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_6 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_6 <= _GEN_4397;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_7 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_7 <= _GEN_4398;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_8 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_8 <= _GEN_4399;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_9 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_9 <= _GEN_4400;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_10 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_10 <= _GEN_4401;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_11 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_11 <= _GEN_4402;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_12 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_12 <= _GEN_4403;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_13 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_13 <= _GEN_4404;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_14 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_14 <= _GEN_4405;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_15 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          tag_3_15 <= _GEN_4406;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_0 <= _GEN_4247;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_1 <= _GEN_4248;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_2 <= _GEN_4249;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_3 <= _GEN_4250;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_4 <= _GEN_4251;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_5 <= _GEN_4252;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_6 <= _GEN_4253;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_7 <= _GEN_4254;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_8 <= _GEN_4255;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_9 <= _GEN_4256;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_10 <= _GEN_4257;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_11 <= _GEN_4258;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_12 <= _GEN_4259;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_13 <= _GEN_4260;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_14 <= _GEN_4261;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_0_15 <= _GEN_4262;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_0 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_0 <= _GEN_4311;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_1 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_1 <= _GEN_4312;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_2 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_2 <= _GEN_4313;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_3 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_3 <= _GEN_4314;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_4 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_4 <= _GEN_4315;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_5 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_5 <= _GEN_4316;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_6 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_6 <= _GEN_4317;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_7 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_7 <= _GEN_4318;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_8 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_8 <= _GEN_4319;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_9 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_9 <= _GEN_4320;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_10 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_10 <= _GEN_4321;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_11 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_11 <= _GEN_4322;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_12 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_12 <= _GEN_4323;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_13 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_13 <= _GEN_4324;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_14 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_14 <= _GEN_4325;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_15 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_1_15 <= _GEN_4326;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_0 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_0 <= _GEN_4359;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_1 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_1 <= _GEN_4360;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_2 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_2 <= _GEN_4361;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_3 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_3 <= _GEN_4362;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_4 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_4 <= _GEN_4363;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_5 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_5 <= _GEN_4364;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_6 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_6 <= _GEN_4365;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_7 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_7 <= _GEN_4366;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_8 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_8 <= _GEN_4367;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_9 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_9 <= _GEN_4368;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_10 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_10 <= _GEN_4369;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_11 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_11 <= _GEN_4370;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_12 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_12 <= _GEN_4371;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_13 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_13 <= _GEN_4372;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_14 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_14 <= _GEN_4373;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_15 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_2_15 <= _GEN_4374;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_0 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_0 <= _GEN_4407;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_1 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_1 <= _GEN_4408;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_2 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_2 <= _GEN_4409;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_3 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_3 <= _GEN_4410;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_4 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_4 <= _GEN_4411;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_5 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_5 <= _GEN_4412;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_6 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_6 <= _GEN_4413;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_7 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_7 <= _GEN_4414;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_8 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_8 <= _GEN_4415;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_9 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_9 <= _GEN_4416;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_10 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_10 <= _GEN_4417;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_11 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_11 <= _GEN_4418;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_12 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_12 <= _GEN_4419;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_13 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_13 <= _GEN_4420;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_14 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_14 <= _GEN_4421;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_15 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          valid_3_15 <= _GEN_4422;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_0 <= _GEN_539;
        end else begin
          dirty_0_0 <= _GEN_4425;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_1 <= _GEN_540;
        end else begin
          dirty_0_1 <= _GEN_4426;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_2 <= _GEN_541;
        end else begin
          dirty_0_2 <= _GEN_4427;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_3 <= _GEN_542;
        end else begin
          dirty_0_3 <= _GEN_4428;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_4 <= _GEN_543;
        end else begin
          dirty_0_4 <= _GEN_4429;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_5 <= _GEN_544;
        end else begin
          dirty_0_5 <= _GEN_4430;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_6 <= _GEN_545;
        end else begin
          dirty_0_6 <= _GEN_4431;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_7 <= _GEN_546;
        end else begin
          dirty_0_7 <= _GEN_4432;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_8 <= _GEN_547;
        end else begin
          dirty_0_8 <= _GEN_4433;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_9 <= _GEN_548;
        end else begin
          dirty_0_9 <= _GEN_4434;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_10 <= _GEN_549;
        end else begin
          dirty_0_10 <= _GEN_4435;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_11 <= _GEN_550;
        end else begin
          dirty_0_11 <= _GEN_4436;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_12 <= _GEN_551;
        end else begin
          dirty_0_12 <= _GEN_4437;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_13 <= _GEN_552;
        end else begin
          dirty_0_13 <= _GEN_4438;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_14 <= _GEN_553;
        end else begin
          dirty_0_14 <= _GEN_4439;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_0_15 <= _GEN_554;
        end else begin
          dirty_0_15 <= _GEN_4440;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_0 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_0 <= _GEN_571;
        end else begin
          dirty_1_0 <= _GEN_4441;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_1 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_1 <= _GEN_572;
        end else begin
          dirty_1_1 <= _GEN_4442;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_2 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_2 <= _GEN_573;
        end else begin
          dirty_1_2 <= _GEN_4443;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_3 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_3 <= _GEN_574;
        end else begin
          dirty_1_3 <= _GEN_4444;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_4 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_4 <= _GEN_575;
        end else begin
          dirty_1_4 <= _GEN_4445;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_5 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_5 <= _GEN_576;
        end else begin
          dirty_1_5 <= _GEN_4446;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_6 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_6 <= _GEN_577;
        end else begin
          dirty_1_6 <= _GEN_4447;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_7 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_7 <= _GEN_578;
        end else begin
          dirty_1_7 <= _GEN_4448;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_8 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_8 <= _GEN_579;
        end else begin
          dirty_1_8 <= _GEN_4449;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_9 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_9 <= _GEN_580;
        end else begin
          dirty_1_9 <= _GEN_4450;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_10 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_10 <= _GEN_581;
        end else begin
          dirty_1_10 <= _GEN_4451;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_11 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_11 <= _GEN_582;
        end else begin
          dirty_1_11 <= _GEN_4452;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_12 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_12 <= _GEN_583;
        end else begin
          dirty_1_12 <= _GEN_4453;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_13 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_13 <= _GEN_584;
        end else begin
          dirty_1_13 <= _GEN_4454;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_14 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_14 <= _GEN_585;
        end else begin
          dirty_1_14 <= _GEN_4455;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_15 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_1_15 <= _GEN_586;
        end else begin
          dirty_1_15 <= _GEN_4456;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_0 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_0 <= _GEN_603;
        end else begin
          dirty_2_0 <= _GEN_4457;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_1 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_1 <= _GEN_604;
        end else begin
          dirty_2_1 <= _GEN_4458;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_2 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_2 <= _GEN_605;
        end else begin
          dirty_2_2 <= _GEN_4459;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_3 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_3 <= _GEN_606;
        end else begin
          dirty_2_3 <= _GEN_4460;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_4 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_4 <= _GEN_607;
        end else begin
          dirty_2_4 <= _GEN_4461;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_5 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_5 <= _GEN_608;
        end else begin
          dirty_2_5 <= _GEN_4462;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_6 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_6 <= _GEN_609;
        end else begin
          dirty_2_6 <= _GEN_4463;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_7 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_7 <= _GEN_610;
        end else begin
          dirty_2_7 <= _GEN_4464;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_8 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_8 <= _GEN_611;
        end else begin
          dirty_2_8 <= _GEN_4465;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_9 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_9 <= _GEN_612;
        end else begin
          dirty_2_9 <= _GEN_4466;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_10 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_10 <= _GEN_613;
        end else begin
          dirty_2_10 <= _GEN_4467;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_11 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_11 <= _GEN_614;
        end else begin
          dirty_2_11 <= _GEN_4468;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_12 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_12 <= _GEN_615;
        end else begin
          dirty_2_12 <= _GEN_4469;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_13 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_13 <= _GEN_616;
        end else begin
          dirty_2_13 <= _GEN_4470;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_14 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_14 <= _GEN_617;
        end else begin
          dirty_2_14 <= _GEN_4471;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_15 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_2_15 <= _GEN_618;
        end else begin
          dirty_2_15 <= _GEN_4472;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_0 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_0 <= _GEN_635;
        end else begin
          dirty_3_0 <= _GEN_4473;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_1 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_1 <= _GEN_636;
        end else begin
          dirty_3_1 <= _GEN_4474;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_2 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_2 <= _GEN_637;
        end else begin
          dirty_3_2 <= _GEN_4475;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_3 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_3 <= _GEN_638;
        end else begin
          dirty_3_3 <= _GEN_4476;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_4 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_4 <= _GEN_639;
        end else begin
          dirty_3_4 <= _GEN_4477;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_5 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_5 <= _GEN_640;
        end else begin
          dirty_3_5 <= _GEN_4478;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_6 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_6 <= _GEN_641;
        end else begin
          dirty_3_6 <= _GEN_4479;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_7 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_7 <= _GEN_642;
        end else begin
          dirty_3_7 <= _GEN_4480;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_8 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_8 <= _GEN_643;
        end else begin
          dirty_3_8 <= _GEN_4481;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_9 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_9 <= _GEN_644;
        end else begin
          dirty_3_9 <= _GEN_4482;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_10 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_10 <= _GEN_645;
        end else begin
          dirty_3_10 <= _GEN_4483;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_11 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_11 <= _GEN_646;
        end else begin
          dirty_3_11 <= _GEN_4484;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_12 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_12 <= _GEN_647;
        end else begin
          dirty_3_12 <= _GEN_4485;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_13 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_13 <= _GEN_648;
        end else begin
          dirty_3_13 <= _GEN_4486;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_14 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_14 <= _GEN_649;
        end else begin
          dirty_3_14 <= _GEN_4487;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_15 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (4'h2 == state) begin // @[d_cache.scala 87:18]
          dirty_3_15 <= _GEN_650;
        end else begin
          dirty_3_15 <= _GEN_4488;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 44:34]
      write_back_data <= 512'h0; // @[d_cache.scala 44:34]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          write_back_data <= _GEN_4423;
        end
      end
    end
    write_back_addr <= _GEN_5703[31:0]; // @[d_cache.scala 45:{34,34}]
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_0 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          receive_data_0 <= _GEN_4205;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_1 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          receive_data_1 <= _GEN_4206;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_2 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          receive_data_2 <= _GEN_4207;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_3 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          receive_data_3 <= _GEN_4208;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_4 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          receive_data_4 <= _GEN_4209;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_5 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          receive_data_5 <= _GEN_4210;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_6 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          receive_data_6 <= _GEN_4211;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_7 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          receive_data_7 <= _GEN_4212;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 51:30]
      receive_num <= 3'h0; // @[d_cache.scala 51:30]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (4'h1 == state) begin // @[d_cache.scala 87:18]
        if (!(way0_hit | way1_hit | way2_hit | way3_hit)) begin // @[d_cache.scala 105:57]
          receive_num <= 3'h0; // @[d_cache.scala 111:29]
        end
      end else if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
        receive_num <= _GEN_4213;
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_0 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_0 <= _GEN_4263;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_1 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_1 <= _GEN_4264;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_2 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_2 <= _GEN_4265;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_3 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_3 <= _GEN_4266;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_4 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_4 <= _GEN_4267;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_5 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_5 <= _GEN_4268;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_6 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_6 <= _GEN_4269;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_7 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_7 <= _GEN_4270;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_8 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_8 <= _GEN_4271;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_9 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_9 <= _GEN_4272;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_10 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_10 <= _GEN_4273;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_11 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_11 <= _GEN_4274;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_12 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_12 <= _GEN_4275;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_13 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_13 <= _GEN_4276;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_14 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_14 <= _GEN_4277;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_15 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 87:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 87:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 87:18]
          quene_15 <= _GEN_4278;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 82:24]
      state <= 4'h0; // @[d_cache.scala 82:24]
    end else if (4'h0 == state) begin // @[d_cache.scala 87:18]
      if (io_from_lsu_arvalid) begin // @[d_cache.scala 89:38]
        if (io_from_lsu_araddr >= 32'ha0000000) begin // @[d_cache.scala 90:58]
          state <= 4'h7; // @[d_cache.scala 91:27]
        end else begin
          state <= 4'h1; // @[d_cache.scala 93:27]
        end
      end else if (io_from_lsu_awvalid) begin // @[d_cache.scala 95:44]
        state <= _GEN_129;
      end
    end else if (4'h1 == state) begin // @[d_cache.scala 87:18]
      if (way0_hit | way1_hit | way2_hit | way3_hit) begin // @[d_cache.scala 105:57]
        state <= 4'h0;
      end else begin
        state <= 4'h3; // @[d_cache.scala 110:23]
      end
    end else if (4'h2 == state) begin // @[d_cache.scala 87:18]
      state <= _GEN_522;
    end else begin
      state <= _GEN_4214;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  ram_0_0 = _RAND_0[511:0];
  _RAND_1 = {16{`RANDOM}};
  ram_0_1 = _RAND_1[511:0];
  _RAND_2 = {16{`RANDOM}};
  ram_0_2 = _RAND_2[511:0];
  _RAND_3 = {16{`RANDOM}};
  ram_0_3 = _RAND_3[511:0];
  _RAND_4 = {16{`RANDOM}};
  ram_0_4 = _RAND_4[511:0];
  _RAND_5 = {16{`RANDOM}};
  ram_0_5 = _RAND_5[511:0];
  _RAND_6 = {16{`RANDOM}};
  ram_0_6 = _RAND_6[511:0];
  _RAND_7 = {16{`RANDOM}};
  ram_0_7 = _RAND_7[511:0];
  _RAND_8 = {16{`RANDOM}};
  ram_0_8 = _RAND_8[511:0];
  _RAND_9 = {16{`RANDOM}};
  ram_0_9 = _RAND_9[511:0];
  _RAND_10 = {16{`RANDOM}};
  ram_0_10 = _RAND_10[511:0];
  _RAND_11 = {16{`RANDOM}};
  ram_0_11 = _RAND_11[511:0];
  _RAND_12 = {16{`RANDOM}};
  ram_0_12 = _RAND_12[511:0];
  _RAND_13 = {16{`RANDOM}};
  ram_0_13 = _RAND_13[511:0];
  _RAND_14 = {16{`RANDOM}};
  ram_0_14 = _RAND_14[511:0];
  _RAND_15 = {16{`RANDOM}};
  ram_0_15 = _RAND_15[511:0];
  _RAND_16 = {16{`RANDOM}};
  ram_1_0 = _RAND_16[511:0];
  _RAND_17 = {16{`RANDOM}};
  ram_1_1 = _RAND_17[511:0];
  _RAND_18 = {16{`RANDOM}};
  ram_1_2 = _RAND_18[511:0];
  _RAND_19 = {16{`RANDOM}};
  ram_1_3 = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  ram_1_4 = _RAND_20[511:0];
  _RAND_21 = {16{`RANDOM}};
  ram_1_5 = _RAND_21[511:0];
  _RAND_22 = {16{`RANDOM}};
  ram_1_6 = _RAND_22[511:0];
  _RAND_23 = {16{`RANDOM}};
  ram_1_7 = _RAND_23[511:0];
  _RAND_24 = {16{`RANDOM}};
  ram_1_8 = _RAND_24[511:0];
  _RAND_25 = {16{`RANDOM}};
  ram_1_9 = _RAND_25[511:0];
  _RAND_26 = {16{`RANDOM}};
  ram_1_10 = _RAND_26[511:0];
  _RAND_27 = {16{`RANDOM}};
  ram_1_11 = _RAND_27[511:0];
  _RAND_28 = {16{`RANDOM}};
  ram_1_12 = _RAND_28[511:0];
  _RAND_29 = {16{`RANDOM}};
  ram_1_13 = _RAND_29[511:0];
  _RAND_30 = {16{`RANDOM}};
  ram_1_14 = _RAND_30[511:0];
  _RAND_31 = {16{`RANDOM}};
  ram_1_15 = _RAND_31[511:0];
  _RAND_32 = {16{`RANDOM}};
  ram_2_0 = _RAND_32[511:0];
  _RAND_33 = {16{`RANDOM}};
  ram_2_1 = _RAND_33[511:0];
  _RAND_34 = {16{`RANDOM}};
  ram_2_2 = _RAND_34[511:0];
  _RAND_35 = {16{`RANDOM}};
  ram_2_3 = _RAND_35[511:0];
  _RAND_36 = {16{`RANDOM}};
  ram_2_4 = _RAND_36[511:0];
  _RAND_37 = {16{`RANDOM}};
  ram_2_5 = _RAND_37[511:0];
  _RAND_38 = {16{`RANDOM}};
  ram_2_6 = _RAND_38[511:0];
  _RAND_39 = {16{`RANDOM}};
  ram_2_7 = _RAND_39[511:0];
  _RAND_40 = {16{`RANDOM}};
  ram_2_8 = _RAND_40[511:0];
  _RAND_41 = {16{`RANDOM}};
  ram_2_9 = _RAND_41[511:0];
  _RAND_42 = {16{`RANDOM}};
  ram_2_10 = _RAND_42[511:0];
  _RAND_43 = {16{`RANDOM}};
  ram_2_11 = _RAND_43[511:0];
  _RAND_44 = {16{`RANDOM}};
  ram_2_12 = _RAND_44[511:0];
  _RAND_45 = {16{`RANDOM}};
  ram_2_13 = _RAND_45[511:0];
  _RAND_46 = {16{`RANDOM}};
  ram_2_14 = _RAND_46[511:0];
  _RAND_47 = {16{`RANDOM}};
  ram_2_15 = _RAND_47[511:0];
  _RAND_48 = {16{`RANDOM}};
  ram_3_0 = _RAND_48[511:0];
  _RAND_49 = {16{`RANDOM}};
  ram_3_1 = _RAND_49[511:0];
  _RAND_50 = {16{`RANDOM}};
  ram_3_2 = _RAND_50[511:0];
  _RAND_51 = {16{`RANDOM}};
  ram_3_3 = _RAND_51[511:0];
  _RAND_52 = {16{`RANDOM}};
  ram_3_4 = _RAND_52[511:0];
  _RAND_53 = {16{`RANDOM}};
  ram_3_5 = _RAND_53[511:0];
  _RAND_54 = {16{`RANDOM}};
  ram_3_6 = _RAND_54[511:0];
  _RAND_55 = {16{`RANDOM}};
  ram_3_7 = _RAND_55[511:0];
  _RAND_56 = {16{`RANDOM}};
  ram_3_8 = _RAND_56[511:0];
  _RAND_57 = {16{`RANDOM}};
  ram_3_9 = _RAND_57[511:0];
  _RAND_58 = {16{`RANDOM}};
  ram_3_10 = _RAND_58[511:0];
  _RAND_59 = {16{`RANDOM}};
  ram_3_11 = _RAND_59[511:0];
  _RAND_60 = {16{`RANDOM}};
  ram_3_12 = _RAND_60[511:0];
  _RAND_61 = {16{`RANDOM}};
  ram_3_13 = _RAND_61[511:0];
  _RAND_62 = {16{`RANDOM}};
  ram_3_14 = _RAND_62[511:0];
  _RAND_63 = {16{`RANDOM}};
  ram_3_15 = _RAND_63[511:0];
  _RAND_64 = {1{`RANDOM}};
  tag_0_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  tag_0_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  tag_0_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  tag_0_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  tag_0_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  tag_0_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  tag_0_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  tag_0_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  tag_0_8 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  tag_0_9 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  tag_0_10 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  tag_0_11 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  tag_0_12 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  tag_0_13 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  tag_0_14 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  tag_0_15 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  tag_1_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  tag_1_1 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  tag_1_2 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  tag_1_3 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  tag_1_4 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  tag_1_5 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  tag_1_6 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  tag_1_7 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  tag_1_8 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  tag_1_9 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  tag_1_10 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  tag_1_11 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  tag_1_12 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  tag_1_13 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  tag_1_14 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  tag_1_15 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  tag_2_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  tag_2_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  tag_2_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  tag_2_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  tag_2_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  tag_2_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  tag_2_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  tag_2_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  tag_2_8 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  tag_2_9 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  tag_2_10 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  tag_2_11 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  tag_2_12 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  tag_2_13 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  tag_2_14 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  tag_2_15 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  tag_3_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  tag_3_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  tag_3_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  tag_3_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  tag_3_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  tag_3_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  tag_3_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  tag_3_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  tag_3_8 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  tag_3_9 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  tag_3_10 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  tag_3_11 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  tag_3_12 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  tag_3_13 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  tag_3_14 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  tag_3_15 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_1_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_1_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_1_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_1_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_1_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_1_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_1_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_1_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_1_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_1_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_1_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_1_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_1_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_1_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_1_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_1_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_2_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_2_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_2_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_2_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_2_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_2_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_2_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_2_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_2_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_2_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_2_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_2_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_2_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_2_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_2_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_2_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_3_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_3_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_3_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_3_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_3_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_3_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_3_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_3_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_3_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_3_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_3_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_3_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_3_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_3_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_3_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_3_15 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  dirty_0_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  dirty_0_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dirty_0_2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  dirty_0_3 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  dirty_0_4 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  dirty_0_5 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  dirty_0_6 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  dirty_0_7 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dirty_0_8 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  dirty_0_9 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  dirty_0_10 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  dirty_0_11 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  dirty_0_12 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  dirty_0_13 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dirty_0_14 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  dirty_0_15 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  dirty_1_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  dirty_1_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  dirty_1_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  dirty_1_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dirty_1_4 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  dirty_1_5 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  dirty_1_6 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  dirty_1_7 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  dirty_1_8 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  dirty_1_9 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  dirty_1_10 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  dirty_1_11 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  dirty_1_12 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  dirty_1_13 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  dirty_1_14 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  dirty_1_15 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  dirty_2_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  dirty_2_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  dirty_2_2 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  dirty_2_3 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  dirty_2_4 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  dirty_2_5 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  dirty_2_6 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  dirty_2_7 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  dirty_2_8 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  dirty_2_9 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  dirty_2_10 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  dirty_2_11 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  dirty_2_12 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  dirty_2_13 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  dirty_2_14 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  dirty_2_15 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  dirty_3_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  dirty_3_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  dirty_3_2 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  dirty_3_3 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  dirty_3_4 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  dirty_3_5 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  dirty_3_6 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  dirty_3_7 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  dirty_3_8 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  dirty_3_9 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  dirty_3_10 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  dirty_3_11 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  dirty_3_12 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  dirty_3_13 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  dirty_3_14 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  dirty_3_15 = _RAND_255[0:0];
  _RAND_256 = {16{`RANDOM}};
  write_back_data = _RAND_256[511:0];
  _RAND_257 = {1{`RANDOM}};
  write_back_addr = _RAND_257[31:0];
  _RAND_258 = {2{`RANDOM}};
  receive_data_0 = _RAND_258[63:0];
  _RAND_259 = {2{`RANDOM}};
  receive_data_1 = _RAND_259[63:0];
  _RAND_260 = {2{`RANDOM}};
  receive_data_2 = _RAND_260[63:0];
  _RAND_261 = {2{`RANDOM}};
  receive_data_3 = _RAND_261[63:0];
  _RAND_262 = {2{`RANDOM}};
  receive_data_4 = _RAND_262[63:0];
  _RAND_263 = {2{`RANDOM}};
  receive_data_5 = _RAND_263[63:0];
  _RAND_264 = {2{`RANDOM}};
  receive_data_6 = _RAND_264[63:0];
  _RAND_265 = {2{`RANDOM}};
  receive_data_7 = _RAND_265[63:0];
  _RAND_266 = {1{`RANDOM}};
  receive_num = _RAND_266[2:0];
  _RAND_267 = {1{`RANDOM}};
  quene_0 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  quene_1 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  quene_2 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  quene_3 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  quene_4 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  quene_5 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  quene_6 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  quene_7 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  quene_8 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  quene_9 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  quene_10 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  quene_11 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  quene_12 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  quene_13 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  quene_14 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  quene_15 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  state = _RAND_283[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI(
  input         clock,
  input         reset,
  input  [31:0] io_axi_in_araddr,
  input  [7:0]  io_axi_in_arlen,
  input         io_axi_in_arvalid,
  input         io_axi_in_rready,
  input  [31:0] io_axi_in_awaddr,
  input  [7:0]  io_axi_in_awlen,
  input         io_axi_in_awvalid,
  input  [63:0] io_axi_in_wdata,
  input  [7:0]  io_axi_in_wstrb,
  input         io_axi_in_wvalid,
  input         io_axi_in_bready,
  output [63:0] io_axi_out_rdata,
  output        io_axi_out_rlast,
  output        io_axi_out_rvalid,
  output        io_axi_out_wready,
  output        io_axi_out_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] Mem_modle_Raddr; // @[AXI.scala 30:27]
  wire [63:0] Mem_modle_Rdata; // @[AXI.scala 30:27]
  wire [63:0] Mem_modle_Waddr; // @[AXI.scala 30:27]
  wire [63:0] Mem_modle_Wdata; // @[AXI.scala 30:27]
  wire [7:0] Mem_modle_Wmask; // @[AXI.scala 30:27]
  wire  Mem_modle_Write_en; // @[AXI.scala 30:27]
  wire  Mem_modle_Read_en; // @[AXI.scala 30:27]
  reg  axi_wready; // @[AXI.scala 14:29]
  reg  axi_bvalid; // @[AXI.scala 17:29]
  reg  axi_rvalid; // @[AXI.scala 21:29]
  reg [7:0] arlen; // @[AXI.scala 22:24]
  reg [7:0] awlen; // @[AXI.scala 23:24]
  reg [63:0] araddr; // @[AXI.scala 24:25]
  reg [63:0] awaddr; // @[AXI.scala 25:25]
  reg [2:0] state; // @[AXI.scala 28:24]
  wire  _GEN_4 = io_axi_in_arvalid | axi_rvalid; // @[AXI.scala 55:42 60:28 21:29]
  wire  _GEN_7 = io_axi_in_awvalid & io_axi_in_wvalid | axi_wready; // @[AXI.scala 43:56 46:28 14:29]
  wire [63:0] _awaddr_T_1 = awaddr + 64'h8; // @[AXI.scala 72:38]
  wire [7:0] _awlen_T_1 = awlen - 8'h1; // @[AXI.scala 73:36]
  wire [63:0] _GEN_14 = io_axi_in_wvalid & axi_wready ? _awaddr_T_1 : awaddr; // @[AXI.scala 25:25 71:60 72:28]
  wire [7:0] _GEN_15 = io_axi_in_wvalid & axi_wready ? _awlen_T_1 : awlen; // @[AXI.scala 23:24 71:60 73:27]
  wire  _GEN_18 = awlen == 8'h0 | axi_bvalid; // @[AXI.scala 64:30 68:28 17:29]
  wire  _T_7 = arlen == 8'h0; // @[AXI.scala 78:23]
  wire [2:0] _GEN_22 = io_axi_in_rready ? 3'h0 : state; // @[AXI.scala 28:24 79:39 80:27]
  wire  _GEN_24 = io_axi_in_rready ? 1'h0 : axi_rvalid; // @[AXI.scala 21:29 79:39 82:32]
  wire [63:0] _araddr_T_1 = araddr + 64'h8; // @[AXI.scala 86:38]
  wire [7:0] _arlen_T_1 = arlen - 8'h1; // @[AXI.scala 87:36]
  wire [63:0] _GEN_25 = io_axi_in_rready ? _araddr_T_1 : araddr; // @[AXI.scala 24:25 85:39 86:28]
  wire [7:0] _GEN_26 = io_axi_in_rready ? _arlen_T_1 : arlen; // @[AXI.scala 22:24 85:39 87:27]
  wire [2:0] _GEN_27 = arlen == 8'h0 ? _GEN_22 : state; // @[AXI.scala 28:24 78:30]
  wire  _GEN_29 = arlen == 8'h0 ? _GEN_24 : axi_rvalid; // @[AXI.scala 21:29 78:30]
  wire [63:0] _GEN_30 = arlen == 8'h0 ? araddr : _GEN_25; // @[AXI.scala 24:25 78:30]
  wire [7:0] _GEN_31 = arlen == 8'h0 ? arlen : _GEN_26; // @[AXI.scala 22:24 78:30]
  wire [2:0] _GEN_32 = io_axi_in_bready ? 3'h0 : state; // @[AXI.scala 92:35 93:23 28:24]
  wire  _GEN_33 = io_axi_in_bready ? 1'h0 : axi_bvalid; // @[AXI.scala 92:35 94:28 17:29]
  wire [2:0] _GEN_35 = 3'h3 == state ? _GEN_32 : state; // @[AXI.scala 41:18 28:24]
  wire  _GEN_36 = 3'h3 == state ? _GEN_33 : axi_bvalid; // @[AXI.scala 41:18 17:29]
  MEM Mem_modle ( // @[AXI.scala 30:27]
    .Raddr(Mem_modle_Raddr),
    .Rdata(Mem_modle_Rdata),
    .Waddr(Mem_modle_Waddr),
    .Wdata(Mem_modle_Wdata),
    .Wmask(Mem_modle_Wmask),
    .Write_en(Mem_modle_Write_en),
    .Read_en(Mem_modle_Read_en)
  );
  assign io_axi_out_rdata = Mem_modle_Rdata; // @[AXI.scala 108:22]
  assign io_axi_out_rlast = state == 3'h1 & _T_7; // @[AXI.scala 110:41]
  assign io_axi_out_rvalid = axi_rvalid; // @[AXI.scala 109:23]
  assign io_axi_out_wready = axi_wready; // @[AXI.scala 112:23]
  assign io_axi_out_bvalid = axi_bvalid; // @[AXI.scala 113:23]
  assign Mem_modle_Raddr = araddr; // @[AXI.scala 31:24]
  assign Mem_modle_Waddr = awaddr; // @[AXI.scala 32:24]
  assign Mem_modle_Wdata = io_axi_in_wdata; // @[AXI.scala 33:24]
  assign Mem_modle_Wmask = io_axi_in_wstrb; // @[AXI.scala 34:24]
  assign Mem_modle_Write_en = axi_wready; // @[AXI.scala 35:27]
  assign Mem_modle_Read_en = axi_rvalid; // @[AXI.scala 36:26]
  always @(posedge clock) begin
    if (reset) begin // @[AXI.scala 14:29]
      axi_wready <= 1'h0; // @[AXI.scala 14:29]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      axi_wready <= _GEN_7;
    end else if (3'h2 == state) begin // @[AXI.scala 41:18]
      if (awlen == 8'h0) begin // @[AXI.scala 64:30]
        axi_wready <= 1'h0; // @[AXI.scala 65:28]
      end
    end
    if (reset) begin // @[AXI.scala 17:29]
      axi_bvalid <= 1'h0; // @[AXI.scala 17:29]
    end else if (!(3'h0 == state)) begin // @[AXI.scala 41:18]
      if (3'h2 == state) begin // @[AXI.scala 41:18]
        axi_bvalid <= _GEN_18;
      end else if (!(3'h1 == state)) begin // @[AXI.scala 41:18]
        axi_bvalid <= _GEN_36;
      end
    end
    if (reset) begin // @[AXI.scala 21:29]
      axi_rvalid <= 1'h0; // @[AXI.scala 21:29]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 43:56]
        axi_rvalid <= _GEN_4;
      end
    end else if (!(3'h2 == state)) begin // @[AXI.scala 41:18]
      if (3'h1 == state) begin // @[AXI.scala 41:18]
        axi_rvalid <= _GEN_29;
      end
    end
    if (reset) begin // @[AXI.scala 22:24]
      arlen <= 8'h0; // @[AXI.scala 22:24]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 43:56]
        if (io_axi_in_arvalid) begin // @[AXI.scala 55:42]
          arlen <= io_axi_in_arlen; // @[AXI.scala 57:23]
        end
      end
    end else if (!(3'h2 == state)) begin // @[AXI.scala 41:18]
      if (3'h1 == state) begin // @[AXI.scala 41:18]
        arlen <= _GEN_31;
      end
    end
    if (reset) begin // @[AXI.scala 23:24]
      awlen <= 8'h0; // @[AXI.scala 23:24]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 43:56]
        awlen <= io_axi_in_awlen; // @[AXI.scala 48:23]
      end
    end else if (3'h2 == state) begin // @[AXI.scala 41:18]
      if (!(awlen == 8'h0)) begin // @[AXI.scala 64:30]
        awlen <= _GEN_15;
      end
    end
    if (reset) begin // @[AXI.scala 24:25]
      araddr <= 64'h0; // @[AXI.scala 24:25]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 43:56]
        if (io_axi_in_arvalid) begin // @[AXI.scala 55:42]
          araddr <= {{32'd0}, io_axi_in_araddr}; // @[AXI.scala 58:24]
        end
      end
    end else if (!(3'h2 == state)) begin // @[AXI.scala 41:18]
      if (3'h1 == state) begin // @[AXI.scala 41:18]
        araddr <= _GEN_30;
      end
    end
    if (reset) begin // @[AXI.scala 25:25]
      awaddr <= 64'h0; // @[AXI.scala 25:25]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 43:56]
        awaddr <= {{32'd0}, io_axi_in_awaddr}; // @[AXI.scala 49:24]
      end
    end else if (3'h2 == state) begin // @[AXI.scala 41:18]
      if (!(awlen == 8'h0)) begin // @[AXI.scala 64:30]
        awaddr <= _GEN_14;
      end
    end
    if (reset) begin // @[AXI.scala 28:24]
      state <= 3'h0; // @[AXI.scala 28:24]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 43:56]
        state <= 3'h2; // @[AXI.scala 44:23]
      end else if (io_axi_in_arvalid) begin // @[AXI.scala 55:42]
        state <= 3'h1; // @[AXI.scala 56:23]
      end
    end else if (3'h2 == state) begin // @[AXI.scala 41:18]
      if (awlen == 8'h0) begin // @[AXI.scala 64:30]
        state <= 3'h3; // @[AXI.scala 69:23]
      end
    end else if (3'h1 == state) begin // @[AXI.scala 41:18]
      state <= _GEN_27;
    end else begin
      state <= _GEN_35;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_wready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_bvalid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_rvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  arlen = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  awlen = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  araddr = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  awaddr = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input         clock,
  input         reset,
  output [31:0] io_inst,
  output [63:0] io_pc,
  output        io_step
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  Register_clock; // @[top.scala 15:25]
  wire [4:0] Register_io_raddr1; // @[top.scala 15:25]
  wire [4:0] Register_io_raddr2; // @[top.scala 15:25]
  wire [63:0] Register_io_rdata1; // @[top.scala 15:25]
  wire [63:0] Register_io_rdata2; // @[top.scala 15:25]
  wire  Register_io_we; // @[top.scala 15:25]
  wire [4:0] Register_io_waddr; // @[top.scala 15:25]
  wire [63:0] Register_io_wdata; // @[top.scala 15:25]
  wire  IFU_clock; // @[top.scala 16:21]
  wire  IFU_reset; // @[top.scala 16:21]
  wire  IFU_io_ds_allowin; // @[top.scala 16:21]
  wire  IFU_io_br_taken; // @[top.scala 16:21]
  wire [63:0] IFU_io_br_target; // @[top.scala 16:21]
  wire [63:0] IFU_io_to_ds_pc; // @[top.scala 16:21]
  wire  IFU_io_fs_to_ds_valid; // @[top.scala 16:21]
  wire [31:0] IFU_io_inst; // @[top.scala 16:21]
  wire [63:0] IFU_io_axi_in_rdata; // @[top.scala 16:21]
  wire  IFU_io_axi_in_rlast; // @[top.scala 16:21]
  wire  IFU_io_axi_in_rvalid; // @[top.scala 16:21]
  wire [31:0] IFU_io_axi_out_araddr; // @[top.scala 16:21]
  wire  IFU_io_axi_out_arvalid; // @[top.scala 16:21]
  wire  IFU_io_axi_out_rready; // @[top.scala 16:21]
  wire  IFU_io_fence; // @[top.scala 16:21]
  wire  IFU_io_clear_cache; // @[top.scala 16:21]
  wire  IFU_io_cache_init; // @[top.scala 16:21]
  wire  IDU_clock; // @[top.scala 17:21]
  wire  IDU_reset; // @[top.scala 17:21]
  wire [63:0] IDU_io_pc; // @[top.scala 17:21]
  wire  IDU_io_fs_to_ds_valid; // @[top.scala 17:21]
  wire  IDU_io_ds_to_es_valid; // @[top.scala 17:21]
  wire  IDU_io_es_allowin; // @[top.scala 17:21]
  wire [31:0] IDU_io_from_fs_inst; // @[top.scala 17:21]
  wire  IDU_io_br_taken; // @[top.scala 17:21]
  wire [63:0] IDU_io_br_target; // @[top.scala 17:21]
  wire  IDU_io_ds_allowin; // @[top.scala 17:21]
  wire  IDU_io_fence; // @[top.scala 17:21]
  wire [4:0] IDU_io_raddr1; // @[top.scala 17:21]
  wire [4:0] IDU_io_raddr2; // @[top.scala 17:21]
  wire [63:0] IDU_io_rdata1; // @[top.scala 17:21]
  wire [63:0] IDU_io_rdata2; // @[top.scala 17:21]
  wire [63:0] IDU_io_to_es_pc; // @[top.scala 17:21]
  wire [31:0] IDU_io_ALUop; // @[top.scala 17:21]
  wire [63:0] IDU_io_src1; // @[top.scala 17:21]
  wire [63:0] IDU_io_src2; // @[top.scala 17:21]
  wire [4:0] IDU_io_rf_dst; // @[top.scala 17:21]
  wire [63:0] IDU_io_store_data; // @[top.scala 17:21]
  wire  IDU_io_ctrl_sign_reg_write; // @[top.scala 17:21]
  wire  IDU_io_ctrl_sign_Writemem_en; // @[top.scala 17:21]
  wire  IDU_io_ctrl_sign_Readmem_en; // @[top.scala 17:21]
  wire [7:0] IDU_io_ctrl_sign_Wmask; // @[top.scala 17:21]
  wire [2:0] IDU_io_load_type; // @[top.scala 17:21]
  wire  IDU_io_es_ld; // @[top.scala 17:21]
  wire [63:0] IDU_io_es_fwd_res; // @[top.scala 17:21]
  wire [63:0] IDU_io_ms_fwd_res; // @[top.scala 17:21]
  wire [63:0] IDU_io_ws_fwd_res; // @[top.scala 17:21]
  wire  IDU_io_es_fwd_ready; // @[top.scala 17:21]
  wire  IDU_io_ms_fwd_ready; // @[top.scala 17:21]
  wire  IDU_io_es_rf_we; // @[top.scala 17:21]
  wire  IDU_io_ms_rf_we; // @[top.scala 17:21]
  wire  IDU_io_ws_rf_we; // @[top.scala 17:21]
  wire  IDU_io_es_valid; // @[top.scala 17:21]
  wire  IDU_io_ms_valid; // @[top.scala 17:21]
  wire  IDU_io_ws_valid; // @[top.scala 17:21]
  wire [4:0] IDU_io_es_rf_dst; // @[top.scala 17:21]
  wire [4:0] IDU_io_ms_rf_dst; // @[top.scala 17:21]
  wire [4:0] IDU_io_ws_rf_dst; // @[top.scala 17:21]
  wire  IDU_io_ds_valid; // @[top.scala 17:21]
  wire  EXU_clock; // @[top.scala 18:21]
  wire  EXU_reset; // @[top.scala 18:21]
  wire [63:0] EXU_io_pc; // @[top.scala 18:21]
  wire  EXU_io_ds_to_es_valid; // @[top.scala 18:21]
  wire  EXU_io_ms_allowin; // @[top.scala 18:21]
  wire  EXU_io_es_allowin; // @[top.scala 18:21]
  wire [31:0] EXU_io_ALUop; // @[top.scala 18:21]
  wire [63:0] EXU_io_src1_value; // @[top.scala 18:21]
  wire [63:0] EXU_io_src2_value; // @[top.scala 18:21]
  wire [4:0] EXU_io_rf_dst; // @[top.scala 18:21]
  wire [63:0] EXU_io_store_data; // @[top.scala 18:21]
  wire  EXU_io_es_to_ms_valid; // @[top.scala 18:21]
  wire [2:0] EXU_io_load_type; // @[top.scala 18:21]
  wire [63:0] EXU_io_to_ms_pc; // @[top.scala 18:21]
  wire [63:0] EXU_io_to_ms_alures; // @[top.scala 18:21]
  wire [63:0] EXU_io_to_ms_store_data; // @[top.scala 18:21]
  wire  EXU_io_to_ms_wen; // @[top.scala 18:21]
  wire [7:0] EXU_io_to_ms_wstrb; // @[top.scala 18:21]
  wire  EXU_io_to_ms_ren; // @[top.scala 18:21]
  wire [63:0] EXU_io_to_ms_maddr; // @[top.scala 18:21]
  wire [4:0] EXU_io_to_ms_rf_dst; // @[top.scala 18:21]
  wire  EXU_io_to_ms_rf_we; // @[top.scala 18:21]
  wire [2:0] EXU_io_to_ms_load_type; // @[top.scala 18:21]
  wire  EXU_io_ctrl_sign_reg_write; // @[top.scala 18:21]
  wire  EXU_io_ctrl_sign_Writemem_en; // @[top.scala 18:21]
  wire  EXU_io_ctrl_sign_Readmem_en; // @[top.scala 18:21]
  wire [7:0] EXU_io_ctrl_sign_Wmask; // @[top.scala 18:21]
  wire  EXU_io_es_valid; // @[top.scala 18:21]
  wire  EXU_io_es_rf_we; // @[top.scala 18:21]
  wire [4:0] EXU_io_es_rf_dst; // @[top.scala 18:21]
  wire  EXU_io_es_fwd_ready; // @[top.scala 18:21]
  wire [63:0] EXU_io_es_fwd_res; // @[top.scala 18:21]
  wire  EXU_io_es_ld; // @[top.scala 18:21]
  wire  LSU_clock; // @[top.scala 19:21]
  wire  LSU_reset; // @[top.scala 19:21]
  wire [63:0] LSU_io_pc; // @[top.scala 19:21]
  wire  LSU_io_es_to_ms_valid; // @[top.scala 19:21]
  wire  LSU_io_ms_allowin; // @[top.scala 19:21]
  wire  LSU_io_rf_we; // @[top.scala 19:21]
  wire [4:0] LSU_io_rf_dst; // @[top.scala 19:21]
  wire [63:0] LSU_io_alu_res; // @[top.scala 19:21]
  wire [63:0] LSU_io_store_data; // @[top.scala 19:21]
  wire [2:0] LSU_io_load_type; // @[top.scala 19:21]
  wire  LSU_io_wen; // @[top.scala 19:21]
  wire [7:0] LSU_io_wstrb; // @[top.scala 19:21]
  wire  LSU_io_ren; // @[top.scala 19:21]
  wire [63:0] LSU_io_maddr; // @[top.scala 19:21]
  wire [63:0] LSU_io_to_ws_pc; // @[top.scala 19:21]
  wire [63:0] LSU_io_ms_final_res; // @[top.scala 19:21]
  wire  LSU_io_ms_to_ws_valid; // @[top.scala 19:21]
  wire  LSU_io_to_ws_rf_we; // @[top.scala 19:21]
  wire [4:0] LSU_io_to_ws_rf_dst; // @[top.scala 19:21]
  wire  LSU_io_ms_valid; // @[top.scala 19:21]
  wire  LSU_io_ms_rf_we; // @[top.scala 19:21]
  wire [4:0] LSU_io_ms_rf_dst; // @[top.scala 19:21]
  wire  LSU_io_ms_fwd_ready; // @[top.scala 19:21]
  wire [63:0] LSU_io_ms_fwd_res; // @[top.scala 19:21]
  wire [63:0] LSU_io_axi_in_rdata; // @[top.scala 19:21]
  wire  LSU_io_axi_in_rvalid; // @[top.scala 19:21]
  wire  LSU_io_axi_in_wready; // @[top.scala 19:21]
  wire [31:0] LSU_io_axi_out_araddr; // @[top.scala 19:21]
  wire  LSU_io_axi_out_arvalid; // @[top.scala 19:21]
  wire [31:0] LSU_io_axi_out_awaddr; // @[top.scala 19:21]
  wire  LSU_io_axi_out_awvalid; // @[top.scala 19:21]
  wire [63:0] LSU_io_axi_out_wdata; // @[top.scala 19:21]
  wire [7:0] LSU_io_axi_out_wstrb; // @[top.scala 19:21]
  wire  LSU_io_axi_out_wvalid; // @[top.scala 19:21]
  wire  WBU_clock; // @[top.scala 20:21]
  wire  WBU_reset; // @[top.scala 20:21]
  wire [63:0] WBU_io_pc; // @[top.scala 20:21]
  wire  WBU_io_ms_to_ws_valid; // @[top.scala 20:21]
  wire [63:0] WBU_io_ms_final_res; // @[top.scala 20:21]
  wire  WBU_io_rf_we; // @[top.scala 20:21]
  wire [4:0] WBU_io_rf_dst; // @[top.scala 20:21]
  wire  WBU_io_we; // @[top.scala 20:21]
  wire [4:0] WBU_io_waddr; // @[top.scala 20:21]
  wire [63:0] WBU_io_wdata; // @[top.scala 20:21]
  wire  WBU_io_ws_valid; // @[top.scala 20:21]
  wire  WBU_io_ws_rf_we; // @[top.scala 20:21]
  wire [4:0] WBU_io_ws_rf_dst; // @[top.scala 20:21]
  wire [63:0] WBU_io_ws_fwd_res; // @[top.scala 20:21]
  wire [63:0] WBU_io_ws_pc; // @[top.scala 20:21]
  wire  arbiter_clock; // @[top.scala 21:25]
  wire  arbiter_reset; // @[top.scala 21:25]
  wire [31:0] arbiter_io_ifu_axi_in_araddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_ifu_axi_in_arlen; // @[top.scala 21:25]
  wire  arbiter_io_ifu_axi_in_arvalid; // @[top.scala 21:25]
  wire  arbiter_io_ifu_axi_in_rready; // @[top.scala 21:25]
  wire [63:0] arbiter_io_ifu_axi_out_rdata; // @[top.scala 21:25]
  wire  arbiter_io_ifu_axi_out_rlast; // @[top.scala 21:25]
  wire  arbiter_io_ifu_axi_out_rvalid; // @[top.scala 21:25]
  wire [31:0] arbiter_io_lsu_axi_in_araddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_lsu_axi_in_arlen; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_arvalid; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_rready; // @[top.scala 21:25]
  wire [31:0] arbiter_io_lsu_axi_in_awaddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_lsu_axi_in_awlen; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_awvalid; // @[top.scala 21:25]
  wire [63:0] arbiter_io_lsu_axi_in_wdata; // @[top.scala 21:25]
  wire [7:0] arbiter_io_lsu_axi_in_wstrb; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_wvalid; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_bready; // @[top.scala 21:25]
  wire [63:0] arbiter_io_lsu_axi_out_rdata; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_out_rlast; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_out_rvalid; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_out_wready; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_out_bvalid; // @[top.scala 21:25]
  wire [63:0] arbiter_io_axi_in_rdata; // @[top.scala 21:25]
  wire  arbiter_io_axi_in_rlast; // @[top.scala 21:25]
  wire  arbiter_io_axi_in_rvalid; // @[top.scala 21:25]
  wire  arbiter_io_axi_in_wready; // @[top.scala 21:25]
  wire  arbiter_io_axi_in_bvalid; // @[top.scala 21:25]
  wire [31:0] arbiter_io_axi_out_araddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_axi_out_arlen; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_arvalid; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_rready; // @[top.scala 21:25]
  wire [31:0] arbiter_io_axi_out_awaddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_axi_out_awlen; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_awvalid; // @[top.scala 21:25]
  wire [63:0] arbiter_io_axi_out_wdata; // @[top.scala 21:25]
  wire [7:0] arbiter_io_axi_out_wstrb; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_wvalid; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_bready; // @[top.scala 21:25]
  wire  i_cache_clock; // @[top.scala 22:25]
  wire  i_cache_reset; // @[top.scala 22:25]
  wire [31:0] i_cache_io_from_ifu_araddr; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_rready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_to_ifu_rdata; // @[top.scala 22:25]
  wire  i_cache_io_to_ifu_rlast; // @[top.scala 22:25]
  wire  i_cache_io_to_ifu_rvalid; // @[top.scala 22:25]
  wire [31:0] i_cache_io_to_axi_araddr; // @[top.scala 22:25]
  wire [7:0] i_cache_io_to_axi_arlen; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_rready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_from_axi_rdata; // @[top.scala 22:25]
  wire  i_cache_io_from_axi_rlast; // @[top.scala 22:25]
  wire  i_cache_io_from_axi_rvalid; // @[top.scala 22:25]
  wire  i_cache_io_cache_init; // @[top.scala 22:25]
  wire  i_cache_io_clear_cache; // @[top.scala 22:25]
  wire  d_cache_clock; // @[top.scala 23:25]
  wire  d_cache_reset; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_araddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_arvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_awaddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_awvalid; // @[top.scala 23:25]
  wire [63:0] d_cache_io_from_lsu_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_from_lsu_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_wvalid; // @[top.scala 23:25]
  wire [63:0] d_cache_io_to_lsu_rdata; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_wready; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_araddr; // @[top.scala 23:25]
  wire [7:0] d_cache_io_to_axi_arlen; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_arvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_rready; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_awaddr; // @[top.scala 23:25]
  wire [7:0] d_cache_io_to_axi_awlen; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_awvalid; // @[top.scala 23:25]
  wire [63:0] d_cache_io_to_axi_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_to_axi_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_wvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_bready; // @[top.scala 23:25]
  wire [63:0] d_cache_io_from_axi_rdata; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_rlast; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_wready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_bvalid; // @[top.scala 23:25]
  wire  axi_clock; // @[top.scala 24:21]
  wire  axi_reset; // @[top.scala 24:21]
  wire [31:0] axi_io_axi_in_araddr; // @[top.scala 24:21]
  wire [7:0] axi_io_axi_in_arlen; // @[top.scala 24:21]
  wire  axi_io_axi_in_arvalid; // @[top.scala 24:21]
  wire  axi_io_axi_in_rready; // @[top.scala 24:21]
  wire [31:0] axi_io_axi_in_awaddr; // @[top.scala 24:21]
  wire [7:0] axi_io_axi_in_awlen; // @[top.scala 24:21]
  wire  axi_io_axi_in_awvalid; // @[top.scala 24:21]
  wire [63:0] axi_io_axi_in_wdata; // @[top.scala 24:21]
  wire [7:0] axi_io_axi_in_wstrb; // @[top.scala 24:21]
  wire  axi_io_axi_in_wvalid; // @[top.scala 24:21]
  wire  axi_io_axi_in_bready; // @[top.scala 24:21]
  wire [63:0] axi_io_axi_out_rdata; // @[top.scala 24:21]
  wire  axi_io_axi_out_rlast; // @[top.scala 24:21]
  wire  axi_io_axi_out_rvalid; // @[top.scala 24:21]
  wire  axi_io_axi_out_wready; // @[top.scala 24:21]
  wire  axi_io_axi_out_bvalid; // @[top.scala 24:21]
  wire [31:0] dpi_flag; // @[top.scala 114:21]
  wire [31:0] dpi_ecall_flag; // @[top.scala 114:21]
  wire [63:0] dpi_pc; // @[top.scala 114:21]
  reg  diff_step; // @[top.scala 111:28]
  wire [63:0] _dpi_io_pc_T = IDU_io_ds_valid ? EXU_io_pc : IDU_io_pc; // @[top.scala 117:96]
  wire [63:0] _dpi_io_pc_T_1 = EXU_io_es_valid ? LSU_io_pc : _dpi_io_pc_T; // @[top.scala 117:72]
  wire [63:0] _dpi_io_pc_T_2 = LSU_io_ms_valid ? WBU_io_pc : _dpi_io_pc_T_1; // @[top.scala 117:48]
  Register Register ( // @[top.scala 15:25]
    .clock(Register_clock),
    .io_raddr1(Register_io_raddr1),
    .io_raddr2(Register_io_raddr2),
    .io_rdata1(Register_io_rdata1),
    .io_rdata2(Register_io_rdata2),
    .io_we(Register_io_we),
    .io_waddr(Register_io_waddr),
    .io_wdata(Register_io_wdata)
  );
  IFU IFU ( // @[top.scala 16:21]
    .clock(IFU_clock),
    .reset(IFU_reset),
    .io_ds_allowin(IFU_io_ds_allowin),
    .io_br_taken(IFU_io_br_taken),
    .io_br_target(IFU_io_br_target),
    .io_to_ds_pc(IFU_io_to_ds_pc),
    .io_fs_to_ds_valid(IFU_io_fs_to_ds_valid),
    .io_inst(IFU_io_inst),
    .io_axi_in_rdata(IFU_io_axi_in_rdata),
    .io_axi_in_rlast(IFU_io_axi_in_rlast),
    .io_axi_in_rvalid(IFU_io_axi_in_rvalid),
    .io_axi_out_araddr(IFU_io_axi_out_araddr),
    .io_axi_out_arvalid(IFU_io_axi_out_arvalid),
    .io_axi_out_rready(IFU_io_axi_out_rready),
    .io_fence(IFU_io_fence),
    .io_clear_cache(IFU_io_clear_cache),
    .io_cache_init(IFU_io_cache_init)
  );
  IDU IDU ( // @[top.scala 17:21]
    .clock(IDU_clock),
    .reset(IDU_reset),
    .io_pc(IDU_io_pc),
    .io_fs_to_ds_valid(IDU_io_fs_to_ds_valid),
    .io_ds_to_es_valid(IDU_io_ds_to_es_valid),
    .io_es_allowin(IDU_io_es_allowin),
    .io_from_fs_inst(IDU_io_from_fs_inst),
    .io_br_taken(IDU_io_br_taken),
    .io_br_target(IDU_io_br_target),
    .io_ds_allowin(IDU_io_ds_allowin),
    .io_fence(IDU_io_fence),
    .io_raddr1(IDU_io_raddr1),
    .io_raddr2(IDU_io_raddr2),
    .io_rdata1(IDU_io_rdata1),
    .io_rdata2(IDU_io_rdata2),
    .io_to_es_pc(IDU_io_to_es_pc),
    .io_ALUop(IDU_io_ALUop),
    .io_src1(IDU_io_src1),
    .io_src2(IDU_io_src2),
    .io_rf_dst(IDU_io_rf_dst),
    .io_store_data(IDU_io_store_data),
    .io_ctrl_sign_reg_write(IDU_io_ctrl_sign_reg_write),
    .io_ctrl_sign_Writemem_en(IDU_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(IDU_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(IDU_io_ctrl_sign_Wmask),
    .io_load_type(IDU_io_load_type),
    .io_es_ld(IDU_io_es_ld),
    .io_es_fwd_res(IDU_io_es_fwd_res),
    .io_ms_fwd_res(IDU_io_ms_fwd_res),
    .io_ws_fwd_res(IDU_io_ws_fwd_res),
    .io_es_fwd_ready(IDU_io_es_fwd_ready),
    .io_ms_fwd_ready(IDU_io_ms_fwd_ready),
    .io_es_rf_we(IDU_io_es_rf_we),
    .io_ms_rf_we(IDU_io_ms_rf_we),
    .io_ws_rf_we(IDU_io_ws_rf_we),
    .io_es_valid(IDU_io_es_valid),
    .io_ms_valid(IDU_io_ms_valid),
    .io_ws_valid(IDU_io_ws_valid),
    .io_es_rf_dst(IDU_io_es_rf_dst),
    .io_ms_rf_dst(IDU_io_ms_rf_dst),
    .io_ws_rf_dst(IDU_io_ws_rf_dst),
    .io_ds_valid(IDU_io_ds_valid)
  );
  EXU EXU ( // @[top.scala 18:21]
    .clock(EXU_clock),
    .reset(EXU_reset),
    .io_pc(EXU_io_pc),
    .io_ds_to_es_valid(EXU_io_ds_to_es_valid),
    .io_ms_allowin(EXU_io_ms_allowin),
    .io_es_allowin(EXU_io_es_allowin),
    .io_ALUop(EXU_io_ALUop),
    .io_src1_value(EXU_io_src1_value),
    .io_src2_value(EXU_io_src2_value),
    .io_rf_dst(EXU_io_rf_dst),
    .io_store_data(EXU_io_store_data),
    .io_es_to_ms_valid(EXU_io_es_to_ms_valid),
    .io_load_type(EXU_io_load_type),
    .io_to_ms_pc(EXU_io_to_ms_pc),
    .io_to_ms_alures(EXU_io_to_ms_alures),
    .io_to_ms_store_data(EXU_io_to_ms_store_data),
    .io_to_ms_wen(EXU_io_to_ms_wen),
    .io_to_ms_wstrb(EXU_io_to_ms_wstrb),
    .io_to_ms_ren(EXU_io_to_ms_ren),
    .io_to_ms_maddr(EXU_io_to_ms_maddr),
    .io_to_ms_rf_dst(EXU_io_to_ms_rf_dst),
    .io_to_ms_rf_we(EXU_io_to_ms_rf_we),
    .io_to_ms_load_type(EXU_io_to_ms_load_type),
    .io_ctrl_sign_reg_write(EXU_io_ctrl_sign_reg_write),
    .io_ctrl_sign_Writemem_en(EXU_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(EXU_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(EXU_io_ctrl_sign_Wmask),
    .io_es_valid(EXU_io_es_valid),
    .io_es_rf_we(EXU_io_es_rf_we),
    .io_es_rf_dst(EXU_io_es_rf_dst),
    .io_es_fwd_ready(EXU_io_es_fwd_ready),
    .io_es_fwd_res(EXU_io_es_fwd_res),
    .io_es_ld(EXU_io_es_ld)
  );
  LSU LSU ( // @[top.scala 19:21]
    .clock(LSU_clock),
    .reset(LSU_reset),
    .io_pc(LSU_io_pc),
    .io_es_to_ms_valid(LSU_io_es_to_ms_valid),
    .io_ms_allowin(LSU_io_ms_allowin),
    .io_rf_we(LSU_io_rf_we),
    .io_rf_dst(LSU_io_rf_dst),
    .io_alu_res(LSU_io_alu_res),
    .io_store_data(LSU_io_store_data),
    .io_load_type(LSU_io_load_type),
    .io_wen(LSU_io_wen),
    .io_wstrb(LSU_io_wstrb),
    .io_ren(LSU_io_ren),
    .io_maddr(LSU_io_maddr),
    .io_to_ws_pc(LSU_io_to_ws_pc),
    .io_ms_final_res(LSU_io_ms_final_res),
    .io_ms_to_ws_valid(LSU_io_ms_to_ws_valid),
    .io_to_ws_rf_we(LSU_io_to_ws_rf_we),
    .io_to_ws_rf_dst(LSU_io_to_ws_rf_dst),
    .io_ms_valid(LSU_io_ms_valid),
    .io_ms_rf_we(LSU_io_ms_rf_we),
    .io_ms_rf_dst(LSU_io_ms_rf_dst),
    .io_ms_fwd_ready(LSU_io_ms_fwd_ready),
    .io_ms_fwd_res(LSU_io_ms_fwd_res),
    .io_axi_in_rdata(LSU_io_axi_in_rdata),
    .io_axi_in_rvalid(LSU_io_axi_in_rvalid),
    .io_axi_in_wready(LSU_io_axi_in_wready),
    .io_axi_out_araddr(LSU_io_axi_out_araddr),
    .io_axi_out_arvalid(LSU_io_axi_out_arvalid),
    .io_axi_out_awaddr(LSU_io_axi_out_awaddr),
    .io_axi_out_awvalid(LSU_io_axi_out_awvalid),
    .io_axi_out_wdata(LSU_io_axi_out_wdata),
    .io_axi_out_wstrb(LSU_io_axi_out_wstrb),
    .io_axi_out_wvalid(LSU_io_axi_out_wvalid)
  );
  WBU WBU ( // @[top.scala 20:21]
    .clock(WBU_clock),
    .reset(WBU_reset),
    .io_pc(WBU_io_pc),
    .io_ms_to_ws_valid(WBU_io_ms_to_ws_valid),
    .io_ms_final_res(WBU_io_ms_final_res),
    .io_rf_we(WBU_io_rf_we),
    .io_rf_dst(WBU_io_rf_dst),
    .io_we(WBU_io_we),
    .io_waddr(WBU_io_waddr),
    .io_wdata(WBU_io_wdata),
    .io_ws_valid(WBU_io_ws_valid),
    .io_ws_rf_we(WBU_io_ws_rf_we),
    .io_ws_rf_dst(WBU_io_ws_rf_dst),
    .io_ws_fwd_res(WBU_io_ws_fwd_res),
    .io_ws_pc(WBU_io_ws_pc)
  );
  AXI_ARBITER arbiter ( // @[top.scala 21:25]
    .clock(arbiter_clock),
    .reset(arbiter_reset),
    .io_ifu_axi_in_araddr(arbiter_io_ifu_axi_in_araddr),
    .io_ifu_axi_in_arlen(arbiter_io_ifu_axi_in_arlen),
    .io_ifu_axi_in_arvalid(arbiter_io_ifu_axi_in_arvalid),
    .io_ifu_axi_in_rready(arbiter_io_ifu_axi_in_rready),
    .io_ifu_axi_out_rdata(arbiter_io_ifu_axi_out_rdata),
    .io_ifu_axi_out_rlast(arbiter_io_ifu_axi_out_rlast),
    .io_ifu_axi_out_rvalid(arbiter_io_ifu_axi_out_rvalid),
    .io_lsu_axi_in_araddr(arbiter_io_lsu_axi_in_araddr),
    .io_lsu_axi_in_arlen(arbiter_io_lsu_axi_in_arlen),
    .io_lsu_axi_in_arvalid(arbiter_io_lsu_axi_in_arvalid),
    .io_lsu_axi_in_rready(arbiter_io_lsu_axi_in_rready),
    .io_lsu_axi_in_awaddr(arbiter_io_lsu_axi_in_awaddr),
    .io_lsu_axi_in_awlen(arbiter_io_lsu_axi_in_awlen),
    .io_lsu_axi_in_awvalid(arbiter_io_lsu_axi_in_awvalid),
    .io_lsu_axi_in_wdata(arbiter_io_lsu_axi_in_wdata),
    .io_lsu_axi_in_wstrb(arbiter_io_lsu_axi_in_wstrb),
    .io_lsu_axi_in_wvalid(arbiter_io_lsu_axi_in_wvalid),
    .io_lsu_axi_in_bready(arbiter_io_lsu_axi_in_bready),
    .io_lsu_axi_out_rdata(arbiter_io_lsu_axi_out_rdata),
    .io_lsu_axi_out_rlast(arbiter_io_lsu_axi_out_rlast),
    .io_lsu_axi_out_rvalid(arbiter_io_lsu_axi_out_rvalid),
    .io_lsu_axi_out_wready(arbiter_io_lsu_axi_out_wready),
    .io_lsu_axi_out_bvalid(arbiter_io_lsu_axi_out_bvalid),
    .io_axi_in_rdata(arbiter_io_axi_in_rdata),
    .io_axi_in_rlast(arbiter_io_axi_in_rlast),
    .io_axi_in_rvalid(arbiter_io_axi_in_rvalid),
    .io_axi_in_wready(arbiter_io_axi_in_wready),
    .io_axi_in_bvalid(arbiter_io_axi_in_bvalid),
    .io_axi_out_araddr(arbiter_io_axi_out_araddr),
    .io_axi_out_arlen(arbiter_io_axi_out_arlen),
    .io_axi_out_arvalid(arbiter_io_axi_out_arvalid),
    .io_axi_out_rready(arbiter_io_axi_out_rready),
    .io_axi_out_awaddr(arbiter_io_axi_out_awaddr),
    .io_axi_out_awlen(arbiter_io_axi_out_awlen),
    .io_axi_out_awvalid(arbiter_io_axi_out_awvalid),
    .io_axi_out_wdata(arbiter_io_axi_out_wdata),
    .io_axi_out_wstrb(arbiter_io_axi_out_wstrb),
    .io_axi_out_wvalid(arbiter_io_axi_out_wvalid),
    .io_axi_out_bready(arbiter_io_axi_out_bready)
  );
  I_CACHE i_cache ( // @[top.scala 22:25]
    .clock(i_cache_clock),
    .reset(i_cache_reset),
    .io_from_ifu_araddr(i_cache_io_from_ifu_araddr),
    .io_from_ifu_arvalid(i_cache_io_from_ifu_arvalid),
    .io_from_ifu_rready(i_cache_io_from_ifu_rready),
    .io_to_ifu_rdata(i_cache_io_to_ifu_rdata),
    .io_to_ifu_rlast(i_cache_io_to_ifu_rlast),
    .io_to_ifu_rvalid(i_cache_io_to_ifu_rvalid),
    .io_to_axi_araddr(i_cache_io_to_axi_araddr),
    .io_to_axi_arlen(i_cache_io_to_axi_arlen),
    .io_to_axi_arvalid(i_cache_io_to_axi_arvalid),
    .io_to_axi_rready(i_cache_io_to_axi_rready),
    .io_from_axi_rdata(i_cache_io_from_axi_rdata),
    .io_from_axi_rlast(i_cache_io_from_axi_rlast),
    .io_from_axi_rvalid(i_cache_io_from_axi_rvalid),
    .io_cache_init(i_cache_io_cache_init),
    .io_clear_cache(i_cache_io_clear_cache)
  );
  D_CACHE d_cache ( // @[top.scala 23:25]
    .clock(d_cache_clock),
    .reset(d_cache_reset),
    .io_from_lsu_araddr(d_cache_io_from_lsu_araddr),
    .io_from_lsu_arvalid(d_cache_io_from_lsu_arvalid),
    .io_from_lsu_awaddr(d_cache_io_from_lsu_awaddr),
    .io_from_lsu_awvalid(d_cache_io_from_lsu_awvalid),
    .io_from_lsu_wdata(d_cache_io_from_lsu_wdata),
    .io_from_lsu_wstrb(d_cache_io_from_lsu_wstrb),
    .io_from_lsu_wvalid(d_cache_io_from_lsu_wvalid),
    .io_to_lsu_rdata(d_cache_io_to_lsu_rdata),
    .io_to_lsu_rvalid(d_cache_io_to_lsu_rvalid),
    .io_to_lsu_wready(d_cache_io_to_lsu_wready),
    .io_to_axi_araddr(d_cache_io_to_axi_araddr),
    .io_to_axi_arlen(d_cache_io_to_axi_arlen),
    .io_to_axi_arvalid(d_cache_io_to_axi_arvalid),
    .io_to_axi_rready(d_cache_io_to_axi_rready),
    .io_to_axi_awaddr(d_cache_io_to_axi_awaddr),
    .io_to_axi_awlen(d_cache_io_to_axi_awlen),
    .io_to_axi_awvalid(d_cache_io_to_axi_awvalid),
    .io_to_axi_wdata(d_cache_io_to_axi_wdata),
    .io_to_axi_wstrb(d_cache_io_to_axi_wstrb),
    .io_to_axi_wvalid(d_cache_io_to_axi_wvalid),
    .io_to_axi_bready(d_cache_io_to_axi_bready),
    .io_from_axi_rdata(d_cache_io_from_axi_rdata),
    .io_from_axi_rlast(d_cache_io_from_axi_rlast),
    .io_from_axi_rvalid(d_cache_io_from_axi_rvalid),
    .io_from_axi_wready(d_cache_io_from_axi_wready),
    .io_from_axi_bvalid(d_cache_io_from_axi_bvalid)
  );
  AXI axi ( // @[top.scala 24:21]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_axi_in_araddr(axi_io_axi_in_araddr),
    .io_axi_in_arlen(axi_io_axi_in_arlen),
    .io_axi_in_arvalid(axi_io_axi_in_arvalid),
    .io_axi_in_rready(axi_io_axi_in_rready),
    .io_axi_in_awaddr(axi_io_axi_in_awaddr),
    .io_axi_in_awlen(axi_io_axi_in_awlen),
    .io_axi_in_awvalid(axi_io_axi_in_awvalid),
    .io_axi_in_wdata(axi_io_axi_in_wdata),
    .io_axi_in_wstrb(axi_io_axi_in_wstrb),
    .io_axi_in_wvalid(axi_io_axi_in_wvalid),
    .io_axi_in_bready(axi_io_axi_in_bready),
    .io_axi_out_rdata(axi_io_axi_out_rdata),
    .io_axi_out_rlast(axi_io_axi_out_rlast),
    .io_axi_out_rvalid(axi_io_axi_out_rvalid),
    .io_axi_out_wready(axi_io_axi_out_wready),
    .io_axi_out_bvalid(axi_io_axi_out_bvalid)
  );
  DPI dpi ( // @[top.scala 114:21]
    .flag(dpi_flag),
    .ecall_flag(dpi_ecall_flag),
    .pc(dpi_pc)
  );
  assign io_inst = IFU_io_inst; // @[top.scala 110:13]
  assign io_pc = IFU_io_to_ds_pc; // @[top.scala 108:11]
  assign io_step = diff_step; // @[top.scala 113:13]
  assign Register_clock = clock;
  assign Register_io_raddr1 = IDU_io_raddr1; // @[top.scala 54:20]
  assign Register_io_raddr2 = IDU_io_raddr2; // @[top.scala 55:20]
  assign Register_io_we = WBU_io_we; // @[top.scala 104:16]
  assign Register_io_waddr = WBU_io_waddr; // @[top.scala 105:19]
  assign Register_io_wdata = WBU_io_wdata; // @[top.scala 106:19]
  assign IFU_clock = clock;
  assign IFU_reset = reset;
  assign IFU_io_ds_allowin = IDU_io_ds_allowin; // @[top.scala 42:20]
  assign IFU_io_br_taken = IDU_io_br_taken; // @[top.scala 43:18]
  assign IFU_io_br_target = IDU_io_br_target; // @[top.scala 44:19]
  assign IFU_io_axi_in_rdata = i_cache_io_to_ifu_rdata; // @[top.scala 29:16]
  assign IFU_io_axi_in_rlast = i_cache_io_to_ifu_rlast; // @[top.scala 29:16]
  assign IFU_io_axi_in_rvalid = i_cache_io_to_ifu_rvalid; // @[top.scala 29:16]
  assign IFU_io_fence = IDU_io_fence; // @[top.scala 46:15]
  assign IFU_io_cache_init = i_cache_io_cache_init; // @[top.scala 47:20]
  assign IDU_clock = clock;
  assign IDU_reset = reset;
  assign IDU_io_pc = IFU_io_to_ds_pc; // @[top.scala 50:12]
  assign IDU_io_fs_to_ds_valid = IFU_io_fs_to_ds_valid; // @[top.scala 51:24]
  assign IDU_io_es_allowin = EXU_io_es_allowin; // @[top.scala 52:20]
  assign IDU_io_from_fs_inst = IFU_io_inst; // @[top.scala 53:22]
  assign IDU_io_rdata1 = Register_io_rdata1; // @[top.scala 56:16]
  assign IDU_io_rdata2 = Register_io_rdata2; // @[top.scala 57:16]
  assign IDU_io_es_ld = EXU_io_es_ld; // @[top.scala 73:15]
  assign IDU_io_es_fwd_res = EXU_io_es_fwd_res; // @[top.scala 68:20]
  assign IDU_io_ms_fwd_res = LSU_io_ms_fwd_res; // @[top.scala 70:20]
  assign IDU_io_ws_fwd_res = WBU_io_ws_fwd_res; // @[top.scala 72:20]
  assign IDU_io_es_fwd_ready = EXU_io_es_fwd_ready; // @[top.scala 67:22]
  assign IDU_io_ms_fwd_ready = LSU_io_ms_fwd_ready; // @[top.scala 69:22]
  assign IDU_io_es_rf_we = EXU_io_es_rf_we; // @[top.scala 60:18]
  assign IDU_io_ms_rf_we = LSU_io_ms_rf_we; // @[top.scala 63:18]
  assign IDU_io_ws_rf_we = WBU_io_ws_rf_we; // @[top.scala 66:18]
  assign IDU_io_es_valid = EXU_io_es_valid; // @[top.scala 58:18]
  assign IDU_io_ms_valid = LSU_io_ms_valid; // @[top.scala 61:18]
  assign IDU_io_ws_valid = WBU_io_ws_valid; // @[top.scala 64:18]
  assign IDU_io_es_rf_dst = EXU_io_es_rf_dst; // @[top.scala 59:19]
  assign IDU_io_ms_rf_dst = LSU_io_ms_rf_dst; // @[top.scala 62:19]
  assign IDU_io_ws_rf_dst = WBU_io_ws_rf_dst; // @[top.scala 65:19]
  assign EXU_clock = clock;
  assign EXU_reset = reset;
  assign EXU_io_pc = IDU_io_to_es_pc; // @[top.scala 75:12]
  assign EXU_io_ds_to_es_valid = IDU_io_ds_to_es_valid; // @[top.scala 76:24]
  assign EXU_io_ms_allowin = LSU_io_ms_allowin; // @[top.scala 77:20]
  assign EXU_io_ALUop = IDU_io_ALUop; // @[top.scala 78:15]
  assign EXU_io_src1_value = IDU_io_src1; // @[top.scala 79:20]
  assign EXU_io_src2_value = IDU_io_src2; // @[top.scala 80:20]
  assign EXU_io_rf_dst = IDU_io_rf_dst; // @[top.scala 81:16]
  assign EXU_io_store_data = IDU_io_store_data; // @[top.scala 82:20]
  assign EXU_io_load_type = IDU_io_load_type; // @[top.scala 84:19]
  assign EXU_io_ctrl_sign_reg_write = IDU_io_ctrl_sign_reg_write; // @[top.scala 83:19]
  assign EXU_io_ctrl_sign_Writemem_en = IDU_io_ctrl_sign_Writemem_en; // @[top.scala 83:19]
  assign EXU_io_ctrl_sign_Readmem_en = IDU_io_ctrl_sign_Readmem_en; // @[top.scala 83:19]
  assign EXU_io_ctrl_sign_Wmask = IDU_io_ctrl_sign_Wmask; // @[top.scala 83:19]
  assign LSU_clock = clock;
  assign LSU_reset = reset;
  assign LSU_io_pc = EXU_io_to_ms_pc; // @[top.scala 86:12]
  assign LSU_io_es_to_ms_valid = EXU_io_es_to_ms_valid; // @[top.scala 87:24]
  assign LSU_io_rf_we = EXU_io_to_ms_rf_we; // @[top.scala 89:15]
  assign LSU_io_rf_dst = EXU_io_to_ms_rf_dst; // @[top.scala 90:16]
  assign LSU_io_alu_res = EXU_io_to_ms_alures; // @[top.scala 91:17]
  assign LSU_io_store_data = EXU_io_to_ms_store_data; // @[top.scala 92:20]
  assign LSU_io_load_type = EXU_io_to_ms_load_type; // @[top.scala 97:19]
  assign LSU_io_wen = EXU_io_to_ms_wen; // @[top.scala 93:13]
  assign LSU_io_wstrb = EXU_io_to_ms_wstrb; // @[top.scala 94:15]
  assign LSU_io_ren = EXU_io_to_ms_ren; // @[top.scala 95:13]
  assign LSU_io_maddr = EXU_io_to_ms_maddr; // @[top.scala 96:15]
  assign LSU_io_axi_in_rdata = d_cache_io_to_lsu_rdata; // @[top.scala 34:16]
  assign LSU_io_axi_in_rvalid = d_cache_io_to_lsu_rvalid; // @[top.scala 34:16]
  assign LSU_io_axi_in_wready = d_cache_io_to_lsu_wready; // @[top.scala 34:16]
  assign WBU_clock = clock;
  assign WBU_reset = reset;
  assign WBU_io_pc = LSU_io_to_ws_pc; // @[top.scala 99:12]
  assign WBU_io_ms_to_ws_valid = LSU_io_ms_to_ws_valid; // @[top.scala 100:24]
  assign WBU_io_ms_final_res = LSU_io_ms_final_res; // @[top.scala 101:22]
  assign WBU_io_rf_we = LSU_io_to_ws_rf_we; // @[top.scala 102:15]
  assign WBU_io_rf_dst = LSU_io_to_ws_rf_dst; // @[top.scala 103:16]
  assign arbiter_clock = clock;
  assign arbiter_reset = reset;
  assign arbiter_io_ifu_axi_in_araddr = i_cache_io_to_axi_araddr; // @[top.scala 27:27]
  assign arbiter_io_ifu_axi_in_arlen = i_cache_io_to_axi_arlen; // @[top.scala 27:27]
  assign arbiter_io_ifu_axi_in_arvalid = i_cache_io_to_axi_arvalid; // @[top.scala 27:27]
  assign arbiter_io_ifu_axi_in_rready = i_cache_io_to_axi_rready; // @[top.scala 27:27]
  assign arbiter_io_lsu_axi_in_araddr = d_cache_io_to_axi_araddr; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_arlen = d_cache_io_to_axi_arlen; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_arvalid = d_cache_io_to_axi_arvalid; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_rready = d_cache_io_to_axi_rready; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_awaddr = d_cache_io_to_axi_awaddr; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_awlen = d_cache_io_to_axi_awlen; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_awvalid = d_cache_io_to_axi_awvalid; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_wdata = d_cache_io_to_axi_wdata; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_wstrb = d_cache_io_to_axi_wstrb; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_wvalid = d_cache_io_to_axi_wvalid; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_bready = d_cache_io_to_axi_bready; // @[top.scala 32:27]
  assign arbiter_io_axi_in_rdata = axi_io_axi_out_rdata; // @[top.scala 37:23]
  assign arbiter_io_axi_in_rlast = axi_io_axi_out_rlast; // @[top.scala 37:23]
  assign arbiter_io_axi_in_rvalid = axi_io_axi_out_rvalid; // @[top.scala 37:23]
  assign arbiter_io_axi_in_wready = axi_io_axi_out_wready; // @[top.scala 37:23]
  assign arbiter_io_axi_in_bvalid = axi_io_axi_out_bvalid; // @[top.scala 37:23]
  assign i_cache_clock = clock;
  assign i_cache_reset = reset;
  assign i_cache_io_from_ifu_araddr = IFU_io_axi_out_araddr; // @[top.scala 30:25]
  assign i_cache_io_from_ifu_arvalid = IFU_io_axi_out_arvalid; // @[top.scala 30:25]
  assign i_cache_io_from_ifu_rready = IFU_io_axi_out_rready; // @[top.scala 30:25]
  assign i_cache_io_from_axi_rdata = arbiter_io_ifu_axi_out_rdata; // @[top.scala 28:25]
  assign i_cache_io_from_axi_rlast = arbiter_io_ifu_axi_out_rlast; // @[top.scala 28:25]
  assign i_cache_io_from_axi_rvalid = arbiter_io_ifu_axi_out_rvalid; // @[top.scala 28:25]
  assign i_cache_io_clear_cache = IFU_io_clear_cache; // @[top.scala 48:28]
  assign d_cache_clock = clock;
  assign d_cache_reset = reset;
  assign d_cache_io_from_lsu_araddr = LSU_io_axi_out_araddr; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_arvalid = LSU_io_axi_out_arvalid; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_awaddr = LSU_io_axi_out_awaddr; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_awvalid = LSU_io_axi_out_awvalid; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_wdata = LSU_io_axi_out_wdata; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_wstrb = LSU_io_axi_out_wstrb; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_wvalid = LSU_io_axi_out_wvalid; // @[top.scala 35:25]
  assign d_cache_io_from_axi_rdata = arbiter_io_lsu_axi_out_rdata; // @[top.scala 33:25]
  assign d_cache_io_from_axi_rlast = arbiter_io_lsu_axi_out_rlast; // @[top.scala 33:25]
  assign d_cache_io_from_axi_rvalid = arbiter_io_lsu_axi_out_rvalid; // @[top.scala 33:25]
  assign d_cache_io_from_axi_wready = arbiter_io_lsu_axi_out_wready; // @[top.scala 33:25]
  assign d_cache_io_from_axi_bvalid = arbiter_io_lsu_axi_out_bvalid; // @[top.scala 33:25]
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_axi_in_araddr = arbiter_io_axi_out_araddr; // @[top.scala 38:19]
  assign axi_io_axi_in_arlen = arbiter_io_axi_out_arlen; // @[top.scala 38:19]
  assign axi_io_axi_in_arvalid = arbiter_io_axi_out_arvalid; // @[top.scala 38:19]
  assign axi_io_axi_in_rready = arbiter_io_axi_out_rready; // @[top.scala 38:19]
  assign axi_io_axi_in_awaddr = arbiter_io_axi_out_awaddr; // @[top.scala 38:19]
  assign axi_io_axi_in_awlen = arbiter_io_axi_out_awlen; // @[top.scala 38:19]
  assign axi_io_axi_in_awvalid = arbiter_io_axi_out_awvalid; // @[top.scala 38:19]
  assign axi_io_axi_in_wdata = arbiter_io_axi_out_wdata; // @[top.scala 38:19]
  assign axi_io_axi_in_wstrb = arbiter_io_axi_out_wstrb; // @[top.scala 38:19]
  assign axi_io_axi_in_wvalid = arbiter_io_axi_out_wvalid; // @[top.scala 38:19]
  assign axi_io_axi_in_bready = arbiter_io_axi_out_bready; // @[top.scala 38:19]
  assign dpi_flag = {{31'd0}, IDU_io_ALUop == 32'h2}; // @[top.scala 115:17]
  assign dpi_ecall_flag = {{31'd0}, IDU_io_ALUop == 32'h3d}; // @[top.scala 116:23]
  assign dpi_pc = WBU_io_ws_valid ? WBU_io_ws_pc : _dpi_io_pc_T_2; // @[top.scala 117:21]
  always @(posedge clock) begin
    if (reset) begin // @[top.scala 111:28]
      diff_step <= 1'h0; // @[top.scala 111:28]
    end else begin
      diff_step <= WBU_io_ws_valid; // @[top.scala 112:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  diff_step = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
