module Register(
  input         clock,
  input  [4:0]  io_raddr1,
  input  [4:0]  io_raddr2,
  output [63:0] io_rdata1,
  output [63:0] io_rdata2,
  input         io_we,
  input  [4:0]  io_waddr,
  input  [63:0] io_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [63:0] Reg [0:31]; // @[register.scala 18:18]
  wire  Reg_io_rdata1_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_io_rdata1_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_io_rdata1_MPORT_data; // @[register.scala 18:18]
  wire  Reg_io_rdata2_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_io_rdata2_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_io_rdata2_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_0_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_0_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_0_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_1_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_1_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_1_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_2_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_2_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_2_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_3_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_3_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_3_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_4_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_4_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_4_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_5_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_5_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_5_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_6_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_6_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_6_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_7_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_7_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_7_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_8_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_8_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_8_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_9_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_9_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_9_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_10_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_10_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_10_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_11_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_11_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_11_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_12_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_12_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_12_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_13_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_13_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_13_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_14_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_14_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_14_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_15_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_15_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_15_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_16_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_16_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_16_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_17_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_17_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_17_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_18_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_18_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_18_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_19_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_19_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_19_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_20_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_20_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_20_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_21_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_21_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_21_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_22_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_22_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_22_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_23_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_23_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_23_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_24_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_24_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_24_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_25_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_25_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_25_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_26_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_26_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_26_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_27_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_27_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_27_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_28_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_28_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_28_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_29_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_29_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_29_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_30_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_30_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_30_MPORT_data; // @[register.scala 18:18]
  wire  Reg_reg_trace_io_input_reg_31_MPORT_en; // @[register.scala 18:18]
  wire [4:0] Reg_reg_trace_io_input_reg_31_MPORT_addr; // @[register.scala 18:18]
  wire [63:0] Reg_reg_trace_io_input_reg_31_MPORT_data; // @[register.scala 18:18]
  wire [63:0] Reg_MPORT_data; // @[register.scala 18:18]
  wire [4:0] Reg_MPORT_addr; // @[register.scala 18:18]
  wire  Reg_MPORT_mask; // @[register.scala 18:18]
  wire  Reg_MPORT_en; // @[register.scala 18:18]
  wire [63:0] reg_trace_input_reg_0; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_1; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_2; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_3; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_4; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_5; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_6; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_7; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_8; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_9; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_10; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_11; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_12; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_13; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_14; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_15; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_16; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_17; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_18; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_19; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_20; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_21; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_22; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_23; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_24; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_25; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_26; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_27; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_28; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_29; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_30; // @[register.scala 24:27]
  wire [63:0] reg_trace_input_reg_31; // @[register.scala 24:27]
  wire  _T = io_waddr != 5'h0; // @[register.scala 19:25]
  traceregs reg_trace ( // @[register.scala 24:27]
    .input_reg_0(reg_trace_input_reg_0),
    .input_reg_1(reg_trace_input_reg_1),
    .input_reg_2(reg_trace_input_reg_2),
    .input_reg_3(reg_trace_input_reg_3),
    .input_reg_4(reg_trace_input_reg_4),
    .input_reg_5(reg_trace_input_reg_5),
    .input_reg_6(reg_trace_input_reg_6),
    .input_reg_7(reg_trace_input_reg_7),
    .input_reg_8(reg_trace_input_reg_8),
    .input_reg_9(reg_trace_input_reg_9),
    .input_reg_10(reg_trace_input_reg_10),
    .input_reg_11(reg_trace_input_reg_11),
    .input_reg_12(reg_trace_input_reg_12),
    .input_reg_13(reg_trace_input_reg_13),
    .input_reg_14(reg_trace_input_reg_14),
    .input_reg_15(reg_trace_input_reg_15),
    .input_reg_16(reg_trace_input_reg_16),
    .input_reg_17(reg_trace_input_reg_17),
    .input_reg_18(reg_trace_input_reg_18),
    .input_reg_19(reg_trace_input_reg_19),
    .input_reg_20(reg_trace_input_reg_20),
    .input_reg_21(reg_trace_input_reg_21),
    .input_reg_22(reg_trace_input_reg_22),
    .input_reg_23(reg_trace_input_reg_23),
    .input_reg_24(reg_trace_input_reg_24),
    .input_reg_25(reg_trace_input_reg_25),
    .input_reg_26(reg_trace_input_reg_26),
    .input_reg_27(reg_trace_input_reg_27),
    .input_reg_28(reg_trace_input_reg_28),
    .input_reg_29(reg_trace_input_reg_29),
    .input_reg_30(reg_trace_input_reg_30),
    .input_reg_31(reg_trace_input_reg_31)
  );
  assign Reg_io_rdata1_MPORT_en = 1'h1;
  assign Reg_io_rdata1_MPORT_addr = io_raddr1;
  assign Reg_io_rdata1_MPORT_data = Reg[Reg_io_rdata1_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_io_rdata2_MPORT_en = 1'h1;
  assign Reg_io_rdata2_MPORT_addr = io_raddr2;
  assign Reg_io_rdata2_MPORT_data = Reg[Reg_io_rdata2_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_0_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_0_MPORT_addr = 5'h0;
  assign Reg_reg_trace_io_input_reg_0_MPORT_data = Reg[Reg_reg_trace_io_input_reg_0_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_1_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_1_MPORT_addr = 5'h1;
  assign Reg_reg_trace_io_input_reg_1_MPORT_data = Reg[Reg_reg_trace_io_input_reg_1_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_2_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_2_MPORT_addr = 5'h2;
  assign Reg_reg_trace_io_input_reg_2_MPORT_data = Reg[Reg_reg_trace_io_input_reg_2_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_3_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_3_MPORT_addr = 5'h3;
  assign Reg_reg_trace_io_input_reg_3_MPORT_data = Reg[Reg_reg_trace_io_input_reg_3_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_4_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_4_MPORT_addr = 5'h4;
  assign Reg_reg_trace_io_input_reg_4_MPORT_data = Reg[Reg_reg_trace_io_input_reg_4_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_5_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_5_MPORT_addr = 5'h5;
  assign Reg_reg_trace_io_input_reg_5_MPORT_data = Reg[Reg_reg_trace_io_input_reg_5_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_6_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_6_MPORT_addr = 5'h6;
  assign Reg_reg_trace_io_input_reg_6_MPORT_data = Reg[Reg_reg_trace_io_input_reg_6_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_7_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_7_MPORT_addr = 5'h7;
  assign Reg_reg_trace_io_input_reg_7_MPORT_data = Reg[Reg_reg_trace_io_input_reg_7_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_8_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_8_MPORT_addr = 5'h8;
  assign Reg_reg_trace_io_input_reg_8_MPORT_data = Reg[Reg_reg_trace_io_input_reg_8_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_9_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_9_MPORT_addr = 5'h9;
  assign Reg_reg_trace_io_input_reg_9_MPORT_data = Reg[Reg_reg_trace_io_input_reg_9_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_10_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_10_MPORT_addr = 5'ha;
  assign Reg_reg_trace_io_input_reg_10_MPORT_data = Reg[Reg_reg_trace_io_input_reg_10_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_11_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_11_MPORT_addr = 5'hb;
  assign Reg_reg_trace_io_input_reg_11_MPORT_data = Reg[Reg_reg_trace_io_input_reg_11_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_12_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_12_MPORT_addr = 5'hc;
  assign Reg_reg_trace_io_input_reg_12_MPORT_data = Reg[Reg_reg_trace_io_input_reg_12_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_13_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_13_MPORT_addr = 5'hd;
  assign Reg_reg_trace_io_input_reg_13_MPORT_data = Reg[Reg_reg_trace_io_input_reg_13_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_14_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_14_MPORT_addr = 5'he;
  assign Reg_reg_trace_io_input_reg_14_MPORT_data = Reg[Reg_reg_trace_io_input_reg_14_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_15_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_15_MPORT_addr = 5'hf;
  assign Reg_reg_trace_io_input_reg_15_MPORT_data = Reg[Reg_reg_trace_io_input_reg_15_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_16_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_16_MPORT_addr = 5'h10;
  assign Reg_reg_trace_io_input_reg_16_MPORT_data = Reg[Reg_reg_trace_io_input_reg_16_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_17_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_17_MPORT_addr = 5'h11;
  assign Reg_reg_trace_io_input_reg_17_MPORT_data = Reg[Reg_reg_trace_io_input_reg_17_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_18_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_18_MPORT_addr = 5'h12;
  assign Reg_reg_trace_io_input_reg_18_MPORT_data = Reg[Reg_reg_trace_io_input_reg_18_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_19_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_19_MPORT_addr = 5'h13;
  assign Reg_reg_trace_io_input_reg_19_MPORT_data = Reg[Reg_reg_trace_io_input_reg_19_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_20_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_20_MPORT_addr = 5'h14;
  assign Reg_reg_trace_io_input_reg_20_MPORT_data = Reg[Reg_reg_trace_io_input_reg_20_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_21_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_21_MPORT_addr = 5'h15;
  assign Reg_reg_trace_io_input_reg_21_MPORT_data = Reg[Reg_reg_trace_io_input_reg_21_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_22_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_22_MPORT_addr = 5'h16;
  assign Reg_reg_trace_io_input_reg_22_MPORT_data = Reg[Reg_reg_trace_io_input_reg_22_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_23_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_23_MPORT_addr = 5'h17;
  assign Reg_reg_trace_io_input_reg_23_MPORT_data = Reg[Reg_reg_trace_io_input_reg_23_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_24_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_24_MPORT_addr = 5'h18;
  assign Reg_reg_trace_io_input_reg_24_MPORT_data = Reg[Reg_reg_trace_io_input_reg_24_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_25_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_25_MPORT_addr = 5'h19;
  assign Reg_reg_trace_io_input_reg_25_MPORT_data = Reg[Reg_reg_trace_io_input_reg_25_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_26_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_26_MPORT_addr = 5'h1a;
  assign Reg_reg_trace_io_input_reg_26_MPORT_data = Reg[Reg_reg_trace_io_input_reg_26_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_27_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_27_MPORT_addr = 5'h1b;
  assign Reg_reg_trace_io_input_reg_27_MPORT_data = Reg[Reg_reg_trace_io_input_reg_27_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_28_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_28_MPORT_addr = 5'h1c;
  assign Reg_reg_trace_io_input_reg_28_MPORT_data = Reg[Reg_reg_trace_io_input_reg_28_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_29_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_29_MPORT_addr = 5'h1d;
  assign Reg_reg_trace_io_input_reg_29_MPORT_data = Reg[Reg_reg_trace_io_input_reg_29_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_30_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_30_MPORT_addr = 5'h1e;
  assign Reg_reg_trace_io_input_reg_30_MPORT_data = Reg[Reg_reg_trace_io_input_reg_30_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_reg_trace_io_input_reg_31_MPORT_en = 1'h1;
  assign Reg_reg_trace_io_input_reg_31_MPORT_addr = 5'h1f;
  assign Reg_reg_trace_io_input_reg_31_MPORT_data = Reg[Reg_reg_trace_io_input_reg_31_MPORT_addr]; // @[register.scala 18:18]
  assign Reg_MPORT_data = io_wdata;
  assign Reg_MPORT_addr = io_waddr;
  assign Reg_MPORT_mask = 1'h1;
  assign Reg_MPORT_en = io_we & _T;
  assign io_rdata1 = io_raddr1 == 5'h0 ? 64'h0 : Reg_io_rdata1_MPORT_data; // @[register.scala 22:21]
  assign io_rdata2 = io_raddr2 == 5'h0 ? 64'h0 : Reg_io_rdata2_MPORT_data; // @[register.scala 23:21]
  assign reg_trace_input_reg_0 = Reg_reg_trace_io_input_reg_0_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_1 = Reg_reg_trace_io_input_reg_1_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_2 = Reg_reg_trace_io_input_reg_2_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_3 = Reg_reg_trace_io_input_reg_3_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_4 = Reg_reg_trace_io_input_reg_4_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_5 = Reg_reg_trace_io_input_reg_5_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_6 = Reg_reg_trace_io_input_reg_6_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_7 = Reg_reg_trace_io_input_reg_7_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_8 = Reg_reg_trace_io_input_reg_8_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_9 = Reg_reg_trace_io_input_reg_9_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_10 = Reg_reg_trace_io_input_reg_10_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_11 = Reg_reg_trace_io_input_reg_11_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_12 = Reg_reg_trace_io_input_reg_12_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_13 = Reg_reg_trace_io_input_reg_13_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_14 = Reg_reg_trace_io_input_reg_14_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_15 = Reg_reg_trace_io_input_reg_15_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_16 = Reg_reg_trace_io_input_reg_16_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_17 = Reg_reg_trace_io_input_reg_17_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_18 = Reg_reg_trace_io_input_reg_18_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_19 = Reg_reg_trace_io_input_reg_19_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_20 = Reg_reg_trace_io_input_reg_20_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_21 = Reg_reg_trace_io_input_reg_21_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_22 = Reg_reg_trace_io_input_reg_22_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_23 = Reg_reg_trace_io_input_reg_23_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_24 = Reg_reg_trace_io_input_reg_24_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_25 = Reg_reg_trace_io_input_reg_25_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_26 = Reg_reg_trace_io_input_reg_26_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_27 = Reg_reg_trace_io_input_reg_27_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_28 = Reg_reg_trace_io_input_reg_28_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_29 = Reg_reg_trace_io_input_reg_29_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_30 = Reg_reg_trace_io_input_reg_30_MPORT_data; // @[register.scala 26:57]
  assign reg_trace_input_reg_31 = Reg_reg_trace_io_input_reg_31_MPORT_data; // @[register.scala 26:57]
  always @(posedge clock) begin
    if (Reg_MPORT_en & Reg_MPORT_mask) begin
      Reg[Reg_MPORT_addr] <= Reg_MPORT_data; // @[register.scala 18:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    Reg[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU(
  input         clock,
  input         reset,
  input         io_ds_allowin,
  input         io_ds_ready_go,
  input         io_ds_valid,
  input         io_br_taken,
  input  [63:0] io_br_target,
  output [63:0] io_to_ds_pc,
  output        io_fs_to_ds_valid,
  output [31:0] io_inst,
  input         io_axi_in_arready,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  input         io_fence,
  output        io_clear_cache,
  input         io_cache_init
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] br_target; // @[IFU.scala 31:28]
  reg  fs_valid; // @[IFU.scala 36:27]
  reg [63:0] fs_pc_next; // @[IFU.scala 42:29]
  reg  cache_init; // @[IFU.scala 43:29]
  wire  _T_1 = fs_valid & io_ds_allowin; // @[IFU.scala 46:31]
  wire  _GEN_1 = fs_valid & io_ds_allowin & cache_init ? 1'h0 : cache_init; // @[IFU.scala 46:60 47:20 43:29]
  wire  _GEN_2 = io_cache_init | _GEN_1; // @[IFU.scala 44:24 45:20]
  reg [63:0] fs_pc; // @[IFU.scala 50:24]
  reg [31:0] fs_inst; // @[IFU.scala 51:26]
  wire [63:0] seq_pc = fs_pc + 64'h4; // @[IFU.scala 74:24]
  wire [63:0] _pc_next_T = io_ds_valid ? io_br_target : br_target; // @[IFU.scala 75:35]
  wire [63:0] pc_next = io_br_taken ? _pc_next_T : seq_pc; // @[IFU.scala 75:19]
  wire  fs_allowin = ~fs_valid | _T_1; // @[IFU.scala 83:29]
  assign io_to_ds_pc = fs_pc; // @[IFU.scala 95:17]
  assign io_fs_to_ds_valid = fs_valid; // @[IFU.scala 82:33]
  assign io_inst = fs_inst; // @[IFU.scala 121:13]
  assign io_axi_out_araddr = pc_next[31:0]; // @[IFU.scala 105:23]
  assign io_axi_out_arvalid = io_ds_ready_go; // @[IFU.scala 106:24]
  assign io_axi_out_rready = ~fs_valid | _T_1; // @[IFU.scala 83:29]
  assign io_clear_cache = io_fence & ~cache_init; // @[IFU.scala 55:32]
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 31:28]
      br_target <= 64'h0; // @[IFU.scala 31:28]
    end else if (io_ds_valid & io_ds_ready_go) begin // @[IFU.scala 32:40]
      br_target <= io_br_target; // @[IFU.scala 33:19]
    end
    if (reset) begin // @[IFU.scala 36:27]
      fs_valid <= 1'h0; // @[IFU.scala 36:27]
    end else if (fs_allowin) begin // @[IFU.scala 84:21]
      fs_valid <= io_axi_in_rvalid; // @[IFU.scala 85:18]
    end
    if (reset) begin // @[IFU.scala 42:29]
      fs_pc_next <= 64'h0; // @[IFU.scala 42:29]
    end else if (io_axi_in_arready & io_ds_ready_go) begin // @[IFU.scala 76:46]
      if (io_br_taken) begin // @[IFU.scala 75:19]
        if (io_ds_valid) begin // @[IFU.scala 75:35]
          fs_pc_next <= io_br_target;
        end else begin
          fs_pc_next <= br_target;
        end
      end else begin
        fs_pc_next <= seq_pc;
      end
    end
    if (reset) begin // @[IFU.scala 43:29]
      cache_init <= 1'h0; // @[IFU.scala 43:29]
    end else begin
      cache_init <= _GEN_2;
    end
    if (reset) begin // @[IFU.scala 50:24]
      fs_pc <= 64'h7ffffffc; // @[IFU.scala 50:24]
    end else if (io_axi_in_rvalid & fs_allowin) begin // @[IFU.scala 87:36]
      fs_pc <= fs_pc_next; // @[IFU.scala 88:15]
    end
    if (reset) begin // @[IFU.scala 51:26]
      fs_inst <= 32'h0; // @[IFU.scala 51:26]
    end else if (io_axi_in_rvalid & fs_allowin) begin // @[IFU.scala 87:36]
      fs_inst <= io_axi_in_rdata[31:0]; // @[IFU.scala 89:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  br_target = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  fs_valid = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  fs_pc_next = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  cache_init = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  fs_pc = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  fs_inst = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module csr_reg(
  input         clock,
  input         io_wen1,
  input         io_wen2,
  input  [1:0]  io_waddr1,
  input  [63:0] io_wdata1,
  input  [63:0] io_wdata2,
  input  [1:0]  io_raddr,
  output [63:0] io_rdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [63:0] CSR_Reg [0:3]; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_io_rdata_MPORT_en; // @[csr_reg.scala 19:22]
  wire [1:0] CSR_Reg_io_rdata_MPORT_addr; // @[csr_reg.scala 19:22]
  wire [63:0] CSR_Reg_io_rdata_MPORT_data; // @[csr_reg.scala 19:22]
  wire [63:0] CSR_Reg_MPORT_data; // @[csr_reg.scala 19:22]
  wire [1:0] CSR_Reg_MPORT_addr; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_MPORT_mask; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_MPORT_en; // @[csr_reg.scala 19:22]
  wire [63:0] CSR_Reg_MPORT_1_data; // @[csr_reg.scala 19:22]
  wire [1:0] CSR_Reg_MPORT_1_addr; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_MPORT_1_mask; // @[csr_reg.scala 19:22]
  wire  CSR_Reg_MPORT_1_en; // @[csr_reg.scala 19:22]
  assign CSR_Reg_io_rdata_MPORT_en = 1'h1;
  assign CSR_Reg_io_rdata_MPORT_addr = io_raddr;
  assign CSR_Reg_io_rdata_MPORT_data = CSR_Reg[CSR_Reg_io_rdata_MPORT_addr]; // @[csr_reg.scala 19:22]
  assign CSR_Reg_MPORT_data = io_wdata1;
  assign CSR_Reg_MPORT_addr = io_waddr1;
  assign CSR_Reg_MPORT_mask = 1'h1;
  assign CSR_Reg_MPORT_en = io_wen1;
  assign CSR_Reg_MPORT_1_data = io_wdata2;
  assign CSR_Reg_MPORT_1_addr = 2'h3;
  assign CSR_Reg_MPORT_1_mask = 1'h1;
  assign CSR_Reg_MPORT_1_en = io_wen2;
  assign io_rdata = CSR_Reg_io_rdata_MPORT_data; // @[csr_reg.scala 26:14]
  always @(posedge clock) begin
    if (CSR_Reg_MPORT_en & CSR_Reg_MPORT_mask) begin
      CSR_Reg[CSR_Reg_MPORT_addr] <= CSR_Reg_MPORT_data; // @[csr_reg.scala 19:22]
    end
    if (CSR_Reg_MPORT_1_en & CSR_Reg_MPORT_1_mask) begin
      CSR_Reg[CSR_Reg_MPORT_1_addr] <= CSR_Reg_MPORT_1_data; // @[csr_reg.scala 19:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    CSR_Reg[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_fs_to_ds_valid,
  output        io_ds_to_es_valid,
  input         io_es_allowin,
  input  [31:0] io_from_fs_inst,
  output        io_br_taken,
  output [63:0] io_br_target,
  output        io_ds_allowin,
  output        io_ds_ready_go,
  output        io_fence,
  output [4:0]  io_raddr1,
  output [4:0]  io_raddr2,
  input  [63:0] io_rdata1,
  input  [63:0] io_rdata2,
  output [63:0] io_to_es_pc,
  output [31:0] io_ALUop,
  output [63:0] io_src1,
  output [63:0] io_src2,
  output [4:0]  io_rf_dst,
  output [63:0] io_store_data,
  output        io_ctrl_sign_reg_write,
  output        io_ctrl_sign_Writemem_en,
  output        io_ctrl_sign_Readmem_en,
  output [7:0]  io_ctrl_sign_Wmask,
  output [2:0]  io_load_type,
  input         io_es_ld,
  input  [63:0] io_es_fwd_res,
  input  [63:0] io_ms_fwd_res,
  input  [63:0] io_ws_fwd_res,
  input         io_es_fwd_ready,
  input         io_ms_fwd_ready,
  input         io_es_rf_we,
  input         io_ms_rf_we,
  input         io_ws_rf_we,
  input         io_es_valid,
  input         io_ms_valid,
  input         io_ws_valid,
  input  [4:0]  io_es_rf_dst,
  input  [4:0]  io_ms_rf_dst,
  input  [4:0]  io_ws_rf_dst,
  output        io_ds_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  csr_reg_clock; // @[IDU.scala 449:21]
  wire  csr_reg_io_wen1; // @[IDU.scala 449:21]
  wire  csr_reg_io_wen2; // @[IDU.scala 449:21]
  wire [1:0] csr_reg_io_waddr1; // @[IDU.scala 449:21]
  wire [63:0] csr_reg_io_wdata1; // @[IDU.scala 449:21]
  wire [63:0] csr_reg_io_wdata2; // @[IDU.scala 449:21]
  wire [1:0] csr_reg_io_raddr; // @[IDU.scala 449:21]
  wire [63:0] csr_reg_io_rdata; // @[IDU.scala 449:21]
  reg  ds_valid; // @[IDU.scala 112:27]
  reg [63:0] ds_pc; // @[IDU.scala 116:24]
  reg [31:0] inst; // @[IDU.scala 118:23]
  reg  br_taken_cancel; // @[IDU.scala 122:34]
  wire [31:0] _src1_is_pc_T = inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_1 = 32'h6f == _src1_is_pc_T; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_3 = 32'h17 == _src1_is_pc_T; // @[Lookup.scala 31:38]
  wire [31:0] _src1_is_pc_T_4 = inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_5 = 32'h1063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_7 = 32'h63 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_9 = 32'h5063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_11 = 32'h4063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_13 = 32'h6063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _src1_is_pc_T_15 = 32'h7063 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  src1_is_pc = _src1_is_pc_T_1 | (_src1_is_pc_T_3 | (_src1_is_pc_T_5 | (_src1_is_pc_T_7 | (_src1_is_pc_T_9 | (
    _src1_is_pc_T_11 | (_src1_is_pc_T_13 | _src1_is_pc_T_15)))))); // @[Lookup.scala 34:39]
  wire  _inst_type_T_1 = 32'h13 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_5 = 32'h37 == _src1_is_pc_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_9 = 32'h67 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_11 = 32'h3023 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_13 = 32'h3013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_15 = 32'h2003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_16 = inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_17 = 32'h3b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_19 = 32'h40000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_25 = 32'h3003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_27 = 32'h1b == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_29 = 32'h33 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_30 = inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_31 = 32'h40005013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_33 = 32'h4003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_35 = 32'h1023 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_37 = 32'h23 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_39 = 32'h6033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_41 = 32'h4013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_43 = 32'h7033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_45 = 32'h7013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_47 = 32'h4000003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_49 = 32'h103b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_51 = 32'h1013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_53 = 32'h5013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_55 = 32'h101b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_57 = 32'h4000501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_59 = 32'h501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_61 = 32'h4000503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_63 = 32'h503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_65 = 32'h3033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_67 = 32'h2033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_75 = 32'h2023 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_77 = 32'h1003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_79 = 32'h5003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_81 = 32'h2000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_83 = 32'h200003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_85 = 32'h200403b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_87 = 32'h200603b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_89 = 32'h4033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_91 = 32'h6013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_93 = 32'h2005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_95 = 32'h2004033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_97 = 32'h200503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_99 = 32'h200703b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_101 = 32'h2007033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_103 = 32'h2006033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_105 = 32'h1033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_107 = 32'h5033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_109 = 32'h40005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_111 = 32'h2013 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_113 = 32'h6003 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_115 = 32'h3 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_119 = 32'h73 == inst; // @[Lookup.scala 31:38]
  wire  _inst_type_T_121 = 32'h1073 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_123 = 32'h2073 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_125 = 32'h3073 == _src1_is_pc_T_4; // @[Lookup.scala 31:38]
  wire [6:0] _inst_type_T_126 = _inst_type_T_125 ? 7'h40 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_127 = _inst_type_T_123 ? 7'h40 : _inst_type_T_126; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_128 = _inst_type_T_121 ? 7'h40 : _inst_type_T_127; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_129 = _inst_type_T_119 ? 7'h40 : _inst_type_T_128; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_130 = _src1_is_pc_T_15 ? 7'h45 : _inst_type_T_129; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_131 = _inst_type_T_115 ? 7'h40 : _inst_type_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_132 = _inst_type_T_113 ? 7'h40 : _inst_type_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_133 = _inst_type_T_111 ? 7'h40 : _inst_type_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_134 = _inst_type_T_109 ? 7'h41 : _inst_type_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_135 = _inst_type_T_107 ? 7'h41 : _inst_type_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_136 = _inst_type_T_105 ? 7'h41 : _inst_type_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_137 = _inst_type_T_103 ? 7'h41 : _inst_type_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_138 = _inst_type_T_101 ? 7'h41 : _inst_type_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_139 = _inst_type_T_99 ? 7'h41 : _inst_type_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_140 = _inst_type_T_97 ? 7'h41 : _inst_type_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_141 = _inst_type_T_95 ? 7'h41 : _inst_type_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_142 = _inst_type_T_93 ? 7'h41 : _inst_type_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_143 = _inst_type_T_91 ? 7'h40 : _inst_type_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_144 = _inst_type_T_89 ? 7'h41 : _inst_type_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_145 = _inst_type_T_87 ? 7'h41 : _inst_type_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_146 = _inst_type_T_85 ? 7'h41 : _inst_type_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_147 = _inst_type_T_83 ? 7'h41 : _inst_type_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_148 = _inst_type_T_81 ? 7'h41 : _inst_type_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_149 = _inst_type_T_79 ? 7'h40 : _inst_type_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_150 = _inst_type_T_77 ? 7'h40 : _inst_type_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_151 = _inst_type_T_75 ? 7'h44 : _inst_type_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_152 = _src1_is_pc_T_13 ? 7'h45 : _inst_type_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_153 = _src1_is_pc_T_11 ? 7'h45 : _inst_type_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_154 = _src1_is_pc_T_9 ? 7'h45 : _inst_type_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_155 = _inst_type_T_67 ? 7'h41 : _inst_type_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_156 = _inst_type_T_65 ? 7'h41 : _inst_type_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_157 = _inst_type_T_63 ? 7'h41 : _inst_type_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_158 = _inst_type_T_61 ? 7'h41 : _inst_type_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_159 = _inst_type_T_59 ? 7'h40 : _inst_type_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_160 = _inst_type_T_57 ? 7'h40 : _inst_type_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_161 = _inst_type_T_55 ? 7'h40 : _inst_type_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_162 = _inst_type_T_53 ? 7'h40 : _inst_type_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_163 = _inst_type_T_51 ? 7'h40 : _inst_type_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_164 = _inst_type_T_49 ? 7'h41 : _inst_type_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_165 = _inst_type_T_47 ? 7'h41 : _inst_type_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_166 = _inst_type_T_45 ? 7'h40 : _inst_type_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_167 = _inst_type_T_43 ? 7'h41 : _inst_type_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_168 = _inst_type_T_41 ? 7'h40 : _inst_type_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_169 = _inst_type_T_39 ? 7'h41 : _inst_type_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_170 = _inst_type_T_37 ? 7'h44 : _inst_type_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_171 = _inst_type_T_35 ? 7'h44 : _inst_type_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_172 = _inst_type_T_33 ? 7'h40 : _inst_type_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_173 = _inst_type_T_31 ? 7'h40 : _inst_type_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_174 = _inst_type_T_29 ? 7'h41 : _inst_type_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_175 = _inst_type_T_27 ? 7'h40 : _inst_type_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_176 = _inst_type_T_25 ? 7'h40 : _inst_type_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_177 = _src1_is_pc_T_7 ? 7'h45 : _inst_type_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_178 = _src1_is_pc_T_5 ? 7'h45 : _inst_type_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_179 = _inst_type_T_19 ? 7'h41 : _inst_type_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_180 = _inst_type_T_17 ? 7'h41 : _inst_type_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_181 = _inst_type_T_15 ? 7'h40 : _inst_type_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_182 = _inst_type_T_13 ? 7'h40 : _inst_type_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_183 = _inst_type_T_11 ? 7'h44 : _inst_type_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_184 = _inst_type_T_9 ? 7'h40 : _inst_type_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_185 = _src1_is_pc_T_1 ? 7'h43 : _inst_type_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_186 = _inst_type_T_5 ? 7'h42 : _inst_type_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_187 = _src1_is_pc_T_3 ? 7'h42 : _inst_type_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_188 = _inst_type_T_1 ? 7'h40 : _inst_type_T_187; // @[Lookup.scala 34:39]
  wire [31:0] inst_type = {{25'd0}, _inst_type_T_188}; // @[IDU.scala 237:15 66:25]
  wire  _conflict_es_rs1_T_1 = inst_type == 32'h45; // @[IDU.scala 492:47]
  wire  _csr_write_T_10 = _inst_type_T_121 | (_inst_type_T_123 | _inst_type_T_125); // @[Lookup.scala 34:39]
  wire [1:0] csr_write = _inst_type_T_119 ? 2'h3 : {{1'd0}, _csr_write_T_10}; // @[Lookup.scala 34:39]
  wire  _conflict_es_rs1_T_3 = csr_write == 2'h1; // @[IDU.scala 492:72]
  wire  _conflict_es_rs1_T_4 = ~src1_is_pc | inst_type == 32'h45 | csr_write == 2'h1; // @[IDU.scala 492:59]
  wire [4:0] rs1 = inst[19:15]; // @[IDU.scala 227:16]
  wire  _conflict_es_rs1_T_6 = rs1 != 5'h0; // @[IDU.scala 492:111]
  wire  conflict_es_rs1 = (~src1_is_pc | inst_type == 32'h45 | csr_write == 2'h1) & (rs1 == io_es_rf_dst & rs1 != 5'h0
     & io_es_rf_we & io_es_valid); // @[IDU.scala 492:81]
  wire  conflict_ms_rs1 = _conflict_es_rs1_T_4 & (rs1 == io_ms_rf_dst & _conflict_es_rs1_T_6 & io_ms_rf_we & io_ms_valid
    ); // @[IDU.scala 493:81]
  wire  conflict_ws_rs1 = _conflict_es_rs1_T_4 & (rs1 == io_ws_rf_dst & _conflict_es_rs1_T_6 & io_ws_rf_we & io_ws_valid
    ); // @[IDU.scala 494:81]
  wire  src2_is_imm = 32'h45 == inst_type | (32'h43 == inst_type | (32'h44 == inst_type | (32'h42 == inst_type | 32'h40
     == inst_type))); // @[Mux.scala 81:58]
  wire  _conflict_es_rs2_T_5 = csr_write == 2'h3; // @[IDU.scala 495:92]
  wire  _conflict_es_rs2_T_6 = ~src2_is_imm | inst_type == 32'h44 | _conflict_es_rs1_T_1 | csr_write == 2'h3; // @[IDU.scala 495:81]
  wire [4:0] rs2 = csr_write[0] ? 5'h11 : inst[24:20]; // @[IDU.scala 226:15]
  wire  _conflict_es_rs2_T_8 = rs2 != 5'h0; // @[IDU.scala 495:130]
  wire  conflict_es_rs2 = (~src2_is_imm | inst_type == 32'h44 | _conflict_es_rs1_T_1 | csr_write == 2'h3) & (rs2 ==
    io_es_rf_dst & rs2 != 5'h0 & io_es_rf_we & io_es_valid); // @[IDU.scala 495:100]
  wire  conflict_ms_rs2 = _conflict_es_rs2_T_6 & (rs2 == io_ms_rf_dst & _conflict_es_rs2_T_8 & io_ms_rf_we & io_ms_valid
    ); // @[IDU.scala 496:100]
  wire  conflict_ws_rs2 = _conflict_es_rs2_T_6 & (rs2 == io_ws_rf_dst & _conflict_es_rs2_T_8 & io_ws_rf_we & io_ws_valid
    ); // @[IDU.scala 497:100]
  wire  _ds_ready_go_T_33 = conflict_es_rs2 & (io_es_fwd_ready & ~io_es_ld) | ~conflict_es_rs2 & conflict_ms_rs2 &
    io_ms_fwd_ready | ~conflict_es_rs2 & ~conflict_ms_rs2 & conflict_ws_rs2 | ~(conflict_es_rs2 | conflict_ms_rs2 |
    conflict_ws_rs2); // @[IDU.scala 150:459]
  wire  ds_ready_go = (conflict_es_rs1 & (io_es_fwd_ready & ~io_es_ld) | ~conflict_es_rs1 & conflict_ms_rs1 &
    io_ms_fwd_ready | ~conflict_es_rs1 & ~conflict_ms_rs1 & conflict_ws_rs1 | ~(conflict_es_rs1 | conflict_ms_rs1 |
    conflict_ws_rs1)) & _ds_ready_go_T_33; // @[IDU.scala 150:265]
  wire  ds_allowin = ~ds_valid | ds_ready_go & io_es_allowin; // @[IDU.scala 152:29]
  wire  _T = ds_allowin & io_fs_to_ds_valid; // @[IDU.scala 133:21]
  wire [63:0] _rdata1_T = conflict_ws_rs1 ? io_ws_fwd_res : io_rdata1; // @[IDU.scala 498:86]
  wire [63:0] _rdata1_T_1 = conflict_ms_rs1 ? io_ms_fwd_res : _rdata1_T; // @[IDU.scala 498:52]
  wire [63:0] rdata1 = conflict_es_rs1 ? io_es_fwd_res : _rdata1_T_1; // @[IDU.scala 498:18]
  wire [63:0] _br_taken_T = conflict_es_rs1 ? io_es_fwd_res : _rdata1_T_1; // @[IDU.scala 483:27]
  wire [63:0] _rdata2_T = conflict_ws_rs2 ? io_ws_fwd_res : io_rdata2; // @[IDU.scala 499:86]
  wire [63:0] _rdata2_T_1 = conflict_ms_rs2 ? io_ms_fwd_res : _rdata2_T; // @[IDU.scala 499:52]
  wire [63:0] rdata2 = conflict_es_rs2 ? io_es_fwd_res : _rdata2_T_1; // @[IDU.scala 499:18]
  wire [63:0] _br_taken_T_1 = conflict_es_rs2 ? io_es_fwd_res : _rdata2_T_1; // @[IDU.scala 483:45]
  wire  _br_taken_T_2 = $signed(_br_taken_T) != $signed(_br_taken_T_1); // @[IDU.scala 483:34]
  wire  _br_taken_T_6 = $signed(_br_taken_T) == $signed(_br_taken_T_1); // @[IDU.scala 484:34]
  wire  _br_taken_T_10 = $signed(_br_taken_T) >= $signed(_br_taken_T_1); // @[IDU.scala 485:34]
  wire  _br_taken_T_14 = $signed(_br_taken_T) < $signed(_br_taken_T_1); // @[IDU.scala 486:34]
  wire  _br_taken_T_16 = rdata1 < rdata2; // @[IDU.scala 487:28]
  wire  _br_taken_T_18 = rdata1 >= rdata2; // @[IDU.scala 488:28]
  wire  _br_taken_T_39 = 32'h30200073 == inst; // @[Lookup.scala 31:38]
  wire  _br_taken_T_42 = _src1_is_pc_T_15 ? _br_taken_T_18 : _inst_type_T_119 | _br_taken_T_39; // @[Lookup.scala 34:39]
  wire  _br_taken_T_43 = _src1_is_pc_T_13 ? _br_taken_T_16 : _br_taken_T_42; // @[Lookup.scala 34:39]
  wire  _br_taken_T_44 = _src1_is_pc_T_11 ? _br_taken_T_14 : _br_taken_T_43; // @[Lookup.scala 34:39]
  wire  _br_taken_T_45 = _src1_is_pc_T_9 ? _br_taken_T_10 : _br_taken_T_44; // @[Lookup.scala 34:39]
  wire  _br_taken_T_46 = _src1_is_pc_T_7 ? _br_taken_T_6 : _br_taken_T_45; // @[Lookup.scala 34:39]
  wire  _br_taken_T_47 = _src1_is_pc_T_5 ? _br_taken_T_2 : _br_taken_T_46; // @[Lookup.scala 34:39]
  wire  br_taken = _src1_is_pc_T_1 | (_inst_type_T_9 | _br_taken_T_47); // @[Lookup.scala 34:39]
  wire  _T_2 = ~br_taken_cancel; // @[IDU.scala 133:57]
  wire  _GEN_0 = _T & br_taken_cancel ? 1'h0 : br_taken_cancel; // @[IDU.scala 135:67 136:25 122:34]
  wire  _GEN_1 = ds_allowin & io_fs_to_ds_valid & br_taken & ~br_taken_cancel | _GEN_0; // @[IDU.scala 133:74 134:25]
  wire  _T_7 = br_taken & _T_2; // @[IDU.scala 140:19]
  wire [4:0] rd = inst[11:7]; // @[IDU.scala 228:15]
  wire  fence = 32'h100f == inst; // @[Lookup.scala 31:38]
  wire [11:0] imm_imm = inst[31:20]; // @[IDU.scala 83:23]
  wire [51:0] _imm_T_2 = imm_imm[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_3 = {_imm_T_2,imm_imm}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_1 = {inst[31],inst[19:12],inst[20],inst[30:21]}; // @[Cat.scala 31:58]
  wire [42:0] _imm_T_6 = imm_imm_1[19] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_7 = {_imm_T_6,inst[31],inst[19:12],inst[20],inst[30:21],1'h0}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_2 = inst[31:12]; // @[IDU.scala 87:23]
  wire [31:0] _imm_T_10 = imm_imm_2[19] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_12 = {_imm_T_10,imm_imm_2,12'h0}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_3 = {inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [51:0] _imm_T_15 = imm_imm_3[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_16 = {_imm_T_15,inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_4 = {inst[31],inst[7],inst[30:25],inst[11:8]}; // @[Cat.scala 31:58]
  wire [50:0] _imm_T_19 = imm_imm_4[11] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_20 = {_imm_T_19,inst[31],inst[7],inst[30:25],inst[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [63:0] _imm_T_22 = 32'h40 == inst_type ? _imm_T_3 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_24 = 32'h43 == inst_type ? _imm_T_7 : _imm_T_22; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_26 = 32'h42 == inst_type ? _imm_T_12 : _imm_T_24; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_28 = 32'h44 == inst_type ? _imm_T_16 : _imm_T_26; // @[Mux.scala 81:58]
  wire [63:0] imm = 32'h45 == inst_type ? _imm_T_20 : _imm_T_28; // @[Mux.scala 81:58]
  wire  _ALUop_T_3 = 32'h100073 == inst; // @[Lookup.scala 31:38]
  wire [6:0] _ALUop_T_118 = _inst_type_T_125 ? 7'h47 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_119 = _inst_type_T_123 ? 7'h46 : _ALUop_T_118; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_120 = _inst_type_T_121 ? 7'h3f : _ALUop_T_119; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_121 = _br_taken_T_39 ? 7'h3e : _ALUop_T_120; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_122 = _inst_type_T_119 ? 7'h3d : _ALUop_T_121; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_123 = _inst_type_T_115 ? 7'hf : _ALUop_T_122; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_124 = _inst_type_T_113 ? 7'hf : _ALUop_T_123; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_125 = _inst_type_T_111 ? 7'h1f : _ALUop_T_124; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_126 = _inst_type_T_109 ? 7'h39 : _ALUop_T_125; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_127 = _inst_type_T_107 ? 7'h38 : _ALUop_T_126; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_128 = _inst_type_T_105 ? 7'h37 : _ALUop_T_127; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_129 = _inst_type_T_103 ? 7'h34 : _ALUop_T_128; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_130 = _inst_type_T_101 ? 7'h33 : _ALUop_T_129; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_131 = _inst_type_T_99 ? 7'h32 : _ALUop_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_132 = _inst_type_T_97 ? 7'h35 : _ALUop_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_133 = _inst_type_T_95 ? 7'h31 : _ALUop_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_134 = _inst_type_T_93 ? 7'h30 : _ALUop_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_135 = _inst_type_T_91 ? 7'hb : _ALUop_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_136 = _inst_type_T_89 ? 7'h2e : _ALUop_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_137 = _inst_type_T_87 ? 7'h14 : _ALUop_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_138 = _inst_type_T_85 ? 7'h13 : _ALUop_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_139 = _inst_type_T_83 ? 7'h12 : _ALUop_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_140 = _inst_type_T_81 ? 7'h11 : _ALUop_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_141 = _inst_type_T_79 ? 7'hf : _ALUop_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_142 = _inst_type_T_77 ? 7'hf : _ALUop_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_143 = _inst_type_T_75 ? 7'hf : _ALUop_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_144 = _inst_type_T_67 ? 7'h1f : _ALUop_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_145 = _inst_type_T_65 ? 7'h1e : _ALUop_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_146 = _inst_type_T_63 ? 7'h1d : _ALUop_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_147 = _inst_type_T_61 ? 7'h1c : _ALUop_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_148 = _inst_type_T_59 ? 7'h1d : _ALUop_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_149 = _inst_type_T_57 ? 7'h1c : _ALUop_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_150 = _inst_type_T_55 ? 7'h16 : _ALUop_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_151 = _inst_type_T_53 ? 7'h38 : _ALUop_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_152 = _inst_type_T_51 ? 7'h37 : _ALUop_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_153 = _inst_type_T_49 ? 7'h16 : _ALUop_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_154 = _inst_type_T_47 ? 7'hd : _ALUop_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_155 = _inst_type_T_45 ? 7'h8 : _ALUop_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_156 = _inst_type_T_43 ? 7'h8 : _ALUop_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_157 = _inst_type_T_41 ? 7'h2e : _ALUop_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_158 = _inst_type_T_39 ? 7'hb : _ALUop_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_159 = _inst_type_T_37 ? 7'hf : _ALUop_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_160 = _inst_type_T_35 ? 7'hf : _ALUop_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_161 = _inst_type_T_33 ? 7'hf : _ALUop_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_162 = _inst_type_T_31 ? 7'h15 : _ALUop_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_163 = _inst_type_T_29 ? 7'hf : _ALUop_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_164 = _inst_type_T_27 ? 7'hc : _ALUop_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_165 = _inst_type_T_25 ? 7'hf : _ALUop_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_166 = _inst_type_T_19 ? 7'he : _ALUop_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_167 = _inst_type_T_17 ? 7'hc : _ALUop_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_168 = _inst_type_T_15 ? 7'hf : _ALUop_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_169 = _inst_type_T_13 ? 7'h1e : _ALUop_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_170 = _inst_type_T_11 ? 7'hf : _ALUop_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_171 = _inst_type_T_9 ? 7'h6 : _ALUop_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_172 = _src1_is_pc_T_1 ? 7'h5 : _ALUop_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_173 = _inst_type_T_5 ? 7'h4 : _ALUop_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_174 = _src1_is_pc_T_3 ? 7'hf : _ALUop_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_175 = _ALUop_T_3 ? 7'h2 : _ALUop_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _ALUop_T_176 = _inst_type_T_1 ? 7'hf : _ALUop_T_175; // @[Lookup.scala 34:39]
  wire  _reg_write_T_28 = fence ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _reg_write_T_29 = _br_taken_T_39 ? 1'h0 : _reg_write_T_28; // @[Lookup.scala 34:39]
  wire  _reg_write_T_30 = _inst_type_T_119 ? 1'h0 : _reg_write_T_29; // @[Lookup.scala 34:39]
  wire  _reg_write_T_31 = _src1_is_pc_T_15 ? 1'h0 : _reg_write_T_30; // @[Lookup.scala 34:39]
  wire  _reg_write_T_32 = _src1_is_pc_T_13 ? 1'h0 : _reg_write_T_31; // @[Lookup.scala 34:39]
  wire  _reg_write_T_33 = _src1_is_pc_T_11 ? 1'h0 : _reg_write_T_32; // @[Lookup.scala 34:39]
  wire  _reg_write_T_34 = _src1_is_pc_T_9 ? 1'h0 : _reg_write_T_33; // @[Lookup.scala 34:39]
  wire  _reg_write_T_35 = _src1_is_pc_T_7 ? 1'h0 : _reg_write_T_34; // @[Lookup.scala 34:39]
  wire  _reg_write_T_36 = _src1_is_pc_T_5 ? 1'h0 : _reg_write_T_35; // @[Lookup.scala 34:39]
  wire  _reg_write_T_37 = _inst_type_T_75 ? 1'h0 : _reg_write_T_36; // @[Lookup.scala 34:39]
  wire  _reg_write_T_38 = _inst_type_T_37 ? 1'h0 : _reg_write_T_37; // @[Lookup.scala 34:39]
  wire  _reg_write_T_39 = _inst_type_T_35 ? 1'h0 : _reg_write_T_38; // @[Lookup.scala 34:39]
  wire  _reg_write_T_40 = _inst_type_T_11 ? 1'h0 : _reg_write_T_39; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_14 = _inst_type_T_79 ? 3'h7 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_15 = _inst_type_T_115 ? 3'h6 : _load_type_T_14; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_16 = _inst_type_T_77 ? 3'h5 : _load_type_T_15; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_17 = _inst_type_T_113 ? 3'h4 : _load_type_T_16; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_18 = _inst_type_T_33 ? 3'h3 : _load_type_T_17; // @[Lookup.scala 34:39]
  wire [2:0] _load_type_T_19 = _inst_type_T_25 ? 3'h2 : _load_type_T_18; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_8 = _inst_type_T_75 ? 4'hf : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_9 = _inst_type_T_37 ? 4'h1 : _Wmask_T_8; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_10 = _inst_type_T_35 ? 4'h3 : _Wmask_T_9; // @[Lookup.scala 34:39]
  wire [1:0] _csr_index_T_6 = 12'h300 == imm[11:0] ? 2'h2 : {{1'd0}, 12'h341 == imm[11:0]}; // @[Mux.scala 81:58]
  wire [1:0] csr_index = 12'h342 == imm[11:0] ? 2'h3 : _csr_index_T_6; // @[Mux.scala 81:58]
  wire [63:0] _csr_wdata_T = rdata1 | csr_reg_io_rdata; // @[IDU.scala 458:26]
  wire [63:0] _csr_wdata_T_1 = ~csr_reg_io_rdata; // @[IDU.scala 459:29]
  wire [63:0] _csr_wdata_T_2 = rdata1 & _csr_wdata_T_1; // @[IDU.scala 459:26]
  wire [63:0] _csr_wdata_T_9 = _inst_type_T_125 ? _csr_wdata_T_2 : 64'h0; // @[Lookup.scala 34:39]
  wire [63:0] _csr_wdata_T_10 = _inst_type_T_123 ? _csr_wdata_T : _csr_wdata_T_9; // @[Lookup.scala 34:39]
  wire [63:0] csr_wdata = _inst_type_T_121 ? rdata1 : _csr_wdata_T_10; // @[Lookup.scala 34:39]
  wire [31:0] ALUop = {{25'd0}, _ALUop_T_176}; // @[IDU.scala 311:11 65:21]
  wire [1:0] _T_17 = ALUop == 32'h3e ? 2'h1 : csr_index; // @[IDU.scala 462:48]
  wire [1:0] _T_24 = _conflict_es_rs1_T_3 ? csr_index : 2'h0; // @[IDU.scala 464:46]
  wire [63:0] _T_28 = _conflict_es_rs1_T_3 ? csr_wdata : 64'h0; // @[IDU.scala 465:48]
  wire [63:0] src1 = src1_is_pc ? ds_pc : rdata1; // @[IDU.scala 471:16]
  wire [63:0] src2 = src2_is_imm ? imm : rdata2; // @[IDU.scala 472:16]
  wire [63:0] _br_target_T_1 = src1 + src2; // @[IDU.scala 475:35]
  wire [63:0] _br_target_T_4 = _br_target_T_1 & 64'hfffffffffffffffe; // @[IDU.scala 476:31]
  wire [63:0] _br_target_T_6 = csr_reg_io_rdata + 64'h4; // @[IDU.scala 478:28]
  wire [63:0] _br_target_T_13 = _br_taken_T_39 ? _br_target_T_6 : _br_target_T_1; // @[Lookup.scala 34:39]
  wire [63:0] _br_target_T_14 = _inst_type_T_119 ? csr_reg_io_rdata : _br_target_T_13; // @[Lookup.scala 34:39]
  wire [31:0] _io_store_data_T_11 = _inst_type_T_75 ? rdata2[31:0] : 32'h0; // @[Lookup.scala 34:39]
  wire [31:0] _io_store_data_T_12 = _inst_type_T_37 ? {{24'd0}, rdata2[7:0]} : _io_store_data_T_11; // @[Lookup.scala 34:39]
  wire [31:0] _io_store_data_T_13 = _inst_type_T_35 ? {{16'd0}, rdata2[15:0]} : _io_store_data_T_12; // @[Lookup.scala 34:39]
  csr_reg csr_reg ( // @[IDU.scala 449:21]
    .clock(csr_reg_clock),
    .io_wen1(csr_reg_io_wen1),
    .io_wen2(csr_reg_io_wen2),
    .io_waddr1(csr_reg_io_waddr1),
    .io_wdata1(csr_reg_io_wdata1),
    .io_wdata2(csr_reg_io_wdata2),
    .io_raddr(csr_reg_io_raddr),
    .io_rdata(csr_reg_io_rdata)
  );
  assign io_ds_to_es_valid = ds_valid & ds_ready_go; // @[IDU.scala 151:32]
  assign io_br_taken = br_taken & ds_ready_go & _T_2; // @[IDU.scala 503:44]
  assign io_br_target = _inst_type_T_9 ? _br_target_T_4 : _br_target_T_14; // @[Lookup.scala 34:39]
  assign io_ds_allowin = ~ds_valid | ds_ready_go & io_es_allowin; // @[IDU.scala 152:29]
  assign io_ds_ready_go = (conflict_es_rs1 & (io_es_fwd_ready & ~io_es_ld) | ~conflict_es_rs1 & conflict_ms_rs1 &
    io_ms_fwd_ready | ~conflict_es_rs1 & ~conflict_ms_rs1 & conflict_ws_rs1 | ~(conflict_es_rs1 | conflict_ms_rs1 |
    conflict_ws_rs1)) & _ds_ready_go_T_33; // @[IDU.scala 150:265]
  assign io_fence = 32'h100f == inst; // @[Lookup.scala 31:38]
  assign io_raddr1 = inst[19:15]; // @[IDU.scala 227:16]
  assign io_raddr2 = csr_write[0] ? 5'h11 : inst[24:20]; // @[IDU.scala 226:15]
  assign io_to_es_pc = ds_pc; // @[IDU.scala 526:17]
  assign io_ALUop = {{25'd0}, _ALUop_T_176}; // @[IDU.scala 311:11 65:21]
  assign io_src1 = csr_write[0] ? csr_reg_io_rdata : src1; // @[IDU.scala 515:19]
  assign io_src2 = src2_is_imm ? imm : rdata2; // @[IDU.scala 472:16]
  assign io_rf_dst = inst[11:7]; // @[IDU.scala 228:15]
  assign io_store_data = _inst_type_T_11 ? rdata2 : {{32'd0}, _io_store_data_T_13}; // @[Lookup.scala 34:39]
  assign io_ctrl_sign_reg_write = _ALUop_T_3 ? 1'h0 : _reg_write_T_40; // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Writemem_en = 32'h44 == inst_type; // @[Mux.scala 81:61]
  assign io_ctrl_sign_Readmem_en = _inst_type_T_25 | (_inst_type_T_15 | (_inst_type_T_113 | (_inst_type_T_77 | (
    _inst_type_T_79 | (_inst_type_T_115 | _inst_type_T_33))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Wmask = _inst_type_T_11 ? 8'hff : {{4'd0}, _Wmask_T_10}; // @[Lookup.scala 34:39]
  assign io_load_type = _inst_type_T_15 ? 3'h1 : _load_type_T_19; // @[Lookup.scala 34:39]
  assign io_ds_valid = ds_valid; // @[IDU.scala 528:17]
  assign csr_reg_clock = clock;
  assign csr_reg_io_wen1 = csr_write[0] & ds_valid; // @[IDU.scala 463:38]
  assign csr_reg_io_wen2 = csr_write[1] & ds_valid; // @[IDU.scala 466:38]
  assign csr_reg_io_waddr1 = _conflict_es_rs2_T_5 ? 2'h1 : _T_24; // @[IDU.scala 464:22]
  assign csr_reg_io_wdata1 = _conflict_es_rs2_T_5 ? ds_pc : _T_28; // @[IDU.scala 465:22]
  assign csr_reg_io_wdata2 = conflict_es_rs2 ? io_es_fwd_res : _rdata2_T_1; // @[IDU.scala 499:18]
  assign csr_reg_io_raddr = csr_write[1] ? 2'h0 : _T_17; // @[IDU.scala 462:21]
  always @(posedge clock) begin
    if (reset) begin // @[IDU.scala 112:27]
      ds_valid <= 1'h0; // @[IDU.scala 112:27]
    end else if (br_taken & _T_2 & ds_allowin) begin // @[IDU.scala 140:53]
      ds_valid <= 1'h0; // @[IDU.scala 141:18]
    end else if (ds_allowin) begin // @[IDU.scala 142:27]
      ds_valid <= io_fs_to_ds_valid; // @[IDU.scala 143:18]
    end
    if (reset) begin // @[IDU.scala 116:24]
      ds_pc <= 64'h0; // @[IDU.scala 116:24]
    end else if (io_fs_to_ds_valid & ds_allowin & ~_T_7) begin // @[IDU.scala 145:75]
      ds_pc <= io_pc; // @[IDU.scala 146:15]
    end
    if (reset) begin // @[IDU.scala 118:23]
      inst <= 32'h0; // @[IDU.scala 118:23]
    end else if (io_fs_to_ds_valid & ds_allowin & ~_T_7) begin // @[IDU.scala 145:75]
      inst <= io_from_fs_inst; // @[IDU.scala 147:14]
    end
    if (reset) begin // @[IDU.scala 122:34]
      br_taken_cancel <= 1'h0; // @[IDU.scala 122:34]
    end else begin
      br_taken_cancel <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ds_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  ds_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  br_taken_cancel = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module partial_product(
  input  [2:0]  io_y,
  input  [63:0] io_x,
  output        io_c,
  output [63:0] io_p
);
  wire [64:0] _io_p_T = {io_x, 1'h0}; // @[Mul.scala 24:18]
  wire [64:0] _io_p_T_2 = ~_io_p_T; // @[Mul.scala 25:12]
  wire [63:0] _io_p_T_3 = ~io_x; // @[Mul.scala 26:12]
  wire [63:0] _io_p_T_6 = 3'h1 == io_y ? io_x : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_p_T_8 = 3'h2 == io_y ? io_x : _io_p_T_6; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_10 = 3'h3 == io_y ? _io_p_T : {{1'd0}, _io_p_T_8}; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_12 = 3'h4 == io_y ? _io_p_T_2 : _io_p_T_10; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_14 = 3'h5 == io_y ? {{1'd0}, _io_p_T_3} : _io_p_T_12; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_16 = 3'h6 == io_y ? {{1'd0}, _io_p_T_3} : _io_p_T_14; // @[Mux.scala 81:58]
  wire [64:0] _io_p_T_18 = 3'h7 == io_y ? 65'h0 : _io_p_T_16; // @[Mux.scala 81:58]
  assign io_c = 3'h6 == io_y | (3'h5 == io_y | 3'h4 == io_y); // @[Mux.scala 81:58]
  assign io_p = _io_p_T_18[63:0]; // @[Mul.scala 20:8]
endmodule
module Mul(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input         io_mulw,
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output        io_out_valid,
  input         io_out_ready,
  output [31:0] io_result_hi,
  output [31:0] io_result_lo
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [95:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] booth_partial_io_y; // @[Mul.scala 72:31]
  wire [63:0] booth_partial_io_x; // @[Mul.scala 72:31]
  wire  booth_partial_io_c; // @[Mul.scala 72:31]
  wire [63:0] booth_partial_io_p; // @[Mul.scala 72:31]
  wire  sign = io_multiplicand[63] ^ io_multiplier[63]; // @[Mul.scala 52:33]
  reg [63:0] res; // @[Mul.scala 54:22]
  reg [1:0] state; // @[Mul.scala 56:24]
  reg [127:0] src1; // @[Mul.scala 58:23]
  reg [64:0] src2; // @[Mul.scala 59:23]
  wire [31:0] _src1_32_T_2 = io_multiplicand[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _src1_32_T_4 = {_src1_32_T_2,io_multiplicand[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] src1_32 = io_mulw ? _src1_32_T_4 : io_multiplicand; // @[Mul.scala 66:19]
  wire [31:0] _src2_32_T_2 = io_multiplier[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _src2_32_T_4 = {_src2_32_T_2,io_multiplier[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] src2_32 = io_mulw ? _src2_32_T_4 : io_multiplier; // @[Mul.scala 67:19]
  wire [63:0] _real_cand_T_5 = src1_32[63] ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 74:12]
  wire [127:0] real_cand = {_real_cand_T_5,src1_32}; // @[Cat.scala 31:58]
  wire [64:0] _real_er_T = {src2_32,1'h0}; // @[Cat.scala 31:58]
  wire [127:0] _GEN_1 = io_mul_valid ? real_cand : src1; // @[Mul.scala 78:44 80:22 58:23]
  wire [63:0] real_er = _real_er_T[63:0]; // @[Mul.scala 62:23 70:13]
  wire  _T_4 = src2 != 65'h0; // @[Mul.scala 89:26]
  wire [63:0] _res_T_1 = res + booth_partial_io_p; // @[Mul.scala 90:32]
  wire [63:0] _GEN_21 = {{63'd0}, booth_partial_io_c}; // @[Mul.scala 90:53]
  wire [63:0] _res_T_3 = _res_T_1 + _GEN_21; // @[Mul.scala 90:53]
  wire [129:0] _src1_T = {src1, 2'h0}; // @[Mul.scala 92:34]
  wire [1:0] _GEN_4 = io_out_ready ? 2'h0 : state; // @[Mul.scala 56:24 94:39 95:31]
  wire [129:0] _GEN_7 = src2 != 65'h0 ? _src1_T : {{2'd0}, src1}; // @[Mul.scala 58:23 89:33 92:26]
  wire [129:0] _GEN_16 = 2'h1 == state ? _GEN_7 : {{2'd0}, src1}; // @[Mul.scala 76:18 58:23]
  wire [129:0] _GEN_18 = 2'h0 == state ? {{2'd0}, _GEN_1} : _GEN_16; // @[Mul.scala 76:18]
  wire [31:0] _io_result_hi_T_1 = {sign,res[62:32]}; // @[Cat.scala 31:58]
  wire  _GEN_22 = _T_4 ? 1'h0 : 1'h1; // @[Mul.scala 108:35 110:26 116:26]
  wire [31:0] _GEN_23 = _T_4 ? 32'h0 : _io_result_hi_T_1; // @[Mul.scala 108:35 111:26 114:26]
  wire [31:0] _GEN_24 = _T_4 ? 32'h0 : res[31:0]; // @[Mul.scala 108:35 112:26 115:26]
  wire  _GEN_26 = state == 2'h1 & _GEN_22; // @[Mul.scala 107:33 121:22]
  wire [31:0] _GEN_27 = state == 2'h1 ? _GEN_23 : 32'h0; // @[Mul.scala 107:33 122:22]
  wire [31:0] _GEN_28 = state == 2'h1 ? _GEN_24 : 32'h0; // @[Mul.scala 107:33 123:22]
  wire [129:0] _GEN_25 = reset ? 130'h0 : _GEN_18; // @[Mul.scala 58:{23,23}]
  partial_product booth_partial ( // @[Mul.scala 72:31]
    .io_y(booth_partial_io_y),
    .io_x(booth_partial_io_x),
    .io_c(booth_partial_io_c),
    .io_p(booth_partial_io_p)
  );
  assign io_out_valid = state == 2'h0 ? 1'h0 : _GEN_26; // @[Mul.scala 102:23 104:22]
  assign io_result_hi = state == 2'h0 ? 32'h0 : _GEN_27; // @[Mul.scala 102:23 105:22]
  assign io_result_lo = state == 2'h0 ? 32'h0 : _GEN_28; // @[Mul.scala 102:23 106:22]
  assign booth_partial_io_y = src2[2:0]; // @[Mul.scala 73:31]
  assign booth_partial_io_x = src1[63:0]; // @[Mul.scala 74:24]
  always @(posedge clock) begin
    if (reset) begin // @[Mul.scala 54:22]
      res <= 64'h0; // @[Mul.scala 54:22]
    end else if (2'h0 == state) begin // @[Mul.scala 76:18]
      if (io_mul_valid) begin // @[Mul.scala 78:44]
        res <= 64'h0; // @[Mul.scala 82:21]
      end
    end else if (2'h1 == state) begin // @[Mul.scala 76:18]
      if (src2 != 65'h0) begin // @[Mul.scala 89:33]
        res <= _res_T_3; // @[Mul.scala 90:25]
      end
    end
    if (reset) begin // @[Mul.scala 56:24]
      state <= 2'h0; // @[Mul.scala 56:24]
    end else if (2'h0 == state) begin // @[Mul.scala 76:18]
      if (io_mul_valid) begin // @[Mul.scala 78:44]
        state <= 2'h1; // @[Mul.scala 79:23]
      end
    end else if (2'h1 == state) begin // @[Mul.scala 76:18]
      if (!(src2 != 65'h0)) begin // @[Mul.scala 89:33]
        state <= _GEN_4;
      end
    end
    src1 <= _GEN_25[127:0]; // @[Mul.scala 58:{23,23}]
    if (reset) begin // @[Mul.scala 59:23]
      src2 <= 65'h0; // @[Mul.scala 59:23]
    end else if (2'h0 == state) begin // @[Mul.scala 76:18]
      if (io_mul_valid) begin // @[Mul.scala 78:44]
        src2 <= {{1'd0}, real_er}; // @[Mul.scala 81:22]
      end
    end else if (2'h1 == state) begin // @[Mul.scala 76:18]
      if (src2 != 65'h0) begin // @[Mul.scala 89:33]
        src2 <= {{2'd0}, src2[64:2]}; // @[Mul.scala 91:26]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  res = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  _RAND_2 = {4{`RANDOM}};
  src1 = _RAND_2[127:0];
  _RAND_3 = {3{`RANDOM}};
  src2 = _RAND_3[64:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Div(
  input         clock,
  input         reset,
  input  [63:0] io_dividend,
  input  [63:0] io_divisor,
  input         io_div_valid,
  input         io_divw,
  input         io_div_signed,
  output        io_out_valid,
  input         io_out_ready,
  output [63:0] io_quotient,
  output [63:0] io_remainder
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  dend_neg = io_divw ? io_dividend[31] : io_dividend[63]; // @[Div.scala 26:20]
  wire  sor_neg = io_divw ? io_divisor[31] : io_divisor[63]; // @[Div.scala 27:19]
  wire  quotient_neg = dend_neg & ~sor_neg | ~dend_neg & sor_neg; // @[Div.scala 28:43]
  wire [31:0] _src1_32_s_T_2 = io_dividend[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _src1_32_s_T_4 = {_src1_32_s_T_2,io_dividend[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] src1_32_s = io_divw ? _src1_32_s_T_4 : io_dividend; // @[Div.scala 36:21]
  wire [31:0] _src2_32_s_T_2 = io_divisor[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _src2_32_s_T_4 = {_src2_32_s_T_2,io_divisor[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] src2_32_s = io_divw ? _src2_32_s_T_4 : io_divisor; // @[Div.scala 37:21]
  wire [63:0] src1_32 = io_divw ? {{32'd0}, io_dividend[31:0]} : io_dividend; // @[Div.scala 38:19]
  wire [63:0] src2_32 = io_divw ? {{32'd0}, io_divisor[31:0]} : io_divisor; // @[Div.scala 39:19]
  wire [63:0] _real_cand_T_2 = ~src1_32_s; // @[Div.scala 43:61]
  wire [63:0] _real_cand_T_4 = _real_cand_T_2 + 64'h1; // @[Div.scala 43:71]
  wire [63:0] _real_cand_T_5 = dend_neg ? _real_cand_T_4 : src1_32_s; // @[Div.scala 43:45]
  wire [63:0] real_cand = io_div_signed ? _real_cand_T_5 : src1_32; // @[Div.scala 43:21]
  wire [63:0] _real_er_T_2 = ~src2_32_s; // @[Div.scala 44:58]
  wire [63:0] _real_er_T_4 = _real_er_T_2 + 64'h1; // @[Div.scala 44:68]
  wire [63:0] _real_er_T_5 = sor_neg ? _real_er_T_4 : src2_32_s; // @[Div.scala 44:43]
  wire [63:0] real_er = io_div_signed ? _real_er_T_5 : src2_32; // @[Div.scala 44:19]
  wire [95:0] _src1_T_1 = {32'h0,real_cand}; // @[Cat.scala 31:58]
  wire [64:0] src2 = {1'h0,real_er}; // @[Cat.scala 31:58]
  reg [127:0] div_cand; // @[Div.scala 51:27]
  reg  div_start; // @[Div.scala 52:28]
  reg [63:0] quotient; // @[Div.scala 54:27]
  reg [31:0] step_num; // @[Div.scala 56:27]
  wire  _GEN_0 = io_out_ready ? 1'h0 : div_start; // @[Div.scala 69:33 70:23 52:28]
  wire  _GEN_1 = io_div_valid & ~div_start | _GEN_0; // @[Div.scala 63:41 64:23]
  wire [127:0] src1 = {{32'd0}, _src1_T_1}; // @[Div.scala 46:20 48:10]
  wire [127:0] _GEN_2 = io_div_valid & ~div_start ? src1 : div_cand; // @[Div.scala 63:41 65:22 51:27]
  wire [63:0] _GEN_3 = io_div_valid & ~div_start ? 64'h0 : quotient; // @[Div.scala 63:41 66:22 54:27]
  wire [31:0] _GEN_4 = io_div_valid & ~div_start ? 32'h40 : step_num; // @[Div.scala 63:41 68:22 56:27]
  wire [64:0] sub_res = div_cand[127:63] - src2; // @[Div.scala 78:41]
  wire [64:0] _quotient_T_2 = {quotient, 1'h0}; // @[Div.scala 80:57]
  wire [64:0] _quotient_T_4 = _quotient_T_2 | 65'h1; // @[Div.scala 80:81]
  wire [64:0] _quotient_T_5 = sub_res[64] ? _quotient_T_2 : _quotient_T_4; // @[Div.scala 80:28]
  wire [127:0] update_cand = {sub_res, 63'h0}; // @[Div.scala 81:36]
  wire [127:0] _new_cand_T_2 = div_cand & 128'h7fffffffffffffff; // @[Div.scala 82:68]
  wire [127:0] _new_cand_T_3 = _new_cand_T_2 | update_cand; // @[Div.scala 82:93]
  wire [127:0] new_cand = sub_res[64] ? div_cand : _new_cand_T_3; // @[Div.scala 82:28]
  wire [128:0] _div_cand_T = {new_cand, 1'h0}; // @[Div.scala 83:34]
  wire [31:0] _step_num_T_1 = step_num - 32'h1; // @[Div.scala 84:34]
  wire [63:0] _io_remainder_T_3 = ~div_cand[127:64]; // @[Div.scala 89:77]
  wire [63:0] _io_remainder_T_5 = _io_remainder_T_3 + 64'h1; // @[Div.scala 89:94]
  wire [63:0] _io_remainder_T_7 = dend_neg ? _io_remainder_T_5 : div_cand[127:64]; // @[Div.scala 89:56]
  wire [63:0] _io_remainder_T_9 = io_div_signed ? _io_remainder_T_7 : div_cand[127:64]; // @[Div.scala 89:32]
  wire [63:0] _io_quotient_T_2 = ~quotient; // @[Div.scala 91:75]
  wire [63:0] _io_quotient_T_4 = _io_quotient_T_2 + 64'h1; // @[Div.scala 91:84]
  wire [63:0] _io_quotient_T_5 = quotient_neg ? _io_quotient_T_4 : quotient; // @[Div.scala 91:55]
  wire [63:0] _io_quotient_T_6 = io_div_signed ? _io_quotient_T_5 : quotient; // @[Div.scala 91:31]
  wire [64:0] _GEN_9 = $signed(step_num) > 32'sh0 ? _quotient_T_5 : {{1'd0}, _GEN_3}; // @[Div.scala 74:36 80:22]
  wire [128:0] _GEN_10 = $signed(step_num) > 32'sh0 ? _div_cand_T : {{1'd0}, _GEN_2}; // @[Div.scala 74:36 83:22]
  wire [63:0] _GEN_12 = $signed(step_num) > 32'sh0 ? 64'h0 : _io_remainder_T_9; // @[Div.scala 74:36 85:26 89:26]
  wire  _GEN_13 = $signed(step_num) > 32'sh0 ? 1'h0 : 1'h1; // @[Div.scala 74:36 86:26 90:26]
  wire [63:0] _GEN_14 = $signed(step_num) > 32'sh0 ? 64'h0 : _io_quotient_T_6; // @[Div.scala 74:36 87:25 91:25]
  wire [64:0] _GEN_15 = div_start ? _GEN_9 : {{1'd0}, _GEN_3}; // @[Div.scala 73:20]
  wire [128:0] _GEN_16 = div_start ? _GEN_10 : {{1'd0}, _GEN_2}; // @[Div.scala 73:20]
  wire [128:0] _GEN_21 = reset ? 129'h0 : _GEN_16; // @[Div.scala 51:{27,27}]
  wire [64:0] _GEN_22 = reset ? 65'h0 : _GEN_15; // @[Div.scala 54:{27,27}]
  assign io_out_valid = div_start & _GEN_13; // @[Div.scala 73:20 95:22]
  assign io_quotient = div_start ? _GEN_14 : 64'h0; // @[Div.scala 73:20 96:21]
  assign io_remainder = div_start ? _GEN_12 : 64'h0; // @[Div.scala 73:20 94:22]
  always @(posedge clock) begin
    div_cand <= _GEN_21[127:0]; // @[Div.scala 51:{27,27}]
    if (reset) begin // @[Div.scala 52:28]
      div_start <= 1'h0; // @[Div.scala 52:28]
    end else begin
      div_start <= _GEN_1;
    end
    quotient <= _GEN_22[63:0]; // @[Div.scala 54:{27,27}]
    if (reset) begin // @[Div.scala 56:27]
      step_num <= 32'h0; // @[Div.scala 56:27]
    end else if (div_start) begin // @[Div.scala 73:20]
      if ($signed(step_num) > 32'sh0) begin // @[Div.scala 74:36]
        step_num <= _step_num_T_1; // @[Div.scala 84:22]
      end else begin
        step_num <= _GEN_4;
      end
    end else begin
      step_num <= _GEN_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  div_cand = _RAND_0[127:0];
  _RAND_1 = {1{`RANDOM}};
  div_start = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  quotient = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  step_num = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [63:0] io_src1_value,
  input  [63:0] io_src2_value,
  input  [31:0] io_ALUop,
  input         io_src_valid,
  output        io_alu_busy,
  input         io_res_ready,
  output [63:0] io_alu_res
);
  wire  Mul_clock; // @[ALU.scala 61:28]
  wire  Mul_reset; // @[ALU.scala 61:28]
  wire  Mul_io_mul_valid; // @[ALU.scala 61:28]
  wire  Mul_io_mulw; // @[ALU.scala 61:28]
  wire [63:0] Mul_io_multiplicand; // @[ALU.scala 61:28]
  wire [63:0] Mul_io_multiplier; // @[ALU.scala 61:28]
  wire  Mul_io_out_valid; // @[ALU.scala 61:28]
  wire  Mul_io_out_ready; // @[ALU.scala 61:28]
  wire [31:0] Mul_io_result_hi; // @[ALU.scala 61:28]
  wire [31:0] Mul_io_result_lo; // @[ALU.scala 61:28]
  wire  Div_clock; // @[ALU.scala 62:28]
  wire  Div_reset; // @[ALU.scala 62:28]
  wire [63:0] Div_io_dividend; // @[ALU.scala 62:28]
  wire [63:0] Div_io_divisor; // @[ALU.scala 62:28]
  wire  Div_io_div_valid; // @[ALU.scala 62:28]
  wire  Div_io_divw; // @[ALU.scala 62:28]
  wire  Div_io_div_signed; // @[ALU.scala 62:28]
  wire  Div_io_out_valid; // @[ALU.scala 62:28]
  wire  Div_io_out_ready; // @[ALU.scala 62:28]
  wire [63:0] Div_io_quotient; // @[ALU.scala 62:28]
  wire [63:0] Div_io_remainder; // @[ALU.scala 62:28]
  wire  mul_valid = 32'h12 == io_ALUop | 32'h11 == io_ALUop; // @[Mux.scala 81:58]
  wire  div_valid = 32'h32 == io_ALUop | (32'h14 == io_ALUop | (32'h33 == io_ALUop | (32'h34 == io_ALUop | (32'h35 ==
    io_ALUop | (32'h13 == io_ALUop | (32'h30 == io_ALUop | 32'h31 == io_ALUop)))))); // @[Mux.scala 81:58]
  wire [63:0] add_res = io_src1_value + io_src2_value; // @[ALU.scala 80:30]
  wire [63:0] sub_res = io_src1_value - io_src2_value; // @[ALU.scala 81:30]
  wire [63:0] sra_res = $signed(io_src1_value) >>> io_src2_value[5:0]; // @[ALU.scala 82:60]
  wire [63:0] srl_res = io_src1_value >> io_src2_value[5:0]; // @[ALU.scala 83:30]
  wire [126:0] _GEN_0 = {{63'd0}, io_src1_value}; // @[ALU.scala 84:30]
  wire [126:0] sll_res = _GEN_0 << io_src2_value[5:0]; // @[ALU.scala 84:30]
  wire [31:0] _sraw_res_T_1 = io_src1_value[31:0]; // @[ALU.scala 85:43]
  wire [31:0] sraw_res = $signed(_sraw_res_T_1) >>> io_src2_value[4:0]; // @[ALU.scala 85:46]
  wire [31:0] srlw_res = io_src1_value[31:0] >> io_src2_value[4:0]; // @[ALU.scala 86:37]
  wire [62:0] _GEN_1 = {{31'd0}, io_src1_value[31:0]}; // @[ALU.scala 87:37]
  wire [62:0] sllw_res = _GEN_1 << io_src2_value[4:0]; // @[ALU.scala 87:37]
  wire [63:0] or_res = io_src1_value | io_src2_value; // @[ALU.scala 88:29]
  wire [63:0] xor_res = io_src1_value ^ io_src2_value; // @[ALU.scala 89:30]
  wire [63:0] and_res = io_src1_value & io_src2_value; // @[ALU.scala 90:30]
  wire [63:0] mlu_res = {Mul_io_result_hi,Mul_io_result_lo}; // @[Cat.scala 31:58]
  wire [31:0] divw_res = Div_io_quotient[31:0]; // @[ALU.scala 93:39]
  wire [31:0] remw_res = Div_io_remainder[31:0]; // @[ALU.scala 95:40]
  wire [63:0] _alu_res_T_1 = io_src1_value + 64'h4; // @[ALU.scala 118:29]
  wire  _alu_res_T_4 = io_src1_value < io_src2_value; // @[ALU.scala 121:33]
  wire  _alu_res_T_8 = $signed(io_src1_value) < $signed(io_src2_value); // @[ALU.scala 123:41]
  wire [31:0] _alu_res_T_12 = add_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_14 = {_alu_res_T_12,add_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_17 = sub_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_19 = {_alu_res_T_17,sub_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_22 = sllw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_24 = {_alu_res_T_22,sllw_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_27 = sraw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _alu_res_T_28 = $signed(_sraw_res_T_1) >>> io_src2_value[4:0]; // @[ALU.scala 142:55]
  wire [63:0] _alu_res_T_29 = {_alu_res_T_27,_alu_res_T_28}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_32 = srlw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_34 = {_alu_res_T_32,srlw_res}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_37 = Mul_io_result_lo[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_38 = {_alu_res_T_37,Mul_io_result_lo}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_41 = divw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_42 = {_alu_res_T_41,divw_res}; // @[Cat.scala 31:58]
  wire [31:0] _alu_res_T_49 = remw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_res_T_50 = {_alu_res_T_49,remw_res}; // @[Cat.scala 31:58]
  wire [63:0] _alu_res_T_56 = 32'hf == io_ALUop ? add_res : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_58 = 32'h4 == io_ALUop ? io_src2_value : _alu_res_T_56; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_60 = 32'h5 == io_ALUop ? _alu_res_T_1 : _alu_res_T_58; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_62 = 32'h6 == io_ALUop ? _alu_res_T_1 : _alu_res_T_60; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_64 = 32'h1e == io_ALUop ? {{63'd0}, _alu_res_T_4} : _alu_res_T_62; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_66 = 32'h1f == io_ALUop ? {{63'd0}, _alu_res_T_8} : _alu_res_T_64; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_68 = 32'hc == io_ALUop ? _alu_res_T_14 : _alu_res_T_66; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_70 = 32'he == io_ALUop ? sub_res : _alu_res_T_68; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_72 = 32'h15 == io_ALUop ? sra_res : _alu_res_T_70; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_74 = 32'hb == io_ALUop ? or_res : _alu_res_T_72; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_76 = 32'h2e == io_ALUop ? xor_res : _alu_res_T_74; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_78 = 32'h8 == io_ALUop ? and_res : _alu_res_T_76; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_80 = 32'hd == io_ALUop ? _alu_res_T_19 : _alu_res_T_78; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_82 = 32'h16 == io_ALUop ? _alu_res_T_24 : _alu_res_T_80; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_84 = 32'h1c == io_ALUop ? _alu_res_T_29 : _alu_res_T_82; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_86 = 32'h1d == io_ALUop ? _alu_res_T_34 : _alu_res_T_84; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_88 = 32'h11 == io_ALUop ? mlu_res : _alu_res_T_86; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_90 = 32'h12 == io_ALUop ? _alu_res_T_38 : _alu_res_T_88; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_92 = 32'h13 == io_ALUop ? _alu_res_T_42 : _alu_res_T_90; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_94 = 32'h30 == io_ALUop ? Div_io_quotient : _alu_res_T_92; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_96 = 32'h31 == io_ALUop ? Div_io_quotient : _alu_res_T_94; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_98 = 32'h35 == io_ALUop ? _alu_res_T_42 : _alu_res_T_96; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_100 = 32'h14 == io_ALUop ? _alu_res_T_50 : _alu_res_T_98; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_102 = 32'h32 == io_ALUop ? _alu_res_T_50 : _alu_res_T_100; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_104 = 32'h33 == io_ALUop ? Div_io_remainder : _alu_res_T_102; // @[Mux.scala 81:58]
  wire [63:0] _alu_res_T_106 = 32'h34 == io_ALUop ? Div_io_remainder : _alu_res_T_104; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_108 = 32'h37 == io_ALUop ? sll_res : {{63'd0}, _alu_res_T_106}; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_110 = 32'h39 == io_ALUop ? {{63'd0}, sra_res} : _alu_res_T_108; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_112 = 32'h38 == io_ALUop ? {{63'd0}, srl_res} : _alu_res_T_110; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_114 = 32'h3f == io_ALUop ? {{63'd0}, io_src1_value} : _alu_res_T_112; // @[Mux.scala 81:58]
  wire [126:0] _alu_res_T_116 = 32'h46 == io_ALUop ? {{63'd0}, io_src1_value} : _alu_res_T_114; // @[Mux.scala 81:58]
  wire [126:0] alu_res = 32'h47 == io_ALUop ? {{63'd0}, io_src1_value} : _alu_res_T_116; // @[Mux.scala 81:58]
  Mul Mul ( // @[ALU.scala 61:28]
    .clock(Mul_clock),
    .reset(Mul_reset),
    .io_mul_valid(Mul_io_mul_valid),
    .io_mulw(Mul_io_mulw),
    .io_multiplicand(Mul_io_multiplicand),
    .io_multiplier(Mul_io_multiplier),
    .io_out_valid(Mul_io_out_valid),
    .io_out_ready(Mul_io_out_ready),
    .io_result_hi(Mul_io_result_hi),
    .io_result_lo(Mul_io_result_lo)
  );
  Div Div ( // @[ALU.scala 62:28]
    .clock(Div_clock),
    .reset(Div_reset),
    .io_dividend(Div_io_dividend),
    .io_divisor(Div_io_divisor),
    .io_div_valid(Div_io_div_valid),
    .io_divw(Div_io_divw),
    .io_div_signed(Div_io_div_signed),
    .io_out_valid(Div_io_out_valid),
    .io_out_ready(Div_io_out_ready),
    .io_quotient(Div_io_quotient),
    .io_remainder(Div_io_remainder)
  );
  assign io_alu_busy = mul_valid ? ~Mul_io_out_valid : div_valid & ~Div_io_out_valid; // @[ALU.scala 164:23]
  assign io_alu_res = alu_res[63:0]; // @[ALU.scala 165:16]
  assign Mul_clock = clock;
  assign Mul_reset = reset;
  assign Mul_io_mul_valid = mul_valid & io_src_valid; // @[ALU.scala 63:39]
  assign Mul_io_mulw = io_ALUop == 32'h12; // @[ALU.scala 46:22]
  assign Mul_io_multiplicand = io_src1_value; // @[ALU.scala 67:29]
  assign Mul_io_multiplier = io_src2_value; // @[ALU.scala 68:27]
  assign Mul_io_out_ready = io_res_ready; // @[ALU.scala 69:26]
  assign Div_clock = clock;
  assign Div_reset = reset;
  assign Div_io_dividend = io_src1_value; // @[ALU.scala 71:25]
  assign Div_io_divisor = io_src2_value; // @[ALU.scala 72:24]
  assign Div_io_div_valid = div_valid & io_src_valid; // @[ALU.scala 73:39]
  assign Div_io_divw = 32'h32 == io_ALUop | (32'h14 == io_ALUop | (32'h35 == io_ALUop | 32'h13 == io_ALUop)); // @[Mux.scala 81:58]
  assign Div_io_div_signed = 32'h14 == io_ALUop | (32'h34 == io_ALUop | (32'h13 == io_ALUop | 32'h31 == io_ALUop)); // @[Mux.scala 81:58]
  assign Div_io_out_ready = io_res_ready; // @[ALU.scala 77:26]
endmodule
module EXU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_ds_to_es_valid,
  input         io_ms_allowin,
  output        io_es_allowin,
  input  [31:0] io_ALUop,
  input  [63:0] io_src1_value,
  input  [63:0] io_src2_value,
  input  [4:0]  io_rf_dst,
  input  [63:0] io_store_data,
  output        io_es_to_ms_valid,
  input  [2:0]  io_load_type,
  output [63:0] io_to_ms_pc,
  output [63:0] io_to_ms_alures,
  output [63:0] io_to_ms_store_data,
  output        io_to_ms_wen,
  output [7:0]  io_to_ms_wstrb,
  output        io_to_ms_ren,
  output [63:0] io_to_ms_maddr,
  output [4:0]  io_to_ms_rf_dst,
  output        io_to_ms_rf_we,
  output [2:0]  io_to_ms_load_type,
  input         io_ctrl_sign_reg_write,
  input         io_ctrl_sign_Writemem_en,
  input         io_ctrl_sign_Readmem_en,
  input  [7:0]  io_ctrl_sign_Wmask,
  output        io_es_valid,
  output        io_es_rf_we,
  output [4:0]  io_es_rf_dst,
  output        io_es_fwd_ready,
  output [63:0] io_es_fwd_res,
  output        io_es_ld
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  ALU_clock; // @[EXU.scala 40:21]
  wire  ALU_reset; // @[EXU.scala 40:21]
  wire [63:0] ALU_io_src1_value; // @[EXU.scala 40:21]
  wire [63:0] ALU_io_src2_value; // @[EXU.scala 40:21]
  wire [31:0] ALU_io_ALUop; // @[EXU.scala 40:21]
  wire  ALU_io_src_valid; // @[EXU.scala 40:21]
  wire  ALU_io_alu_busy; // @[EXU.scala 40:21]
  wire  ALU_io_res_ready; // @[EXU.scala 40:21]
  wire [63:0] ALU_io_alu_res; // @[EXU.scala 40:21]
  reg [63:0] es_pc; // @[EXU.scala 42:24]
  reg  es_valid; // @[EXU.scala 43:27]
  reg [4:0] es_rd; // @[EXU.scala 47:24]
  reg  es_rf_we; // @[EXU.scala 48:27]
  reg [63:0] src1_value; // @[EXU.scala 50:29]
  reg [63:0] src2_value; // @[EXU.scala 51:29]
  reg [63:0] store_data; // @[EXU.scala 52:29]
  reg [7:0] st_wstrb; // @[EXU.scala 53:27]
  reg  st_we; // @[EXU.scala 54:24]
  reg  ld_we; // @[EXU.scala 55:24]
  reg [31:0] ALUop; // @[EXU.scala 57:24]
  reg [2:0] load_type; // @[EXU.scala 58:28]
  wire  es_ready_go = ~ALU_io_alu_busy; // @[EXU.scala 78:20]
  wire  es_allowin = ~es_valid | es_ready_go & io_ms_allowin; // @[EXU.scala 80:29]
  ALU ALU ( // @[EXU.scala 40:21]
    .clock(ALU_clock),
    .reset(ALU_reset),
    .io_src1_value(ALU_io_src1_value),
    .io_src2_value(ALU_io_src2_value),
    .io_ALUop(ALU_io_ALUop),
    .io_src_valid(ALU_io_src_valid),
    .io_alu_busy(ALU_io_alu_busy),
    .io_res_ready(ALU_io_res_ready),
    .io_alu_res(ALU_io_alu_res)
  );
  assign io_es_allowin = ~es_valid | es_ready_go & io_ms_allowin; // @[EXU.scala 80:29]
  assign io_es_to_ms_valid = es_valid & es_ready_go; // @[EXU.scala 79:32]
  assign io_to_ms_pc = es_pc; // @[EXU.scala 112:17]
  assign io_to_ms_alures = ALU_io_alu_res; // @[EXU.scala 56:23 98:13]
  assign io_to_ms_store_data = store_data; // @[EXU.scala 115:25]
  assign io_to_ms_wen = st_we; // @[EXU.scala 116:18]
  assign io_to_ms_wstrb = st_wstrb; // @[EXU.scala 117:20]
  assign io_to_ms_ren = ld_we; // @[EXU.scala 118:18]
  assign io_to_ms_maddr = ALU_io_alu_res; // @[EXU.scala 56:23 98:13]
  assign io_to_ms_rf_dst = es_rd; // @[EXU.scala 120:21]
  assign io_to_ms_rf_we = es_rf_we; // @[EXU.scala 121:20]
  assign io_to_ms_load_type = load_type; // @[EXU.scala 125:24]
  assign io_es_valid = es_valid; // @[EXU.scala 122:17]
  assign io_es_rf_we = es_rf_we; // @[EXU.scala 124:17]
  assign io_es_rf_dst = es_rd; // @[EXU.scala 123:18]
  assign io_es_fwd_ready = es_valid & es_ready_go; // @[EXU.scala 79:32]
  assign io_es_fwd_res = ALU_io_alu_res; // @[EXU.scala 56:23 98:13]
  assign io_es_ld = ld_we & es_valid; // @[EXU.scala 128:23]
  assign ALU_clock = clock;
  assign ALU_reset = reset;
  assign ALU_io_src1_value = ALUop == 32'h6 ? es_pc : src1_value; // @[EXU.scala 94:26]
  assign ALU_io_src2_value = src2_value; // @[EXU.scala 95:20]
  assign ALU_io_ALUop = ALUop; // @[EXU.scala 96:15]
  assign ALU_io_src_valid = es_valid; // @[EXU.scala 97:19]
  assign ALU_io_res_ready = io_ms_allowin; // @[EXU.scala 99:19]
  always @(posedge clock) begin
    if (reset) begin // @[EXU.scala 42:24]
      es_pc <= 64'h0; // @[EXU.scala 42:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      es_pc <= io_pc; // @[EXU.scala 64:15]
    end
    if (reset) begin // @[EXU.scala 43:27]
      es_valid <= 1'h0; // @[EXU.scala 43:27]
    end else if (es_allowin) begin // @[EXU.scala 60:21]
      es_valid <= io_ds_to_es_valid; // @[EXU.scala 61:18]
    end
    if (reset) begin // @[EXU.scala 47:24]
      es_rd <= 5'h0; // @[EXU.scala 47:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      es_rd <= io_rf_dst; // @[EXU.scala 69:15]
    end
    if (reset) begin // @[EXU.scala 48:27]
      es_rf_we <= 1'h0; // @[EXU.scala 48:27]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      es_rf_we <= io_ctrl_sign_reg_write; // @[EXU.scala 65:18]
    end
    if (reset) begin // @[EXU.scala 50:29]
      src1_value <= 64'h0; // @[EXU.scala 50:29]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      src1_value <= io_src1_value; // @[EXU.scala 67:20]
    end
    if (reset) begin // @[EXU.scala 51:29]
      src2_value <= 64'h0; // @[EXU.scala 51:29]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      src2_value <= io_src2_value; // @[EXU.scala 68:20]
    end
    if (reset) begin // @[EXU.scala 52:29]
      store_data <= 64'h0; // @[EXU.scala 52:29]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      store_data <= io_store_data; // @[EXU.scala 70:20]
    end
    if (reset) begin // @[EXU.scala 53:27]
      st_wstrb <= 8'h0; // @[EXU.scala 53:27]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      st_wstrb <= io_ctrl_sign_Wmask; // @[EXU.scala 71:18]
    end
    if (reset) begin // @[EXU.scala 54:24]
      st_we <= 1'h0; // @[EXU.scala 54:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      st_we <= io_ctrl_sign_Writemem_en; // @[EXU.scala 72:15]
    end
    if (reset) begin // @[EXU.scala 55:24]
      ld_we <= 1'h0; // @[EXU.scala 55:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      ld_we <= io_ctrl_sign_Readmem_en; // @[EXU.scala 73:15]
    end
    if (reset) begin // @[EXU.scala 57:24]
      ALUop <= 32'h0; // @[EXU.scala 57:24]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      ALUop <= io_ALUop; // @[EXU.scala 74:15]
    end
    if (reset) begin // @[EXU.scala 58:28]
      load_type <= 3'h0; // @[EXU.scala 58:28]
    end else if (io_ds_to_es_valid & es_allowin) begin // @[EXU.scala 63:42]
      load_type <= io_load_type; // @[EXU.scala 75:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  es_pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  es_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  es_rd = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  es_rf_we = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  src1_value = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  src2_value = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  store_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  st_wstrb = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  st_we = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ld_we = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ALUop = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  load_type = _RAND_11[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_es_to_ms_valid,
  output        io_ms_allowin,
  input         io_rf_we,
  input  [4:0]  io_rf_dst,
  input  [63:0] io_alu_res,
  input  [63:0] io_store_data,
  input  [2:0]  io_load_type,
  input         io_wen,
  input  [7:0]  io_wstrb,
  input         io_ren,
  input  [63:0] io_maddr,
  output [63:0] io_to_ws_pc,
  output [63:0] io_ms_final_res,
  output        io_ms_to_ws_valid,
  output        io_to_ws_rf_we,
  output [4:0]  io_to_ws_rf_dst,
  output        io_ms_valid,
  output        io_ms_rf_we,
  output [4:0]  io_ms_rf_dst,
  output        io_ms_fwd_ready,
  output [63:0] io_ms_fwd_res,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [63:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg  ms_valid; // @[LSU.scala 36:27]
  reg [63:0] ms_pc; // @[LSU.scala 37:24]
  reg  ms_rf_we; // @[LSU.scala 41:27]
  reg [4:0] ms_rf_dst; // @[LSU.scala 42:28]
  reg [63:0] ms_res; // @[LSU.scala 43:25]
  reg [63:0] store_data; // @[LSU.scala 45:29]
  reg  wen; // @[LSU.scala 46:22]
  reg [7:0] wstrb; // @[LSU.scala 47:24]
  reg  ren; // @[LSU.scala 48:22]
  reg [63:0] maddr; // @[LSU.scala 49:24]
  reg [2:0] load_type; // @[LSU.scala 50:28]
  wire  ms_ready_go = wen & io_axi_in_bvalid | ren & io_axi_in_rvalid | ~(wen | ren); // @[LSU.scala 70:75]
  wire  ms_allowin = ~ms_valid | ms_ready_go; // @[LSU.scala 71:29]
  wire [31:0] _rdata_T_2 = io_axi_in_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rdata_T_4 = {_rdata_T_2,io_axi_in_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdata_T_7 = {56'h0,io_axi_in_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdata_T_10 = {32'h0,io_axi_in_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [47:0] _rdata_T_13 = io_axi_in_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rdata_T_15 = {_rdata_T_13,io_axi_in_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [55:0] _rdata_T_18 = io_axi_in_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rdata_T_20 = {_rdata_T_18,io_axi_in_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdata_T_23 = {48'h0,io_axi_in_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdata_T_25 = 3'h1 == load_type ? _rdata_T_4 : io_axi_in_rdata; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_27 = 3'h2 == load_type ? io_axi_in_rdata : _rdata_T_25; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_29 = 3'h3 == load_type ? _rdata_T_7 : _rdata_T_27; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_31 = 3'h4 == load_type ? _rdata_T_10 : _rdata_T_29; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_33 = 3'h5 == load_type ? _rdata_T_15 : _rdata_T_31; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_35 = 3'h6 == load_type ? _rdata_T_20 : _rdata_T_33; // @[Mux.scala 81:58]
  wire [63:0] rdata = 3'h7 == load_type ? _rdata_T_23 : _rdata_T_35; // @[Mux.scala 81:58]
  wire  _io_ms_final_res_T = load_type != 3'h0; // @[LSU.scala 115:37]
  assign io_ms_allowin = ~ms_valid | ms_ready_go; // @[LSU.scala 71:29]
  assign io_to_ws_pc = ms_pc; // @[LSU.scala 119:17]
  assign io_ms_final_res = load_type != 3'h0 ? rdata : ms_res; // @[LSU.scala 115:27]
  assign io_ms_to_ws_valid = ms_valid & ms_ready_go; // @[LSU.scala 72:32]
  assign io_to_ws_rf_we = ms_rf_we; // @[LSU.scala 118:20]
  assign io_to_ws_rf_dst = ms_rf_dst; // @[LSU.scala 117:21]
  assign io_ms_valid = ms_valid; // @[LSU.scala 121:17]
  assign io_ms_rf_we = ms_rf_we & ms_valid; // @[LSU.scala 123:28]
  assign io_ms_rf_dst = ms_rf_dst; // @[LSU.scala 122:18]
  assign io_ms_fwd_ready = ms_valid & ms_ready_go; // @[LSU.scala 72:32]
  assign io_ms_fwd_res = _io_ms_final_res_T ? rdata : ms_res; // @[LSU.scala 126:25]
  assign io_axi_out_araddr = maddr[31:0]; // @[LSU.scala 88:23]
  assign io_axi_out_arvalid = ren & ms_valid; // @[LSU.scala 89:31]
  assign io_axi_out_awaddr = maddr[31:0]; // @[LSU.scala 94:23]
  assign io_axi_out_awvalid = wen & ms_valid; // @[LSU.scala 95:31]
  assign io_axi_out_wdata = store_data; // @[LSU.scala 99:22]
  assign io_axi_out_wstrb = wstrb; // @[LSU.scala 100:22]
  assign io_axi_out_wvalid = wen; // @[LSU.scala 102:23]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 36:27]
      ms_valid <= 1'h0; // @[LSU.scala 36:27]
    end else if (ms_allowin) begin // @[LSU.scala 53:21]
      ms_valid <= io_es_to_ms_valid; // @[LSU.scala 54:18]
    end
    if (reset) begin // @[LSU.scala 37:24]
      ms_pc <= 64'h0; // @[LSU.scala 37:24]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      ms_pc <= io_pc; // @[LSU.scala 57:15]
    end
    if (reset) begin // @[LSU.scala 41:27]
      ms_rf_we <= 1'h0; // @[LSU.scala 41:27]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      ms_rf_we <= io_rf_we; // @[LSU.scala 58:18]
    end
    if (reset) begin // @[LSU.scala 42:28]
      ms_rf_dst <= 5'h0; // @[LSU.scala 42:28]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      ms_rf_dst <= io_rf_dst; // @[LSU.scala 59:19]
    end
    if (reset) begin // @[LSU.scala 43:25]
      ms_res <= 64'h0; // @[LSU.scala 43:25]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      ms_res <= io_alu_res; // @[LSU.scala 60:16]
    end
    if (reset) begin // @[LSU.scala 45:29]
      store_data <= 64'h0; // @[LSU.scala 45:29]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      store_data <= io_store_data; // @[LSU.scala 61:20]
    end
    if (reset) begin // @[LSU.scala 46:22]
      wen <= 1'h0; // @[LSU.scala 46:22]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      wen <= io_wen; // @[LSU.scala 62:13]
    end
    if (reset) begin // @[LSU.scala 47:24]
      wstrb <= 8'h0; // @[LSU.scala 47:24]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      wstrb <= io_wstrb; // @[LSU.scala 63:15]
    end
    if (reset) begin // @[LSU.scala 48:22]
      ren <= 1'h0; // @[LSU.scala 48:22]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      ren <= io_ren; // @[LSU.scala 64:13]
    end
    if (reset) begin // @[LSU.scala 49:24]
      maddr <= 64'h0; // @[LSU.scala 49:24]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      maddr <= io_maddr; // @[LSU.scala 65:15]
    end
    if (reset) begin // @[LSU.scala 50:28]
      load_type <= 3'h0; // @[LSU.scala 50:28]
    end else if (io_es_to_ms_valid & ms_allowin) begin // @[LSU.scala 56:40]
      load_type <= io_load_type; // @[LSU.scala 66:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ms_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  ms_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  ms_rf_we = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ms_rf_dst = _RAND_3[4:0];
  _RAND_4 = {2{`RANDOM}};
  ms_res = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  store_data = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  wen = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wstrb = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  ren = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  maddr = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  load_type = _RAND_10[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_ms_to_ws_valid,
  input  [63:0] io_ms_final_res,
  input         io_rf_we,
  input  [4:0]  io_rf_dst,
  output        io_we,
  output [4:0]  io_waddr,
  output [63:0] io_wdata,
  output        io_ws_valid,
  output        io_ws_rf_we,
  output [4:0]  io_ws_rf_dst,
  output [63:0] io_ws_fwd_res,
  output [63:0] io_ws_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  ws_valid; // @[WBU.scala 25:27]
  reg [63:0] ws_pc; // @[WBU.scala 26:24]
  reg  ws_rf_we; // @[WBU.scala 30:27]
  reg [4:0] ws_rf_dst; // @[WBU.scala 31:28]
  reg [63:0] ws_res; // @[WBU.scala 32:25]
  assign io_we = ws_rf_we & ws_valid; // @[WBU.scala 61:22]
  assign io_waddr = ws_rf_dst; // @[WBU.scala 62:14]
  assign io_wdata = ws_res; // @[WBU.scala 63:14]
  assign io_ws_valid = ws_valid; // @[WBU.scala 64:17]
  assign io_ws_rf_we = ws_rf_we; // @[WBU.scala 66:17]
  assign io_ws_rf_dst = ws_rf_dst; // @[WBU.scala 65:18]
  assign io_ws_fwd_res = ws_res; // @[WBU.scala 68:19]
  assign io_ws_pc = ws_pc; // @[WBU.scala 69:14]
  always @(posedge clock) begin
    if (reset) begin // @[WBU.scala 25:27]
      ws_valid <= 1'h0; // @[WBU.scala 25:27]
    end else begin
      ws_valid <= io_ms_to_ws_valid;
    end
    if (reset) begin // @[WBU.scala 26:24]
      ws_pc <= 64'h0; // @[WBU.scala 26:24]
    end else if (io_ms_to_ws_valid) begin // @[WBU.scala 43:40]
      ws_pc <= io_pc; // @[WBU.scala 44:15]
    end
    if (reset) begin // @[WBU.scala 30:27]
      ws_rf_we <= 1'h0; // @[WBU.scala 30:27]
    end else if (io_ms_to_ws_valid) begin // @[WBU.scala 43:40]
      ws_rf_we <= io_rf_we; // @[WBU.scala 45:18]
    end
    if (reset) begin // @[WBU.scala 31:28]
      ws_rf_dst <= 5'h0; // @[WBU.scala 31:28]
    end else if (io_ms_to_ws_valid) begin // @[WBU.scala 43:40]
      ws_rf_dst <= io_rf_dst; // @[WBU.scala 46:19]
    end
    if (reset) begin // @[WBU.scala 32:25]
      ws_res <= 64'h0; // @[WBU.scala 32:25]
    end else if (io_ms_to_ws_valid) begin // @[WBU.scala 43:40]
      ws_res <= io_ms_final_res; // @[WBU.scala 47:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ws_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  ws_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  ws_rf_we = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ws_rf_dst = _RAND_3[4:0];
  _RAND_4 = {2{`RANDOM}};
  ws_res = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI_ARBITER(
  input         clock,
  input         reset,
  input  [31:0] io_ifu_axi_in_araddr,
  input  [7:0]  io_ifu_axi_in_arlen,
  input         io_ifu_axi_in_arvalid,
  input         io_ifu_axi_in_rready,
  output [63:0] io_ifu_axi_out_rdata,
  output        io_ifu_axi_out_rlast,
  output        io_ifu_axi_out_rvalid,
  input  [31:0] io_lsu_axi_in_araddr,
  input  [7:0]  io_lsu_axi_in_arlen,
  input         io_lsu_axi_in_arvalid,
  input         io_lsu_axi_in_rready,
  input  [31:0] io_lsu_axi_in_awaddr,
  input  [7:0]  io_lsu_axi_in_awlen,
  input         io_lsu_axi_in_awvalid,
  input  [63:0] io_lsu_axi_in_wdata,
  input  [7:0]  io_lsu_axi_in_wstrb,
  input         io_lsu_axi_in_wvalid,
  input         io_lsu_axi_in_bready,
  output [63:0] io_lsu_axi_out_rdata,
  output        io_lsu_axi_out_rlast,
  output        io_lsu_axi_out_rvalid,
  output        io_lsu_axi_out_wready,
  output        io_lsu_axi_out_bvalid,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rlast,
  input         io_axi_in_rvalid,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output [7:0]  io_axi_out_arlen,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output [7:0]  io_axi_out_awlen,
  output        io_axi_out_awvalid,
  output [63:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[axi_arbiter.scala 18:24]
  wire [1:0] _GEN_0 = io_ifu_axi_in_arvalid ? 2'h1 : state; // @[axi_arbiter.scala 59:46 60:23 18:24]
  wire [31:0] _GEN_1 = io_ifu_axi_in_arvalid ? io_ifu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 59:46 61:28 65:28]
  wire [7:0] _GEN_2 = io_ifu_axi_in_arvalid ? io_ifu_axi_in_arlen : 8'h0; // @[axi_arbiter.scala 59:46 61:28 65:28]
  wire  _GEN_6 = io_ifu_axi_in_arvalid & io_ifu_axi_in_rready; // @[axi_arbiter.scala 59:46 61:28 65:28]
  wire [63:0] _GEN_18 = io_ifu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 59:46 62:32 67:32]
  wire  _GEN_19 = io_ifu_axi_in_arvalid & io_axi_in_rlast; // @[axi_arbiter.scala 59:46 62:32 67:32]
  wire  _GEN_20 = io_ifu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 59:46 62:32 67:32]
  wire [31:0] _GEN_32 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_araddr : _GEN_1; // @[axi_arbiter.scala 54:46 56:28]
  wire [7:0] _GEN_33 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_arlen : _GEN_2; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_36 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_arvalid : io_ifu_axi_in_arvalid; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_37 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_rready : _GEN_6; // @[axi_arbiter.scala 54:46 56:28]
  wire [31:0] _GEN_38 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 54:46 56:28]
  wire [7:0] _GEN_39 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_awlen : 8'h0; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_42 = io_lsu_axi_in_arvalid & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 54:46 56:28]
  wire [63:0] _GEN_43 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wdata : 64'h0; // @[axi_arbiter.scala 54:46 56:28]
  wire [7:0] _GEN_44 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_46 = io_lsu_axi_in_arvalid & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 54:46 56:28]
  wire  _GEN_47 = io_lsu_axi_in_arvalid & io_lsu_axi_in_bready; // @[axi_arbiter.scala 54:46 56:28]
  wire [63:0] _GEN_49 = io_lsu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 54:46 57:32]
  wire  _GEN_50 = io_lsu_axi_in_arvalid & io_axi_in_rlast; // @[axi_arbiter.scala 54:46 57:32]
  wire  _GEN_51 = io_lsu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 54:46 57:32]
  wire  _GEN_53 = io_lsu_axi_in_arvalid & io_axi_in_wready; // @[axi_arbiter.scala 54:46 57:32]
  wire  _GEN_54 = io_lsu_axi_in_arvalid & io_axi_in_bvalid; // @[axi_arbiter.scala 54:46 57:32]
  wire [63:0] _GEN_56 = io_lsu_axi_in_arvalid ? 64'h0 : _GEN_18; // @[axi_arbiter.scala 54:46 58:32]
  wire  _GEN_57 = io_lsu_axi_in_arvalid ? 1'h0 : _GEN_19; // @[axi_arbiter.scala 54:46 58:32]
  wire  _GEN_58 = io_lsu_axi_in_arvalid ? 1'h0 : _GEN_20; // @[axi_arbiter.scala 54:46 58:32]
  wire [31:0] _GEN_63 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_araddr : _GEN_32; // @[axi_arbiter.scala 49:40 51:28]
  wire [7:0] _GEN_64 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_arlen : _GEN_33; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_67 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_arvalid : _GEN_36; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_68 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_rready : _GEN_37; // @[axi_arbiter.scala 49:40 51:28]
  wire [31:0] _GEN_69 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awaddr : _GEN_38; // @[axi_arbiter.scala 49:40 51:28]
  wire [7:0] _GEN_70 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awlen : _GEN_39; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_73 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awvalid : _GEN_42; // @[axi_arbiter.scala 49:40 51:28]
  wire [63:0] _GEN_74 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wdata : _GEN_43; // @[axi_arbiter.scala 49:40 51:28]
  wire [7:0] _GEN_75 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wstrb : _GEN_44; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_77 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wvalid : _GEN_46; // @[axi_arbiter.scala 49:40 51:28]
  wire  _GEN_78 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_bready : _GEN_47; // @[axi_arbiter.scala 49:40 51:28]
  wire [63:0] _GEN_80 = io_lsu_axi_in_awvalid ? io_axi_in_rdata : _GEN_49; // @[axi_arbiter.scala 49:40 52:32]
  wire  _GEN_81 = io_lsu_axi_in_awvalid ? io_axi_in_rlast : _GEN_50; // @[axi_arbiter.scala 49:40 52:32]
  wire  _GEN_82 = io_lsu_axi_in_awvalid ? io_axi_in_rvalid : _GEN_51; // @[axi_arbiter.scala 49:40 52:32]
  wire  _GEN_84 = io_lsu_axi_in_awvalid ? io_axi_in_wready : _GEN_53; // @[axi_arbiter.scala 49:40 52:32]
  wire  _GEN_85 = io_lsu_axi_in_awvalid ? io_axi_in_bvalid : _GEN_54; // @[axi_arbiter.scala 49:40 52:32]
  wire [63:0] _GEN_87 = io_lsu_axi_in_awvalid ? 64'h0 : _GEN_56; // @[axi_arbiter.scala 49:40 53:32]
  wire  _GEN_88 = io_lsu_axi_in_awvalid ? 1'h0 : _GEN_57; // @[axi_arbiter.scala 49:40 53:32]
  wire  _GEN_89 = io_lsu_axi_in_awvalid ? 1'h0 : _GEN_58; // @[axi_arbiter.scala 49:40 53:32]
  wire [1:0] _GEN_94 = io_lsu_axi_out_rvalid & io_lsu_axi_in_rready & io_lsu_axi_out_rlast ? 2'h0 : state; // @[axi_arbiter.scala 82:88 83:23 18:24]
  wire [1:0] _GEN_95 = io_lsu_axi_out_bvalid & io_lsu_axi_in_bready ? 2'h0 : state; // @[axi_arbiter.scala 90:64 91:23 18:24]
  wire [31:0] _GEN_96 = state == 2'h3 ? io_lsu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [7:0] _GEN_97 = state == 2'h3 ? io_lsu_axi_in_arlen : 8'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_100 = state == 2'h3 & io_lsu_axi_in_arvalid; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_101 = state == 2'h3 & io_lsu_axi_in_rready; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [31:0] _GEN_102 = state == 2'h3 ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [7:0] _GEN_103 = state == 2'h3 ? io_lsu_axi_in_awlen : 8'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_106 = state == 2'h3 & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [63:0] _GEN_107 = state == 2'h3 ? io_lsu_axi_in_wdata : 64'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [7:0] _GEN_108 = state == 2'h3 ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_110 = state == 2'h3 & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire  _GEN_111 = state == 2'h3 & io_lsu_axi_in_bready; // @[axi_arbiter.scala 86:39 87:24 95:24]
  wire [63:0] _GEN_113 = state == 2'h3 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire  _GEN_114 = state == 2'h3 & io_axi_in_rlast; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire  _GEN_115 = state == 2'h3 & io_axi_in_rvalid; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire  _GEN_117 = state == 2'h3 & io_axi_in_wready; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire  _GEN_118 = state == 2'h3 & io_axi_in_bvalid; // @[axi_arbiter.scala 86:39 88:28 96:28]
  wire [1:0] _GEN_126 = state == 2'h3 ? _GEN_95 : state; // @[axi_arbiter.scala 18:24 86:39]
  wire [31:0] _GEN_127 = state == 2'h2 ? io_lsu_axi_in_araddr : _GEN_96; // @[axi_arbiter.scala 78:39 79:24]
  wire [7:0] _GEN_128 = state == 2'h2 ? io_lsu_axi_in_arlen : _GEN_97; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_131 = state == 2'h2 ? io_lsu_axi_in_arvalid : _GEN_100; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_132 = state == 2'h2 ? io_lsu_axi_in_rready : _GEN_101; // @[axi_arbiter.scala 78:39 79:24]
  wire [31:0] _GEN_133 = state == 2'h2 ? io_lsu_axi_in_awaddr : _GEN_102; // @[axi_arbiter.scala 78:39 79:24]
  wire [7:0] _GEN_134 = state == 2'h2 ? io_lsu_axi_in_awlen : _GEN_103; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_137 = state == 2'h2 ? io_lsu_axi_in_awvalid : _GEN_106; // @[axi_arbiter.scala 78:39 79:24]
  wire [63:0] _GEN_138 = state == 2'h2 ? io_lsu_axi_in_wdata : _GEN_107; // @[axi_arbiter.scala 78:39 79:24]
  wire [7:0] _GEN_139 = state == 2'h2 ? io_lsu_axi_in_wstrb : _GEN_108; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_141 = state == 2'h2 ? io_lsu_axi_in_wvalid : _GEN_110; // @[axi_arbiter.scala 78:39 79:24]
  wire  _GEN_142 = state == 2'h2 ? io_lsu_axi_in_bready : _GEN_111; // @[axi_arbiter.scala 78:39 79:24]
  wire [63:0] _GEN_144 = state == 2'h2 ? io_axi_in_rdata : _GEN_113; // @[axi_arbiter.scala 78:39 80:28]
  wire  _GEN_145 = state == 2'h2 ? io_axi_in_rlast : _GEN_114; // @[axi_arbiter.scala 78:39 80:28]
  wire  _GEN_146 = state == 2'h2 ? io_axi_in_rvalid : _GEN_115; // @[axi_arbiter.scala 78:39 80:28]
  wire  _GEN_148 = state == 2'h2 ? io_axi_in_wready : _GEN_117; // @[axi_arbiter.scala 78:39 80:28]
  wire  _GEN_149 = state == 2'h2 ? io_axi_in_bvalid : _GEN_118; // @[axi_arbiter.scala 78:39 80:28]
  wire [31:0] _GEN_158 = state == 2'h1 ? io_ifu_axi_in_araddr : _GEN_127; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_159 = state == 2'h1 ? io_ifu_axi_in_arlen : _GEN_128; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_162 = state == 2'h1 ? io_ifu_axi_in_arvalid : _GEN_131; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_163 = state == 2'h1 ? io_ifu_axi_in_rready : _GEN_132; // @[axi_arbiter.scala 70:39 71:24]
  wire [31:0] _GEN_164 = state == 2'h1 ? 32'h0 : _GEN_133; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_165 = state == 2'h1 ? 8'h0 : _GEN_134; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_168 = state == 2'h1 ? 1'h0 : _GEN_137; // @[axi_arbiter.scala 70:39 71:24]
  wire [63:0] _GEN_169 = state == 2'h1 ? 64'h0 : _GEN_138; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_170 = state == 2'h1 ? 8'h0 : _GEN_139; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_172 = state == 2'h1 ? 1'h0 : _GEN_141; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_173 = state == 2'h1 ? 1'h0 : _GEN_142; // @[axi_arbiter.scala 70:39 71:24]
  wire [63:0] _GEN_175 = state == 2'h1 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_176 = state == 2'h1 & io_axi_in_rlast; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_177 = state == 2'h1 & io_axi_in_rvalid; // @[axi_arbiter.scala 70:39 72:28]
  wire [63:0] _GEN_182 = state == 2'h1 ? 64'h0 : _GEN_144; // @[axi_arbiter.scala 70:39 73:28]
  wire  _GEN_183 = state == 2'h1 ? 1'h0 : _GEN_145; // @[axi_arbiter.scala 70:39 73:28]
  wire  _GEN_184 = state == 2'h1 ? 1'h0 : _GEN_146; // @[axi_arbiter.scala 70:39 73:28]
  wire  _GEN_186 = state == 2'h1 ? 1'h0 : _GEN_148; // @[axi_arbiter.scala 70:39 73:28]
  wire  _GEN_187 = state == 2'h1 ? 1'h0 : _GEN_149; // @[axi_arbiter.scala 70:39 73:28]
  assign io_ifu_axi_out_rdata = state == 2'h0 ? _GEN_87 : _GEN_175; // @[axi_arbiter.scala 48:27]
  assign io_ifu_axi_out_rlast = state == 2'h0 ? _GEN_88 : _GEN_176; // @[axi_arbiter.scala 48:27]
  assign io_ifu_axi_out_rvalid = state == 2'h0 ? _GEN_89 : _GEN_177; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_rdata = state == 2'h0 ? _GEN_80 : _GEN_182; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_rlast = state == 2'h0 ? _GEN_81 : _GEN_183; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_rvalid = state == 2'h0 ? _GEN_82 : _GEN_184; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_wready = state == 2'h0 ? _GEN_84 : _GEN_186; // @[axi_arbiter.scala 48:27]
  assign io_lsu_axi_out_bvalid = state == 2'h0 ? _GEN_85 : _GEN_187; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_araddr = state == 2'h0 ? _GEN_63 : _GEN_158; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_arlen = state == 2'h0 ? _GEN_64 : _GEN_159; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_arvalid = state == 2'h0 ? _GEN_67 : _GEN_162; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_rready = state == 2'h0 ? _GEN_68 : _GEN_163; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_awaddr = state == 2'h0 ? _GEN_69 : _GEN_164; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_awlen = state == 2'h0 ? _GEN_70 : _GEN_165; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_awvalid = state == 2'h0 ? _GEN_73 : _GEN_168; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_wdata = state == 2'h0 ? _GEN_74 : _GEN_169; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_wstrb = state == 2'h0 ? _GEN_75 : _GEN_170; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_wvalid = state == 2'h0 ? _GEN_77 : _GEN_172; // @[axi_arbiter.scala 48:27]
  assign io_axi_out_bready = state == 2'h0 ? _GEN_78 : _GEN_173; // @[axi_arbiter.scala 48:27]
  always @(posedge clock) begin
    if (reset) begin // @[axi_arbiter.scala 18:24]
      state <= 2'h0; // @[axi_arbiter.scala 18:24]
    end else if (state == 2'h0) begin // @[axi_arbiter.scala 48:27]
      if (io_lsu_axi_in_awvalid) begin // @[axi_arbiter.scala 49:40]
        state <= 2'h3; // @[axi_arbiter.scala 50:23]
      end else if (io_lsu_axi_in_arvalid) begin // @[axi_arbiter.scala 54:46]
        state <= 2'h2; // @[axi_arbiter.scala 55:23]
      end else begin
        state <= _GEN_0;
      end
    end else if (state == 2'h1) begin // @[axi_arbiter.scala 70:39]
      if (io_ifu_axi_out_rvalid & io_ifu_axi_in_rready & io_ifu_axi_out_rlast) begin // @[axi_arbiter.scala 74:88]
        state <= 2'h0; // @[axi_arbiter.scala 75:23]
      end
    end else if (state == 2'h2) begin // @[axi_arbiter.scala 78:39]
      state <= _GEN_94;
    end else begin
      state <= _GEN_126;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module I_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_ifu_araddr,
  input         io_from_ifu_arvalid,
  input         io_from_ifu_rready,
  output        io_to_ifu_arready,
  output [63:0] io_to_ifu_rdata,
  output        io_to_ifu_rvalid,
  output [31:0] io_to_axi_araddr,
  output [7:0]  io_to_axi_arlen,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rlast,
  input         io_from_axi_rvalid,
  output        io_cache_init,
  input         io_clear_cache
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] ram_0_0; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_1; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_2; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_3; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_4; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_5; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_6; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_7; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_8; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_9; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_10; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_11; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_12; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_13; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_14; // @[i_cache.scala 19:24]
  reg [127:0] ram_0_15; // @[i_cache.scala 19:24]
  reg [127:0] ram_1_0; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_1; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_2; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_3; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_4; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_5; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_6; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_7; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_8; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_9; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_10; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_11; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_12; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_13; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_14; // @[i_cache.scala 20:24]
  reg [127:0] ram_1_15; // @[i_cache.scala 20:24]
  reg [127:0] ram_2_0; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_1; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_2; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_3; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_4; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_5; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_6; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_7; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_8; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_9; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_10; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_11; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_12; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_13; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_14; // @[i_cache.scala 21:24]
  reg [127:0] ram_2_15; // @[i_cache.scala 21:24]
  reg [127:0] ram_3_0; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_1; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_2; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_3; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_4; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_5; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_6; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_7; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_8; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_9; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_10; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_11; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_12; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_13; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_14; // @[i_cache.scala 22:24]
  reg [127:0] ram_3_15; // @[i_cache.scala 22:24]
  reg [31:0] tag_0_0; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_1; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_2; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_3; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_4; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_5; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_6; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_7; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_8; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_9; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_10; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_11; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_12; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_13; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_14; // @[i_cache.scala 23:24]
  reg [31:0] tag_0_15; // @[i_cache.scala 23:24]
  reg [31:0] tag_1_0; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_1; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_2; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_3; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_4; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_5; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_6; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_7; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_8; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_9; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_10; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_11; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_12; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_13; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_14; // @[i_cache.scala 24:24]
  reg [31:0] tag_1_15; // @[i_cache.scala 24:24]
  reg [31:0] tag_2_0; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_1; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_2; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_3; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_4; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_5; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_6; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_7; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_8; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_9; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_10; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_11; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_12; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_13; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_14; // @[i_cache.scala 25:24]
  reg [31:0] tag_2_15; // @[i_cache.scala 25:24]
  reg [31:0] tag_3_0; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_1; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_2; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_3; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_4; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_5; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_6; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_7; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_8; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_9; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_10; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_11; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_12; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_13; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_14; // @[i_cache.scala 26:24]
  reg [31:0] tag_3_15; // @[i_cache.scala 26:24]
  reg  valid_0_0; // @[i_cache.scala 27:26]
  reg  valid_0_1; // @[i_cache.scala 27:26]
  reg  valid_0_2; // @[i_cache.scala 27:26]
  reg  valid_0_3; // @[i_cache.scala 27:26]
  reg  valid_0_4; // @[i_cache.scala 27:26]
  reg  valid_0_5; // @[i_cache.scala 27:26]
  reg  valid_0_6; // @[i_cache.scala 27:26]
  reg  valid_0_7; // @[i_cache.scala 27:26]
  reg  valid_0_8; // @[i_cache.scala 27:26]
  reg  valid_0_9; // @[i_cache.scala 27:26]
  reg  valid_0_10; // @[i_cache.scala 27:26]
  reg  valid_0_11; // @[i_cache.scala 27:26]
  reg  valid_0_12; // @[i_cache.scala 27:26]
  reg  valid_0_13; // @[i_cache.scala 27:26]
  reg  valid_0_14; // @[i_cache.scala 27:26]
  reg  valid_0_15; // @[i_cache.scala 27:26]
  reg  valid_1_0; // @[i_cache.scala 28:26]
  reg  valid_1_1; // @[i_cache.scala 28:26]
  reg  valid_1_2; // @[i_cache.scala 28:26]
  reg  valid_1_3; // @[i_cache.scala 28:26]
  reg  valid_1_4; // @[i_cache.scala 28:26]
  reg  valid_1_5; // @[i_cache.scala 28:26]
  reg  valid_1_6; // @[i_cache.scala 28:26]
  reg  valid_1_7; // @[i_cache.scala 28:26]
  reg  valid_1_8; // @[i_cache.scala 28:26]
  reg  valid_1_9; // @[i_cache.scala 28:26]
  reg  valid_1_10; // @[i_cache.scala 28:26]
  reg  valid_1_11; // @[i_cache.scala 28:26]
  reg  valid_1_12; // @[i_cache.scala 28:26]
  reg  valid_1_13; // @[i_cache.scala 28:26]
  reg  valid_1_14; // @[i_cache.scala 28:26]
  reg  valid_1_15; // @[i_cache.scala 28:26]
  reg  valid_2_0; // @[i_cache.scala 29:26]
  reg  valid_2_1; // @[i_cache.scala 29:26]
  reg  valid_2_2; // @[i_cache.scala 29:26]
  reg  valid_2_3; // @[i_cache.scala 29:26]
  reg  valid_2_4; // @[i_cache.scala 29:26]
  reg  valid_2_5; // @[i_cache.scala 29:26]
  reg  valid_2_6; // @[i_cache.scala 29:26]
  reg  valid_2_7; // @[i_cache.scala 29:26]
  reg  valid_2_8; // @[i_cache.scala 29:26]
  reg  valid_2_9; // @[i_cache.scala 29:26]
  reg  valid_2_10; // @[i_cache.scala 29:26]
  reg  valid_2_11; // @[i_cache.scala 29:26]
  reg  valid_2_12; // @[i_cache.scala 29:26]
  reg  valid_2_13; // @[i_cache.scala 29:26]
  reg  valid_2_14; // @[i_cache.scala 29:26]
  reg  valid_2_15; // @[i_cache.scala 29:26]
  reg  valid_3_0; // @[i_cache.scala 30:26]
  reg  valid_3_1; // @[i_cache.scala 30:26]
  reg  valid_3_2; // @[i_cache.scala 30:26]
  reg  valid_3_3; // @[i_cache.scala 30:26]
  reg  valid_3_4; // @[i_cache.scala 30:26]
  reg  valid_3_5; // @[i_cache.scala 30:26]
  reg  valid_3_6; // @[i_cache.scala 30:26]
  reg  valid_3_7; // @[i_cache.scala 30:26]
  reg  valid_3_8; // @[i_cache.scala 30:26]
  reg  valid_3_9; // @[i_cache.scala 30:26]
  reg  valid_3_10; // @[i_cache.scala 30:26]
  reg  valid_3_11; // @[i_cache.scala 30:26]
  reg  valid_3_12; // @[i_cache.scala 30:26]
  reg  valid_3_13; // @[i_cache.scala 30:26]
  reg  valid_3_14; // @[i_cache.scala 30:26]
  reg  valid_3_15; // @[i_cache.scala 30:26]
  reg [31:0] addr; // @[i_cache.scala 32:23]
  reg [63:0] receive_data_0; // @[i_cache.scala 40:31]
  reg [63:0] receive_data_1; // @[i_cache.scala 40:31]
  reg [2:0] receive_num; // @[i_cache.scala 41:30]
  reg [7:0] quene_0; // @[i_cache.scala 42:24]
  reg [7:0] quene_1; // @[i_cache.scala 42:24]
  reg [7:0] quene_2; // @[i_cache.scala 42:24]
  reg [7:0] quene_3; // @[i_cache.scala 42:24]
  reg [7:0] quene_4; // @[i_cache.scala 42:24]
  reg [7:0] quene_5; // @[i_cache.scala 42:24]
  reg [7:0] quene_6; // @[i_cache.scala 42:24]
  reg [7:0] quene_7; // @[i_cache.scala 42:24]
  reg [7:0] quene_8; // @[i_cache.scala 42:24]
  reg [7:0] quene_9; // @[i_cache.scala 42:24]
  reg [7:0] quene_10; // @[i_cache.scala 42:24]
  reg [7:0] quene_11; // @[i_cache.scala 42:24]
  reg [7:0] quene_12; // @[i_cache.scala 42:24]
  reg [7:0] quene_13; // @[i_cache.scala 42:24]
  reg [7:0] quene_14; // @[i_cache.scala 42:24]
  reg [7:0] quene_15; // @[i_cache.scala 42:24]
  wire [3:0] offset = addr[3:0]; // @[i_cache.scala 44:22]
  wire [3:0] index = addr[7:4]; // @[i_cache.scala 45:21]
  wire [23:0] tag = addr[31:8]; // @[i_cache.scala 46:19]
  wire [6:0] shift_bit = {offset, 3'h0}; // @[i_cache.scala 47:28]
  wire [31:0] _GEN_1 = 4'h1 == index ? tag_0_1 : tag_0_0; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_2 = 4'h2 == index ? tag_0_2 : _GEN_1; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_3 = 4'h3 == index ? tag_0_3 : _GEN_2; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_4 = 4'h4 == index ? tag_0_4 : _GEN_3; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_5 = 4'h5 == index ? tag_0_5 : _GEN_4; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_6 = 4'h6 == index ? tag_0_6 : _GEN_5; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_7 = 4'h7 == index ? tag_0_7 : _GEN_6; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_8 = 4'h8 == index ? tag_0_8 : _GEN_7; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_9 = 4'h9 == index ? tag_0_9 : _GEN_8; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_10 = 4'ha == index ? tag_0_10 : _GEN_9; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_11 = 4'hb == index ? tag_0_11 : _GEN_10; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_12 = 4'hc == index ? tag_0_12 : _GEN_11; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_13 = 4'hd == index ? tag_0_13 : _GEN_12; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_14 = 4'he == index ? tag_0_14 : _GEN_13; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_15 = 4'hf == index ? tag_0_15 : _GEN_14; // @[i_cache.scala 49:{31,31}]
  wire [31:0] _GEN_2929 = {{8'd0}, tag}; // @[i_cache.scala 49:31]
  wire  _GEN_17 = 4'h1 == index ? valid_0_1 : valid_0_0; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_18 = 4'h2 == index ? valid_0_2 : _GEN_17; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_19 = 4'h3 == index ? valid_0_3 : _GEN_18; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_20 = 4'h4 == index ? valid_0_4 : _GEN_19; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_21 = 4'h5 == index ? valid_0_5 : _GEN_20; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_22 = 4'h6 == index ? valid_0_6 : _GEN_21; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_23 = 4'h7 == index ? valid_0_7 : _GEN_22; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_24 = 4'h8 == index ? valid_0_8 : _GEN_23; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_25 = 4'h9 == index ? valid_0_9 : _GEN_24; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_26 = 4'ha == index ? valid_0_10 : _GEN_25; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_27 = 4'hb == index ? valid_0_11 : _GEN_26; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_28 = 4'hc == index ? valid_0_12 : _GEN_27; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_29 = 4'hd == index ? valid_0_13 : _GEN_28; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_30 = 4'he == index ? valid_0_14 : _GEN_29; // @[i_cache.scala 49:{57,57}]
  wire  _GEN_31 = 4'hf == index ? valid_0_15 : _GEN_30; // @[i_cache.scala 49:{57,57}]
  wire  way0_hit = _GEN_15 == _GEN_2929 & _GEN_31; // @[i_cache.scala 49:40]
  wire [31:0] _GEN_33 = 4'h1 == index ? tag_1_1 : tag_1_0; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_34 = 4'h2 == index ? tag_1_2 : _GEN_33; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_35 = 4'h3 == index ? tag_1_3 : _GEN_34; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_36 = 4'h4 == index ? tag_1_4 : _GEN_35; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_37 = 4'h5 == index ? tag_1_5 : _GEN_36; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_38 = 4'h6 == index ? tag_1_6 : _GEN_37; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_39 = 4'h7 == index ? tag_1_7 : _GEN_38; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_40 = 4'h8 == index ? tag_1_8 : _GEN_39; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_41 = 4'h9 == index ? tag_1_9 : _GEN_40; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_42 = 4'ha == index ? tag_1_10 : _GEN_41; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_43 = 4'hb == index ? tag_1_11 : _GEN_42; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_44 = 4'hc == index ? tag_1_12 : _GEN_43; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_45 = 4'hd == index ? tag_1_13 : _GEN_44; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_46 = 4'he == index ? tag_1_14 : _GEN_45; // @[i_cache.scala 51:{31,31}]
  wire [31:0] _GEN_47 = 4'hf == index ? tag_1_15 : _GEN_46; // @[i_cache.scala 51:{31,31}]
  wire  _GEN_49 = 4'h1 == index ? valid_1_1 : valid_1_0; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_50 = 4'h2 == index ? valid_1_2 : _GEN_49; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_51 = 4'h3 == index ? valid_1_3 : _GEN_50; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_52 = 4'h4 == index ? valid_1_4 : _GEN_51; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_53 = 4'h5 == index ? valid_1_5 : _GEN_52; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_54 = 4'h6 == index ? valid_1_6 : _GEN_53; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_55 = 4'h7 == index ? valid_1_7 : _GEN_54; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_56 = 4'h8 == index ? valid_1_8 : _GEN_55; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_57 = 4'h9 == index ? valid_1_9 : _GEN_56; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_58 = 4'ha == index ? valid_1_10 : _GEN_57; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_59 = 4'hb == index ? valid_1_11 : _GEN_58; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_60 = 4'hc == index ? valid_1_12 : _GEN_59; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_61 = 4'hd == index ? valid_1_13 : _GEN_60; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_62 = 4'he == index ? valid_1_14 : _GEN_61; // @[i_cache.scala 51:{57,57}]
  wire  _GEN_63 = 4'hf == index ? valid_1_15 : _GEN_62; // @[i_cache.scala 51:{57,57}]
  wire  way1_hit = _GEN_47 == _GEN_2929 & _GEN_63; // @[i_cache.scala 51:40]
  wire [31:0] _GEN_65 = 4'h1 == index ? tag_2_1 : tag_2_0; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_66 = 4'h2 == index ? tag_2_2 : _GEN_65; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_67 = 4'h3 == index ? tag_2_3 : _GEN_66; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_68 = 4'h4 == index ? tag_2_4 : _GEN_67; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_69 = 4'h5 == index ? tag_2_5 : _GEN_68; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_70 = 4'h6 == index ? tag_2_6 : _GEN_69; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_71 = 4'h7 == index ? tag_2_7 : _GEN_70; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_72 = 4'h8 == index ? tag_2_8 : _GEN_71; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_73 = 4'h9 == index ? tag_2_9 : _GEN_72; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_74 = 4'ha == index ? tag_2_10 : _GEN_73; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_75 = 4'hb == index ? tag_2_11 : _GEN_74; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_76 = 4'hc == index ? tag_2_12 : _GEN_75; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_77 = 4'hd == index ? tag_2_13 : _GEN_76; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_78 = 4'he == index ? tag_2_14 : _GEN_77; // @[i_cache.scala 52:{31,31}]
  wire [31:0] _GEN_79 = 4'hf == index ? tag_2_15 : _GEN_78; // @[i_cache.scala 52:{31,31}]
  wire  _GEN_81 = 4'h1 == index ? valid_2_1 : valid_2_0; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_82 = 4'h2 == index ? valid_2_2 : _GEN_81; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_83 = 4'h3 == index ? valid_2_3 : _GEN_82; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_84 = 4'h4 == index ? valid_2_4 : _GEN_83; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_85 = 4'h5 == index ? valid_2_5 : _GEN_84; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_86 = 4'h6 == index ? valid_2_6 : _GEN_85; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_87 = 4'h7 == index ? valid_2_7 : _GEN_86; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_88 = 4'h8 == index ? valid_2_8 : _GEN_87; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_89 = 4'h9 == index ? valid_2_9 : _GEN_88; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_90 = 4'ha == index ? valid_2_10 : _GEN_89; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_91 = 4'hb == index ? valid_2_11 : _GEN_90; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_92 = 4'hc == index ? valid_2_12 : _GEN_91; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_93 = 4'hd == index ? valid_2_13 : _GEN_92; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_94 = 4'he == index ? valid_2_14 : _GEN_93; // @[i_cache.scala 52:{57,57}]
  wire  _GEN_95 = 4'hf == index ? valid_2_15 : _GEN_94; // @[i_cache.scala 52:{57,57}]
  wire  way2_hit = _GEN_79 == _GEN_2929 & _GEN_95; // @[i_cache.scala 52:40]
  wire [31:0] _GEN_97 = 4'h1 == index ? tag_3_1 : tag_3_0; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_98 = 4'h2 == index ? tag_3_2 : _GEN_97; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_99 = 4'h3 == index ? tag_3_3 : _GEN_98; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_100 = 4'h4 == index ? tag_3_4 : _GEN_99; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_101 = 4'h5 == index ? tag_3_5 : _GEN_100; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_102 = 4'h6 == index ? tag_3_6 : _GEN_101; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_103 = 4'h7 == index ? tag_3_7 : _GEN_102; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_104 = 4'h8 == index ? tag_3_8 : _GEN_103; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_105 = 4'h9 == index ? tag_3_9 : _GEN_104; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_106 = 4'ha == index ? tag_3_10 : _GEN_105; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_107 = 4'hb == index ? tag_3_11 : _GEN_106; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_108 = 4'hc == index ? tag_3_12 : _GEN_107; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_109 = 4'hd == index ? tag_3_13 : _GEN_108; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_110 = 4'he == index ? tag_3_14 : _GEN_109; // @[i_cache.scala 53:{31,31}]
  wire [31:0] _GEN_111 = 4'hf == index ? tag_3_15 : _GEN_110; // @[i_cache.scala 53:{31,31}]
  wire  _GEN_113 = 4'h1 == index ? valid_3_1 : valid_3_0; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_114 = 4'h2 == index ? valid_3_2 : _GEN_113; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_115 = 4'h3 == index ? valid_3_3 : _GEN_114; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_116 = 4'h4 == index ? valid_3_4 : _GEN_115; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_117 = 4'h5 == index ? valid_3_5 : _GEN_116; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_118 = 4'h6 == index ? valid_3_6 : _GEN_117; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_119 = 4'h7 == index ? valid_3_7 : _GEN_118; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_120 = 4'h8 == index ? valid_3_8 : _GEN_119; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_121 = 4'h9 == index ? valid_3_9 : _GEN_120; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_122 = 4'ha == index ? valid_3_10 : _GEN_121; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_123 = 4'hb == index ? valid_3_11 : _GEN_122; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_124 = 4'hc == index ? valid_3_12 : _GEN_123; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_125 = 4'hd == index ? valid_3_13 : _GEN_124; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_126 = 4'he == index ? valid_3_14 : _GEN_125; // @[i_cache.scala 53:{57,57}]
  wire  _GEN_127 = 4'hf == index ? valid_3_15 : _GEN_126; // @[i_cache.scala 53:{57,57}]
  wire  way3_hit = _GEN_111 == _GEN_2929 & _GEN_127; // @[i_cache.scala 53:40]
  wire [2:0] _unuse_way_T_4 = ~_GEN_127 ? 3'h4 : 3'h0; // @[i_cache.scala 54:108]
  wire [2:0] _unuse_way_T_5 = ~_GEN_95 ? 3'h3 : _unuse_way_T_4; // @[i_cache.scala 54:79]
  wire [2:0] _unuse_way_T_6 = ~_GEN_63 ? 3'h2 : _unuse_way_T_5; // @[i_cache.scala 54:50]
  wire [2:0] unuse_way = ~_GEN_31 ? 3'h1 : _unuse_way_T_6; // @[i_cache.scala 54:21]
  reg [2:0] state; // @[i_cache.scala 56:24]
  wire  _T_4 = way0_hit | way1_hit | way2_hit | way3_hit; // @[i_cache.scala 69:46]
  wire [2:0] _GEN_132 = io_from_ifu_rready ? 3'h0 : state; // @[i_cache.scala 56:24 70:41 71:27]
  wire [63:0] _GEN_135 = ~receive_num[0] ? io_from_axi_rdata : receive_data_0; // @[i_cache.scala 40:31 80:{43,43}]
  wire [63:0] _GEN_136 = receive_num[0] ? io_from_axi_rdata : receive_data_1; // @[i_cache.scala 40:31 80:{43,43}]
  wire [2:0] _receive_num_T_1 = receive_num + 3'h1; // @[i_cache.scala 81:44]
  wire [2:0] _GEN_137 = io_from_axi_rlast ? 3'h3 : state; // @[i_cache.scala 56:24 82:40 83:27]
  wire [63:0] _GEN_138 = io_from_axi_rvalid ? _GEN_135 : receive_data_0; // @[i_cache.scala 40:31 79:37]
  wire [63:0] _GEN_139 = io_from_axi_rvalid ? _GEN_136 : receive_data_1; // @[i_cache.scala 40:31 79:37]
  wire [2:0] _GEN_140 = io_from_axi_rvalid ? _receive_num_T_1 : receive_num; // @[i_cache.scala 79:37 81:29 41:30]
  wire [2:0] _GEN_141 = io_from_axi_rvalid ? _GEN_137 : state; // @[i_cache.scala 56:24 79:37]
  wire [127:0] _ram_0_T = {receive_data_1,receive_data_0}; // @[Cat.scala 31:58]
  wire [127:0] _GEN_142 = 4'h0 == index ? _ram_0_T : ram_0_0; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_143 = 4'h1 == index ? _ram_0_T : ram_0_1; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_144 = 4'h2 == index ? _ram_0_T : ram_0_2; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_145 = 4'h3 == index ? _ram_0_T : ram_0_3; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_146 = 4'h4 == index ? _ram_0_T : ram_0_4; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_147 = 4'h5 == index ? _ram_0_T : ram_0_5; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_148 = 4'h6 == index ? _ram_0_T : ram_0_6; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_149 = 4'h7 == index ? _ram_0_T : ram_0_7; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_150 = 4'h8 == index ? _ram_0_T : ram_0_8; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_151 = 4'h9 == index ? _ram_0_T : ram_0_9; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_152 = 4'ha == index ? _ram_0_T : ram_0_10; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_153 = 4'hb == index ? _ram_0_T : ram_0_11; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_154 = 4'hc == index ? _ram_0_T : ram_0_12; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_155 = 4'hd == index ? _ram_0_T : ram_0_13; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_156 = 4'he == index ? _ram_0_T : ram_0_14; // @[i_cache.scala 19:24 90:{30,30}]
  wire [127:0] _GEN_157 = 4'hf == index ? _ram_0_T : ram_0_15; // @[i_cache.scala 19:24 90:{30,30}]
  wire [31:0] _GEN_158 = 4'h0 == index ? _GEN_2929 : tag_0_0; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_159 = 4'h1 == index ? _GEN_2929 : tag_0_1; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_160 = 4'h2 == index ? _GEN_2929 : tag_0_2; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_161 = 4'h3 == index ? _GEN_2929 : tag_0_3; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_162 = 4'h4 == index ? _GEN_2929 : tag_0_4; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_163 = 4'h5 == index ? _GEN_2929 : tag_0_5; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_164 = 4'h6 == index ? _GEN_2929 : tag_0_6; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_165 = 4'h7 == index ? _GEN_2929 : tag_0_7; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_166 = 4'h8 == index ? _GEN_2929 : tag_0_8; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_167 = 4'h9 == index ? _GEN_2929 : tag_0_9; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_168 = 4'ha == index ? _GEN_2929 : tag_0_10; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_169 = 4'hb == index ? _GEN_2929 : tag_0_11; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_170 = 4'hc == index ? _GEN_2929 : tag_0_12; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_171 = 4'hd == index ? _GEN_2929 : tag_0_13; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_172 = 4'he == index ? _GEN_2929 : tag_0_14; // @[i_cache.scala 23:24 91:{30,30}]
  wire [31:0] _GEN_173 = 4'hf == index ? _GEN_2929 : tag_0_15; // @[i_cache.scala 23:24 91:{30,30}]
  wire  _GEN_2941 = 4'h0 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_174 = 4'h0 == index | valid_0_0; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2942 = 4'h1 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_175 = 4'h1 == index | valid_0_1; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2943 = 4'h2 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_176 = 4'h2 == index | valid_0_2; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2944 = 4'h3 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_177 = 4'h3 == index | valid_0_3; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2945 = 4'h4 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_178 = 4'h4 == index | valid_0_4; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2946 = 4'h5 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_179 = 4'h5 == index | valid_0_5; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2947 = 4'h6 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_180 = 4'h6 == index | valid_0_6; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2948 = 4'h7 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_181 = 4'h7 == index | valid_0_7; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2949 = 4'h8 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_182 = 4'h8 == index | valid_0_8; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2950 = 4'h9 == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_183 = 4'h9 == index | valid_0_9; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2951 = 4'ha == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_184 = 4'ha == index | valid_0_10; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2952 = 4'hb == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_185 = 4'hb == index | valid_0_11; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2953 = 4'hc == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_186 = 4'hc == index | valid_0_12; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2954 = 4'hd == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_187 = 4'hd == index | valid_0_13; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2955 = 4'he == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_188 = 4'he == index | valid_0_14; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_2956 = 4'hf == index; // @[i_cache.scala 27:26 92:{32,32}]
  wire  _GEN_189 = 4'hf == index | valid_0_15; // @[i_cache.scala 27:26 92:{32,32}]
  wire [7:0] _GEN_191 = 4'h1 == index ? quene_1 : quene_0; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_192 = 4'h2 == index ? quene_2 : _GEN_191; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_193 = 4'h3 == index ? quene_3 : _GEN_192; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_194 = 4'h4 == index ? quene_4 : _GEN_193; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_195 = 4'h5 == index ? quene_5 : _GEN_194; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_196 = 4'h6 == index ? quene_6 : _GEN_195; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_197 = 4'h7 == index ? quene_7 : _GEN_196; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_198 = 4'h8 == index ? quene_8 : _GEN_197; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_199 = 4'h9 == index ? quene_9 : _GEN_198; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_200 = 4'ha == index ? quene_10 : _GEN_199; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_201 = 4'hb == index ? quene_11 : _GEN_200; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_202 = 4'hc == index ? quene_12 : _GEN_201; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_203 = 4'hd == index ? quene_13 : _GEN_202; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_204 = 4'he == index ? quene_14 : _GEN_203; // @[i_cache.scala 93:{46,46}]
  wire [7:0] _GEN_205 = 4'hf == index ? quene_15 : _GEN_204; // @[i_cache.scala 93:{46,46}]
  wire [9:0] _GEN_2957 = {_GEN_205, 2'h0}; // @[i_cache.scala 93:46]
  wire [10:0] _quene_T = {{1'd0}, _GEN_2957}; // @[i_cache.scala 93:46]
  wire [7:0] _GEN_206 = 4'h0 == index ? _quene_T[7:0] : quene_0; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_207 = 4'h1 == index ? _quene_T[7:0] : quene_1; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_208 = 4'h2 == index ? _quene_T[7:0] : quene_2; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_209 = 4'h3 == index ? _quene_T[7:0] : quene_3; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_210 = 4'h4 == index ? _quene_T[7:0] : quene_4; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_211 = 4'h5 == index ? _quene_T[7:0] : quene_5; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_212 = 4'h6 == index ? _quene_T[7:0] : quene_6; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_213 = 4'h7 == index ? _quene_T[7:0] : quene_7; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_214 = 4'h8 == index ? _quene_T[7:0] : quene_8; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_215 = 4'h9 == index ? _quene_T[7:0] : quene_9; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_216 = 4'ha == index ? _quene_T[7:0] : quene_10; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_217 = 4'hb == index ? _quene_T[7:0] : quene_11; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_218 = 4'hc == index ? _quene_T[7:0] : quene_12; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_219 = 4'hd == index ? _quene_T[7:0] : quene_13; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_220 = 4'he == index ? _quene_T[7:0] : quene_14; // @[i_cache.scala 42:24 93:{30,30}]
  wire [7:0] _GEN_221 = 4'hf == index ? _quene_T[7:0] : quene_15; // @[i_cache.scala 42:24 93:{30,30}]
  wire [127:0] _GEN_222 = 4'h0 == index ? _ram_0_T : ram_1_0; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_223 = 4'h1 == index ? _ram_0_T : ram_1_1; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_224 = 4'h2 == index ? _ram_0_T : ram_1_2; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_225 = 4'h3 == index ? _ram_0_T : ram_1_3; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_226 = 4'h4 == index ? _ram_0_T : ram_1_4; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_227 = 4'h5 == index ? _ram_0_T : ram_1_5; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_228 = 4'h6 == index ? _ram_0_T : ram_1_6; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_229 = 4'h7 == index ? _ram_0_T : ram_1_7; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_230 = 4'h8 == index ? _ram_0_T : ram_1_8; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_231 = 4'h9 == index ? _ram_0_T : ram_1_9; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_232 = 4'ha == index ? _ram_0_T : ram_1_10; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_233 = 4'hb == index ? _ram_0_T : ram_1_11; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_234 = 4'hc == index ? _ram_0_T : ram_1_12; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_235 = 4'hd == index ? _ram_0_T : ram_1_13; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_236 = 4'he == index ? _ram_0_T : ram_1_14; // @[i_cache.scala 20:24 95:{30,30}]
  wire [127:0] _GEN_237 = 4'hf == index ? _ram_0_T : ram_1_15; // @[i_cache.scala 20:24 95:{30,30}]
  wire [31:0] _GEN_238 = 4'h0 == index ? _GEN_2929 : tag_1_0; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_239 = 4'h1 == index ? _GEN_2929 : tag_1_1; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_240 = 4'h2 == index ? _GEN_2929 : tag_1_2; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_241 = 4'h3 == index ? _GEN_2929 : tag_1_3; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_242 = 4'h4 == index ? _GEN_2929 : tag_1_4; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_243 = 4'h5 == index ? _GEN_2929 : tag_1_5; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_244 = 4'h6 == index ? _GEN_2929 : tag_1_6; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_245 = 4'h7 == index ? _GEN_2929 : tag_1_7; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_246 = 4'h8 == index ? _GEN_2929 : tag_1_8; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_247 = 4'h9 == index ? _GEN_2929 : tag_1_9; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_248 = 4'ha == index ? _GEN_2929 : tag_1_10; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_249 = 4'hb == index ? _GEN_2929 : tag_1_11; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_250 = 4'hc == index ? _GEN_2929 : tag_1_12; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_251 = 4'hd == index ? _GEN_2929 : tag_1_13; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_252 = 4'he == index ? _GEN_2929 : tag_1_14; // @[i_cache.scala 24:24 96:{30,30}]
  wire [31:0] _GEN_253 = 4'hf == index ? _GEN_2929 : tag_1_15; // @[i_cache.scala 24:24 96:{30,30}]
  wire  _GEN_254 = _GEN_2941 | valid_1_0; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_255 = _GEN_2942 | valid_1_1; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_256 = _GEN_2943 | valid_1_2; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_257 = _GEN_2944 | valid_1_3; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_258 = _GEN_2945 | valid_1_4; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_259 = _GEN_2946 | valid_1_5; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_260 = _GEN_2947 | valid_1_6; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_261 = _GEN_2948 | valid_1_7; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_262 = _GEN_2949 | valid_1_8; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_263 = _GEN_2950 | valid_1_9; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_264 = _GEN_2951 | valid_1_10; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_265 = _GEN_2952 | valid_1_11; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_266 = _GEN_2953 | valid_1_12; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_267 = _GEN_2954 | valid_1_13; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_268 = _GEN_2955 | valid_1_14; // @[i_cache.scala 28:26 97:{32,32}]
  wire  _GEN_269 = _GEN_2956 | valid_1_15; // @[i_cache.scala 28:26 97:{32,32}]
  wire [10:0] _quene_T_2 = _quene_T | 11'h1; // @[i_cache.scala 98:55]
  wire [7:0] _GEN_270 = 4'h0 == index ? _quene_T_2[7:0] : quene_0; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_271 = 4'h1 == index ? _quene_T_2[7:0] : quene_1; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_272 = 4'h2 == index ? _quene_T_2[7:0] : quene_2; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_273 = 4'h3 == index ? _quene_T_2[7:0] : quene_3; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_274 = 4'h4 == index ? _quene_T_2[7:0] : quene_4; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_275 = 4'h5 == index ? _quene_T_2[7:0] : quene_5; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_276 = 4'h6 == index ? _quene_T_2[7:0] : quene_6; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_277 = 4'h7 == index ? _quene_T_2[7:0] : quene_7; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_278 = 4'h8 == index ? _quene_T_2[7:0] : quene_8; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_279 = 4'h9 == index ? _quene_T_2[7:0] : quene_9; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_280 = 4'ha == index ? _quene_T_2[7:0] : quene_10; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_281 = 4'hb == index ? _quene_T_2[7:0] : quene_11; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_282 = 4'hc == index ? _quene_T_2[7:0] : quene_12; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_283 = 4'hd == index ? _quene_T_2[7:0] : quene_13; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_284 = 4'he == index ? _quene_T_2[7:0] : quene_14; // @[i_cache.scala 42:24 98:{30,30}]
  wire [7:0] _GEN_285 = 4'hf == index ? _quene_T_2[7:0] : quene_15; // @[i_cache.scala 42:24 98:{30,30}]
  wire [127:0] _GEN_286 = 4'h0 == index ? _ram_0_T : ram_2_0; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_287 = 4'h1 == index ? _ram_0_T : ram_2_1; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_288 = 4'h2 == index ? _ram_0_T : ram_2_2; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_289 = 4'h3 == index ? _ram_0_T : ram_2_3; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_290 = 4'h4 == index ? _ram_0_T : ram_2_4; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_291 = 4'h5 == index ? _ram_0_T : ram_2_5; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_292 = 4'h6 == index ? _ram_0_T : ram_2_6; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_293 = 4'h7 == index ? _ram_0_T : ram_2_7; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_294 = 4'h8 == index ? _ram_0_T : ram_2_8; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_295 = 4'h9 == index ? _ram_0_T : ram_2_9; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_296 = 4'ha == index ? _ram_0_T : ram_2_10; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_297 = 4'hb == index ? _ram_0_T : ram_2_11; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_298 = 4'hc == index ? _ram_0_T : ram_2_12; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_299 = 4'hd == index ? _ram_0_T : ram_2_13; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_300 = 4'he == index ? _ram_0_T : ram_2_14; // @[i_cache.scala 100:{30,30} 21:24]
  wire [127:0] _GEN_301 = 4'hf == index ? _ram_0_T : ram_2_15; // @[i_cache.scala 100:{30,30} 21:24]
  wire [31:0] _GEN_302 = 4'h0 == index ? _GEN_2929 : tag_2_0; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_303 = 4'h1 == index ? _GEN_2929 : tag_2_1; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_304 = 4'h2 == index ? _GEN_2929 : tag_2_2; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_305 = 4'h3 == index ? _GEN_2929 : tag_2_3; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_306 = 4'h4 == index ? _GEN_2929 : tag_2_4; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_307 = 4'h5 == index ? _GEN_2929 : tag_2_5; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_308 = 4'h6 == index ? _GEN_2929 : tag_2_6; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_309 = 4'h7 == index ? _GEN_2929 : tag_2_7; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_310 = 4'h8 == index ? _GEN_2929 : tag_2_8; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_311 = 4'h9 == index ? _GEN_2929 : tag_2_9; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_312 = 4'ha == index ? _GEN_2929 : tag_2_10; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_313 = 4'hb == index ? _GEN_2929 : tag_2_11; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_314 = 4'hc == index ? _GEN_2929 : tag_2_12; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_315 = 4'hd == index ? _GEN_2929 : tag_2_13; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_316 = 4'he == index ? _GEN_2929 : tag_2_14; // @[i_cache.scala 101:{30,30} 25:24]
  wire [31:0] _GEN_317 = 4'hf == index ? _GEN_2929 : tag_2_15; // @[i_cache.scala 101:{30,30} 25:24]
  wire  _GEN_318 = _GEN_2941 | valid_2_0; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_319 = _GEN_2942 | valid_2_1; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_320 = _GEN_2943 | valid_2_2; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_321 = _GEN_2944 | valid_2_3; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_322 = _GEN_2945 | valid_2_4; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_323 = _GEN_2946 | valid_2_5; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_324 = _GEN_2947 | valid_2_6; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_325 = _GEN_2948 | valid_2_7; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_326 = _GEN_2949 | valid_2_8; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_327 = _GEN_2950 | valid_2_9; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_328 = _GEN_2951 | valid_2_10; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_329 = _GEN_2952 | valid_2_11; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_330 = _GEN_2953 | valid_2_12; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_331 = _GEN_2954 | valid_2_13; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_332 = _GEN_2955 | valid_2_14; // @[i_cache.scala 102:{32,32} 29:26]
  wire  _GEN_333 = _GEN_2956 | valid_2_15; // @[i_cache.scala 102:{32,32} 29:26]
  wire [10:0] _quene_T_4 = _quene_T | 11'h2; // @[i_cache.scala 103:55]
  wire [7:0] _GEN_334 = 4'h0 == index ? _quene_T_4[7:0] : quene_0; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_335 = 4'h1 == index ? _quene_T_4[7:0] : quene_1; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_336 = 4'h2 == index ? _quene_T_4[7:0] : quene_2; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_337 = 4'h3 == index ? _quene_T_4[7:0] : quene_3; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_338 = 4'h4 == index ? _quene_T_4[7:0] : quene_4; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_339 = 4'h5 == index ? _quene_T_4[7:0] : quene_5; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_340 = 4'h6 == index ? _quene_T_4[7:0] : quene_6; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_341 = 4'h7 == index ? _quene_T_4[7:0] : quene_7; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_342 = 4'h8 == index ? _quene_T_4[7:0] : quene_8; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_343 = 4'h9 == index ? _quene_T_4[7:0] : quene_9; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_344 = 4'ha == index ? _quene_T_4[7:0] : quene_10; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_345 = 4'hb == index ? _quene_T_4[7:0] : quene_11; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_346 = 4'hc == index ? _quene_T_4[7:0] : quene_12; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_347 = 4'hd == index ? _quene_T_4[7:0] : quene_13; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_348 = 4'he == index ? _quene_T_4[7:0] : quene_14; // @[i_cache.scala 103:{30,30} 42:24]
  wire [7:0] _GEN_349 = 4'hf == index ? _quene_T_4[7:0] : quene_15; // @[i_cache.scala 103:{30,30} 42:24]
  wire [127:0] _GEN_350 = 4'h0 == index ? _ram_0_T : ram_3_0; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_351 = 4'h1 == index ? _ram_0_T : ram_3_1; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_352 = 4'h2 == index ? _ram_0_T : ram_3_2; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_353 = 4'h3 == index ? _ram_0_T : ram_3_3; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_354 = 4'h4 == index ? _ram_0_T : ram_3_4; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_355 = 4'h5 == index ? _ram_0_T : ram_3_5; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_356 = 4'h6 == index ? _ram_0_T : ram_3_6; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_357 = 4'h7 == index ? _ram_0_T : ram_3_7; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_358 = 4'h8 == index ? _ram_0_T : ram_3_8; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_359 = 4'h9 == index ? _ram_0_T : ram_3_9; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_360 = 4'ha == index ? _ram_0_T : ram_3_10; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_361 = 4'hb == index ? _ram_0_T : ram_3_11; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_362 = 4'hc == index ? _ram_0_T : ram_3_12; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_363 = 4'hd == index ? _ram_0_T : ram_3_13; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_364 = 4'he == index ? _ram_0_T : ram_3_14; // @[i_cache.scala 105:{30,30} 22:24]
  wire [127:0] _GEN_365 = 4'hf == index ? _ram_0_T : ram_3_15; // @[i_cache.scala 105:{30,30} 22:24]
  wire [31:0] _GEN_366 = 4'h0 == index ? _GEN_2929 : tag_3_0; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_367 = 4'h1 == index ? _GEN_2929 : tag_3_1; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_368 = 4'h2 == index ? _GEN_2929 : tag_3_2; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_369 = 4'h3 == index ? _GEN_2929 : tag_3_3; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_370 = 4'h4 == index ? _GEN_2929 : tag_3_4; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_371 = 4'h5 == index ? _GEN_2929 : tag_3_5; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_372 = 4'h6 == index ? _GEN_2929 : tag_3_6; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_373 = 4'h7 == index ? _GEN_2929 : tag_3_7; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_374 = 4'h8 == index ? _GEN_2929 : tag_3_8; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_375 = 4'h9 == index ? _GEN_2929 : tag_3_9; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_376 = 4'ha == index ? _GEN_2929 : tag_3_10; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_377 = 4'hb == index ? _GEN_2929 : tag_3_11; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_378 = 4'hc == index ? _GEN_2929 : tag_3_12; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_379 = 4'hd == index ? _GEN_2929 : tag_3_13; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_380 = 4'he == index ? _GEN_2929 : tag_3_14; // @[i_cache.scala 106:{30,30} 26:24]
  wire [31:0] _GEN_381 = 4'hf == index ? _GEN_2929 : tag_3_15; // @[i_cache.scala 106:{30,30} 26:24]
  wire  _GEN_382 = _GEN_2941 | valid_3_0; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_383 = _GEN_2942 | valid_3_1; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_384 = _GEN_2943 | valid_3_2; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_385 = _GEN_2944 | valid_3_3; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_386 = _GEN_2945 | valid_3_4; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_387 = _GEN_2946 | valid_3_5; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_388 = _GEN_2947 | valid_3_6; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_389 = _GEN_2948 | valid_3_7; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_390 = _GEN_2949 | valid_3_8; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_391 = _GEN_2950 | valid_3_9; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_392 = _GEN_2951 | valid_3_10; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_393 = _GEN_2952 | valid_3_11; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_394 = _GEN_2953 | valid_3_12; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_395 = _GEN_2954 | valid_3_13; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_396 = _GEN_2955 | valid_3_14; // @[i_cache.scala 107:{32,32} 30:26]
  wire  _GEN_397 = _GEN_2956 | valid_3_15; // @[i_cache.scala 107:{32,32} 30:26]
  wire [10:0] _quene_T_6 = _quene_T | 11'h3; // @[i_cache.scala 108:55]
  wire [7:0] _GEN_398 = 4'h0 == index ? _quene_T_6[7:0] : quene_0; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_399 = 4'h1 == index ? _quene_T_6[7:0] : quene_1; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_400 = 4'h2 == index ? _quene_T_6[7:0] : quene_2; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_401 = 4'h3 == index ? _quene_T_6[7:0] : quene_3; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_402 = 4'h4 == index ? _quene_T_6[7:0] : quene_4; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_403 = 4'h5 == index ? _quene_T_6[7:0] : quene_5; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_404 = 4'h6 == index ? _quene_T_6[7:0] : quene_6; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_405 = 4'h7 == index ? _quene_T_6[7:0] : quene_7; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_406 = 4'h8 == index ? _quene_T_6[7:0] : quene_8; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_407 = 4'h9 == index ? _quene_T_6[7:0] : quene_9; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_408 = 4'ha == index ? _quene_T_6[7:0] : quene_10; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_409 = 4'hb == index ? _quene_T_6[7:0] : quene_11; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_410 = 4'hc == index ? _quene_T_6[7:0] : quene_12; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_411 = 4'hd == index ? _quene_T_6[7:0] : quene_13; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_412 = 4'he == index ? _quene_T_6[7:0] : quene_14; // @[i_cache.scala 108:{30,30} 42:24]
  wire [7:0] _GEN_413 = 4'hf == index ? _quene_T_6[7:0] : quene_15; // @[i_cache.scala 108:{30,30} 42:24]
  wire [127:0] _GEN_670 = _GEN_205[7:6] == 2'h2 ? _GEN_286 : ram_2_0; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_671 = _GEN_205[7:6] == 2'h2 ? _GEN_287 : ram_2_1; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_672 = _GEN_205[7:6] == 2'h2 ? _GEN_288 : ram_2_2; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_673 = _GEN_205[7:6] == 2'h2 ? _GEN_289 : ram_2_3; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_674 = _GEN_205[7:6] == 2'h2 ? _GEN_290 : ram_2_4; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_675 = _GEN_205[7:6] == 2'h2 ? _GEN_291 : ram_2_5; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_676 = _GEN_205[7:6] == 2'h2 ? _GEN_292 : ram_2_6; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_677 = _GEN_205[7:6] == 2'h2 ? _GEN_293 : ram_2_7; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_678 = _GEN_205[7:6] == 2'h2 ? _GEN_294 : ram_2_8; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_679 = _GEN_205[7:6] == 2'h2 ? _GEN_295 : ram_2_9; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_680 = _GEN_205[7:6] == 2'h2 ? _GEN_296 : ram_2_10; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_681 = _GEN_205[7:6] == 2'h2 ? _GEN_297 : ram_2_11; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_682 = _GEN_205[7:6] == 2'h2 ? _GEN_298 : ram_2_12; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_683 = _GEN_205[7:6] == 2'h2 ? _GEN_299 : ram_2_13; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_684 = _GEN_205[7:6] == 2'h2 ? _GEN_300 : ram_2_14; // @[i_cache.scala 120:52 21:24]
  wire [127:0] _GEN_685 = _GEN_205[7:6] == 2'h2 ? _GEN_301 : ram_2_15; // @[i_cache.scala 120:52 21:24]
  wire [31:0] _GEN_686 = _GEN_205[7:6] == 2'h2 ? _GEN_302 : tag_2_0; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_687 = _GEN_205[7:6] == 2'h2 ? _GEN_303 : tag_2_1; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_688 = _GEN_205[7:6] == 2'h2 ? _GEN_304 : tag_2_2; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_689 = _GEN_205[7:6] == 2'h2 ? _GEN_305 : tag_2_3; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_690 = _GEN_205[7:6] == 2'h2 ? _GEN_306 : tag_2_4; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_691 = _GEN_205[7:6] == 2'h2 ? _GEN_307 : tag_2_5; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_692 = _GEN_205[7:6] == 2'h2 ? _GEN_308 : tag_2_6; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_693 = _GEN_205[7:6] == 2'h2 ? _GEN_309 : tag_2_7; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_694 = _GEN_205[7:6] == 2'h2 ? _GEN_310 : tag_2_8; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_695 = _GEN_205[7:6] == 2'h2 ? _GEN_311 : tag_2_9; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_696 = _GEN_205[7:6] == 2'h2 ? _GEN_312 : tag_2_10; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_697 = _GEN_205[7:6] == 2'h2 ? _GEN_313 : tag_2_11; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_698 = _GEN_205[7:6] == 2'h2 ? _GEN_314 : tag_2_12; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_699 = _GEN_205[7:6] == 2'h2 ? _GEN_315 : tag_2_13; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_700 = _GEN_205[7:6] == 2'h2 ? _GEN_316 : tag_2_14; // @[i_cache.scala 120:52 25:24]
  wire [31:0] _GEN_701 = _GEN_205[7:6] == 2'h2 ? _GEN_317 : tag_2_15; // @[i_cache.scala 120:52 25:24]
  wire  _GEN_702 = _GEN_205[7:6] == 2'h2 ? _GEN_318 : valid_2_0; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_703 = _GEN_205[7:6] == 2'h2 ? _GEN_319 : valid_2_1; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_704 = _GEN_205[7:6] == 2'h2 ? _GEN_320 : valid_2_2; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_705 = _GEN_205[7:6] == 2'h2 ? _GEN_321 : valid_2_3; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_706 = _GEN_205[7:6] == 2'h2 ? _GEN_322 : valid_2_4; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_707 = _GEN_205[7:6] == 2'h2 ? _GEN_323 : valid_2_5; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_708 = _GEN_205[7:6] == 2'h2 ? _GEN_324 : valid_2_6; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_709 = _GEN_205[7:6] == 2'h2 ? _GEN_325 : valid_2_7; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_710 = _GEN_205[7:6] == 2'h2 ? _GEN_326 : valid_2_8; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_711 = _GEN_205[7:6] == 2'h2 ? _GEN_327 : valid_2_9; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_712 = _GEN_205[7:6] == 2'h2 ? _GEN_328 : valid_2_10; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_713 = _GEN_205[7:6] == 2'h2 ? _GEN_329 : valid_2_11; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_714 = _GEN_205[7:6] == 2'h2 ? _GEN_330 : valid_2_12; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_715 = _GEN_205[7:6] == 2'h2 ? _GEN_331 : valid_2_13; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_716 = _GEN_205[7:6] == 2'h2 ? _GEN_332 : valid_2_14; // @[i_cache.scala 120:52 29:26]
  wire  _GEN_717 = _GEN_205[7:6] == 2'h2 ? _GEN_333 : valid_2_15; // @[i_cache.scala 120:52 29:26]
  wire [7:0] _GEN_718 = _GEN_205[7:6] == 2'h2 ? _GEN_334 : _GEN_398; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_719 = _GEN_205[7:6] == 2'h2 ? _GEN_335 : _GEN_399; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_720 = _GEN_205[7:6] == 2'h2 ? _GEN_336 : _GEN_400; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_721 = _GEN_205[7:6] == 2'h2 ? _GEN_337 : _GEN_401; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_722 = _GEN_205[7:6] == 2'h2 ? _GEN_338 : _GEN_402; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_723 = _GEN_205[7:6] == 2'h2 ? _GEN_339 : _GEN_403; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_724 = _GEN_205[7:6] == 2'h2 ? _GEN_340 : _GEN_404; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_725 = _GEN_205[7:6] == 2'h2 ? _GEN_341 : _GEN_405; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_726 = _GEN_205[7:6] == 2'h2 ? _GEN_342 : _GEN_406; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_727 = _GEN_205[7:6] == 2'h2 ? _GEN_343 : _GEN_407; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_728 = _GEN_205[7:6] == 2'h2 ? _GEN_344 : _GEN_408; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_729 = _GEN_205[7:6] == 2'h2 ? _GEN_345 : _GEN_409; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_730 = _GEN_205[7:6] == 2'h2 ? _GEN_346 : _GEN_410; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_731 = _GEN_205[7:6] == 2'h2 ? _GEN_347 : _GEN_411; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_732 = _GEN_205[7:6] == 2'h2 ? _GEN_348 : _GEN_412; // @[i_cache.scala 120:52]
  wire [7:0] _GEN_733 = _GEN_205[7:6] == 2'h2 ? _GEN_349 : _GEN_413; // @[i_cache.scala 120:52]
  wire [127:0] _GEN_734 = _GEN_205[7:6] == 2'h2 ? ram_3_0 : _GEN_350; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_735 = _GEN_205[7:6] == 2'h2 ? ram_3_1 : _GEN_351; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_736 = _GEN_205[7:6] == 2'h2 ? ram_3_2 : _GEN_352; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_737 = _GEN_205[7:6] == 2'h2 ? ram_3_3 : _GEN_353; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_738 = _GEN_205[7:6] == 2'h2 ? ram_3_4 : _GEN_354; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_739 = _GEN_205[7:6] == 2'h2 ? ram_3_5 : _GEN_355; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_740 = _GEN_205[7:6] == 2'h2 ? ram_3_6 : _GEN_356; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_741 = _GEN_205[7:6] == 2'h2 ? ram_3_7 : _GEN_357; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_742 = _GEN_205[7:6] == 2'h2 ? ram_3_8 : _GEN_358; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_743 = _GEN_205[7:6] == 2'h2 ? ram_3_9 : _GEN_359; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_744 = _GEN_205[7:6] == 2'h2 ? ram_3_10 : _GEN_360; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_745 = _GEN_205[7:6] == 2'h2 ? ram_3_11 : _GEN_361; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_746 = _GEN_205[7:6] == 2'h2 ? ram_3_12 : _GEN_362; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_747 = _GEN_205[7:6] == 2'h2 ? ram_3_13 : _GEN_363; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_748 = _GEN_205[7:6] == 2'h2 ? ram_3_14 : _GEN_364; // @[i_cache.scala 120:52 22:24]
  wire [127:0] _GEN_749 = _GEN_205[7:6] == 2'h2 ? ram_3_15 : _GEN_365; // @[i_cache.scala 120:52 22:24]
  wire [31:0] _GEN_750 = _GEN_205[7:6] == 2'h2 ? tag_3_0 : _GEN_366; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_751 = _GEN_205[7:6] == 2'h2 ? tag_3_1 : _GEN_367; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_752 = _GEN_205[7:6] == 2'h2 ? tag_3_2 : _GEN_368; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_753 = _GEN_205[7:6] == 2'h2 ? tag_3_3 : _GEN_369; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_754 = _GEN_205[7:6] == 2'h2 ? tag_3_4 : _GEN_370; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_755 = _GEN_205[7:6] == 2'h2 ? tag_3_5 : _GEN_371; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_756 = _GEN_205[7:6] == 2'h2 ? tag_3_6 : _GEN_372; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_757 = _GEN_205[7:6] == 2'h2 ? tag_3_7 : _GEN_373; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_758 = _GEN_205[7:6] == 2'h2 ? tag_3_8 : _GEN_374; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_759 = _GEN_205[7:6] == 2'h2 ? tag_3_9 : _GEN_375; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_760 = _GEN_205[7:6] == 2'h2 ? tag_3_10 : _GEN_376; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_761 = _GEN_205[7:6] == 2'h2 ? tag_3_11 : _GEN_377; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_762 = _GEN_205[7:6] == 2'h2 ? tag_3_12 : _GEN_378; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_763 = _GEN_205[7:6] == 2'h2 ? tag_3_13 : _GEN_379; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_764 = _GEN_205[7:6] == 2'h2 ? tag_3_14 : _GEN_380; // @[i_cache.scala 120:52 26:24]
  wire [31:0] _GEN_765 = _GEN_205[7:6] == 2'h2 ? tag_3_15 : _GEN_381; // @[i_cache.scala 120:52 26:24]
  wire  _GEN_766 = _GEN_205[7:6] == 2'h2 ? valid_3_0 : _GEN_382; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_767 = _GEN_205[7:6] == 2'h2 ? valid_3_1 : _GEN_383; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_768 = _GEN_205[7:6] == 2'h2 ? valid_3_2 : _GEN_384; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_769 = _GEN_205[7:6] == 2'h2 ? valid_3_3 : _GEN_385; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_770 = _GEN_205[7:6] == 2'h2 ? valid_3_4 : _GEN_386; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_771 = _GEN_205[7:6] == 2'h2 ? valid_3_5 : _GEN_387; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_772 = _GEN_205[7:6] == 2'h2 ? valid_3_6 : _GEN_388; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_773 = _GEN_205[7:6] == 2'h2 ? valid_3_7 : _GEN_389; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_774 = _GEN_205[7:6] == 2'h2 ? valid_3_8 : _GEN_390; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_775 = _GEN_205[7:6] == 2'h2 ? valid_3_9 : _GEN_391; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_776 = _GEN_205[7:6] == 2'h2 ? valid_3_10 : _GEN_392; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_777 = _GEN_205[7:6] == 2'h2 ? valid_3_11 : _GEN_393; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_778 = _GEN_205[7:6] == 2'h2 ? valid_3_12 : _GEN_394; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_779 = _GEN_205[7:6] == 2'h2 ? valid_3_13 : _GEN_395; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_780 = _GEN_205[7:6] == 2'h2 ? valid_3_14 : _GEN_396; // @[i_cache.scala 120:52 30:26]
  wire  _GEN_781 = _GEN_205[7:6] == 2'h2 ? valid_3_15 : _GEN_397; // @[i_cache.scala 120:52 30:26]
  wire [127:0] _GEN_782 = _GEN_205[7:6] == 2'h1 ? _GEN_222 : ram_1_0; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_783 = _GEN_205[7:6] == 2'h1 ? _GEN_223 : ram_1_1; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_784 = _GEN_205[7:6] == 2'h1 ? _GEN_224 : ram_1_2; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_785 = _GEN_205[7:6] == 2'h1 ? _GEN_225 : ram_1_3; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_786 = _GEN_205[7:6] == 2'h1 ? _GEN_226 : ram_1_4; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_787 = _GEN_205[7:6] == 2'h1 ? _GEN_227 : ram_1_5; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_788 = _GEN_205[7:6] == 2'h1 ? _GEN_228 : ram_1_6; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_789 = _GEN_205[7:6] == 2'h1 ? _GEN_229 : ram_1_7; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_790 = _GEN_205[7:6] == 2'h1 ? _GEN_230 : ram_1_8; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_791 = _GEN_205[7:6] == 2'h1 ? _GEN_231 : ram_1_9; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_792 = _GEN_205[7:6] == 2'h1 ? _GEN_232 : ram_1_10; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_793 = _GEN_205[7:6] == 2'h1 ? _GEN_233 : ram_1_11; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_794 = _GEN_205[7:6] == 2'h1 ? _GEN_234 : ram_1_12; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_795 = _GEN_205[7:6] == 2'h1 ? _GEN_235 : ram_1_13; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_796 = _GEN_205[7:6] == 2'h1 ? _GEN_236 : ram_1_14; // @[i_cache.scala 115:52 20:24]
  wire [127:0] _GEN_797 = _GEN_205[7:6] == 2'h1 ? _GEN_237 : ram_1_15; // @[i_cache.scala 115:52 20:24]
  wire [31:0] _GEN_798 = _GEN_205[7:6] == 2'h1 ? _GEN_238 : tag_1_0; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_799 = _GEN_205[7:6] == 2'h1 ? _GEN_239 : tag_1_1; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_800 = _GEN_205[7:6] == 2'h1 ? _GEN_240 : tag_1_2; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_801 = _GEN_205[7:6] == 2'h1 ? _GEN_241 : tag_1_3; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_802 = _GEN_205[7:6] == 2'h1 ? _GEN_242 : tag_1_4; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_803 = _GEN_205[7:6] == 2'h1 ? _GEN_243 : tag_1_5; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_804 = _GEN_205[7:6] == 2'h1 ? _GEN_244 : tag_1_6; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_805 = _GEN_205[7:6] == 2'h1 ? _GEN_245 : tag_1_7; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_806 = _GEN_205[7:6] == 2'h1 ? _GEN_246 : tag_1_8; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_807 = _GEN_205[7:6] == 2'h1 ? _GEN_247 : tag_1_9; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_808 = _GEN_205[7:6] == 2'h1 ? _GEN_248 : tag_1_10; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_809 = _GEN_205[7:6] == 2'h1 ? _GEN_249 : tag_1_11; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_810 = _GEN_205[7:6] == 2'h1 ? _GEN_250 : tag_1_12; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_811 = _GEN_205[7:6] == 2'h1 ? _GEN_251 : tag_1_13; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_812 = _GEN_205[7:6] == 2'h1 ? _GEN_252 : tag_1_14; // @[i_cache.scala 115:52 24:24]
  wire [31:0] _GEN_813 = _GEN_205[7:6] == 2'h1 ? _GEN_253 : tag_1_15; // @[i_cache.scala 115:52 24:24]
  wire  _GEN_814 = _GEN_205[7:6] == 2'h1 ? _GEN_254 : valid_1_0; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_815 = _GEN_205[7:6] == 2'h1 ? _GEN_255 : valid_1_1; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_816 = _GEN_205[7:6] == 2'h1 ? _GEN_256 : valid_1_2; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_817 = _GEN_205[7:6] == 2'h1 ? _GEN_257 : valid_1_3; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_818 = _GEN_205[7:6] == 2'h1 ? _GEN_258 : valid_1_4; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_819 = _GEN_205[7:6] == 2'h1 ? _GEN_259 : valid_1_5; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_820 = _GEN_205[7:6] == 2'h1 ? _GEN_260 : valid_1_6; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_821 = _GEN_205[7:6] == 2'h1 ? _GEN_261 : valid_1_7; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_822 = _GEN_205[7:6] == 2'h1 ? _GEN_262 : valid_1_8; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_823 = _GEN_205[7:6] == 2'h1 ? _GEN_263 : valid_1_9; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_824 = _GEN_205[7:6] == 2'h1 ? _GEN_264 : valid_1_10; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_825 = _GEN_205[7:6] == 2'h1 ? _GEN_265 : valid_1_11; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_826 = _GEN_205[7:6] == 2'h1 ? _GEN_266 : valid_1_12; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_827 = _GEN_205[7:6] == 2'h1 ? _GEN_267 : valid_1_13; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_828 = _GEN_205[7:6] == 2'h1 ? _GEN_268 : valid_1_14; // @[i_cache.scala 115:52 28:26]
  wire  _GEN_829 = _GEN_205[7:6] == 2'h1 ? _GEN_269 : valid_1_15; // @[i_cache.scala 115:52 28:26]
  wire [7:0] _GEN_830 = _GEN_205[7:6] == 2'h1 ? _GEN_270 : _GEN_718; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_831 = _GEN_205[7:6] == 2'h1 ? _GEN_271 : _GEN_719; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_832 = _GEN_205[7:6] == 2'h1 ? _GEN_272 : _GEN_720; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_833 = _GEN_205[7:6] == 2'h1 ? _GEN_273 : _GEN_721; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_834 = _GEN_205[7:6] == 2'h1 ? _GEN_274 : _GEN_722; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_835 = _GEN_205[7:6] == 2'h1 ? _GEN_275 : _GEN_723; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_836 = _GEN_205[7:6] == 2'h1 ? _GEN_276 : _GEN_724; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_837 = _GEN_205[7:6] == 2'h1 ? _GEN_277 : _GEN_725; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_838 = _GEN_205[7:6] == 2'h1 ? _GEN_278 : _GEN_726; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_839 = _GEN_205[7:6] == 2'h1 ? _GEN_279 : _GEN_727; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_840 = _GEN_205[7:6] == 2'h1 ? _GEN_280 : _GEN_728; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_841 = _GEN_205[7:6] == 2'h1 ? _GEN_281 : _GEN_729; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_842 = _GEN_205[7:6] == 2'h1 ? _GEN_282 : _GEN_730; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_843 = _GEN_205[7:6] == 2'h1 ? _GEN_283 : _GEN_731; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_844 = _GEN_205[7:6] == 2'h1 ? _GEN_284 : _GEN_732; // @[i_cache.scala 115:52]
  wire [7:0] _GEN_845 = _GEN_205[7:6] == 2'h1 ? _GEN_285 : _GEN_733; // @[i_cache.scala 115:52]
  wire [127:0] _GEN_846 = _GEN_205[7:6] == 2'h1 ? ram_2_0 : _GEN_670; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_847 = _GEN_205[7:6] == 2'h1 ? ram_2_1 : _GEN_671; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_848 = _GEN_205[7:6] == 2'h1 ? ram_2_2 : _GEN_672; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_849 = _GEN_205[7:6] == 2'h1 ? ram_2_3 : _GEN_673; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_850 = _GEN_205[7:6] == 2'h1 ? ram_2_4 : _GEN_674; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_851 = _GEN_205[7:6] == 2'h1 ? ram_2_5 : _GEN_675; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_852 = _GEN_205[7:6] == 2'h1 ? ram_2_6 : _GEN_676; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_853 = _GEN_205[7:6] == 2'h1 ? ram_2_7 : _GEN_677; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_854 = _GEN_205[7:6] == 2'h1 ? ram_2_8 : _GEN_678; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_855 = _GEN_205[7:6] == 2'h1 ? ram_2_9 : _GEN_679; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_856 = _GEN_205[7:6] == 2'h1 ? ram_2_10 : _GEN_680; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_857 = _GEN_205[7:6] == 2'h1 ? ram_2_11 : _GEN_681; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_858 = _GEN_205[7:6] == 2'h1 ? ram_2_12 : _GEN_682; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_859 = _GEN_205[7:6] == 2'h1 ? ram_2_13 : _GEN_683; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_860 = _GEN_205[7:6] == 2'h1 ? ram_2_14 : _GEN_684; // @[i_cache.scala 115:52 21:24]
  wire [127:0] _GEN_861 = _GEN_205[7:6] == 2'h1 ? ram_2_15 : _GEN_685; // @[i_cache.scala 115:52 21:24]
  wire [31:0] _GEN_862 = _GEN_205[7:6] == 2'h1 ? tag_2_0 : _GEN_686; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_863 = _GEN_205[7:6] == 2'h1 ? tag_2_1 : _GEN_687; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_864 = _GEN_205[7:6] == 2'h1 ? tag_2_2 : _GEN_688; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_865 = _GEN_205[7:6] == 2'h1 ? tag_2_3 : _GEN_689; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_866 = _GEN_205[7:6] == 2'h1 ? tag_2_4 : _GEN_690; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_867 = _GEN_205[7:6] == 2'h1 ? tag_2_5 : _GEN_691; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_868 = _GEN_205[7:6] == 2'h1 ? tag_2_6 : _GEN_692; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_869 = _GEN_205[7:6] == 2'h1 ? tag_2_7 : _GEN_693; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_870 = _GEN_205[7:6] == 2'h1 ? tag_2_8 : _GEN_694; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_871 = _GEN_205[7:6] == 2'h1 ? tag_2_9 : _GEN_695; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_872 = _GEN_205[7:6] == 2'h1 ? tag_2_10 : _GEN_696; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_873 = _GEN_205[7:6] == 2'h1 ? tag_2_11 : _GEN_697; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_874 = _GEN_205[7:6] == 2'h1 ? tag_2_12 : _GEN_698; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_875 = _GEN_205[7:6] == 2'h1 ? tag_2_13 : _GEN_699; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_876 = _GEN_205[7:6] == 2'h1 ? tag_2_14 : _GEN_700; // @[i_cache.scala 115:52 25:24]
  wire [31:0] _GEN_877 = _GEN_205[7:6] == 2'h1 ? tag_2_15 : _GEN_701; // @[i_cache.scala 115:52 25:24]
  wire  _GEN_878 = _GEN_205[7:6] == 2'h1 ? valid_2_0 : _GEN_702; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_879 = _GEN_205[7:6] == 2'h1 ? valid_2_1 : _GEN_703; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_880 = _GEN_205[7:6] == 2'h1 ? valid_2_2 : _GEN_704; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_881 = _GEN_205[7:6] == 2'h1 ? valid_2_3 : _GEN_705; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_882 = _GEN_205[7:6] == 2'h1 ? valid_2_4 : _GEN_706; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_883 = _GEN_205[7:6] == 2'h1 ? valid_2_5 : _GEN_707; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_884 = _GEN_205[7:6] == 2'h1 ? valid_2_6 : _GEN_708; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_885 = _GEN_205[7:6] == 2'h1 ? valid_2_7 : _GEN_709; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_886 = _GEN_205[7:6] == 2'h1 ? valid_2_8 : _GEN_710; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_887 = _GEN_205[7:6] == 2'h1 ? valid_2_9 : _GEN_711; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_888 = _GEN_205[7:6] == 2'h1 ? valid_2_10 : _GEN_712; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_889 = _GEN_205[7:6] == 2'h1 ? valid_2_11 : _GEN_713; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_890 = _GEN_205[7:6] == 2'h1 ? valid_2_12 : _GEN_714; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_891 = _GEN_205[7:6] == 2'h1 ? valid_2_13 : _GEN_715; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_892 = _GEN_205[7:6] == 2'h1 ? valid_2_14 : _GEN_716; // @[i_cache.scala 115:52 29:26]
  wire  _GEN_893 = _GEN_205[7:6] == 2'h1 ? valid_2_15 : _GEN_717; // @[i_cache.scala 115:52 29:26]
  wire [127:0] _GEN_894 = _GEN_205[7:6] == 2'h1 ? ram_3_0 : _GEN_734; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_895 = _GEN_205[7:6] == 2'h1 ? ram_3_1 : _GEN_735; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_896 = _GEN_205[7:6] == 2'h1 ? ram_3_2 : _GEN_736; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_897 = _GEN_205[7:6] == 2'h1 ? ram_3_3 : _GEN_737; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_898 = _GEN_205[7:6] == 2'h1 ? ram_3_4 : _GEN_738; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_899 = _GEN_205[7:6] == 2'h1 ? ram_3_5 : _GEN_739; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_900 = _GEN_205[7:6] == 2'h1 ? ram_3_6 : _GEN_740; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_901 = _GEN_205[7:6] == 2'h1 ? ram_3_7 : _GEN_741; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_902 = _GEN_205[7:6] == 2'h1 ? ram_3_8 : _GEN_742; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_903 = _GEN_205[7:6] == 2'h1 ? ram_3_9 : _GEN_743; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_904 = _GEN_205[7:6] == 2'h1 ? ram_3_10 : _GEN_744; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_905 = _GEN_205[7:6] == 2'h1 ? ram_3_11 : _GEN_745; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_906 = _GEN_205[7:6] == 2'h1 ? ram_3_12 : _GEN_746; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_907 = _GEN_205[7:6] == 2'h1 ? ram_3_13 : _GEN_747; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_908 = _GEN_205[7:6] == 2'h1 ? ram_3_14 : _GEN_748; // @[i_cache.scala 115:52 22:24]
  wire [127:0] _GEN_909 = _GEN_205[7:6] == 2'h1 ? ram_3_15 : _GEN_749; // @[i_cache.scala 115:52 22:24]
  wire [31:0] _GEN_910 = _GEN_205[7:6] == 2'h1 ? tag_3_0 : _GEN_750; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_911 = _GEN_205[7:6] == 2'h1 ? tag_3_1 : _GEN_751; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_912 = _GEN_205[7:6] == 2'h1 ? tag_3_2 : _GEN_752; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_913 = _GEN_205[7:6] == 2'h1 ? tag_3_3 : _GEN_753; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_914 = _GEN_205[7:6] == 2'h1 ? tag_3_4 : _GEN_754; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_915 = _GEN_205[7:6] == 2'h1 ? tag_3_5 : _GEN_755; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_916 = _GEN_205[7:6] == 2'h1 ? tag_3_6 : _GEN_756; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_917 = _GEN_205[7:6] == 2'h1 ? tag_3_7 : _GEN_757; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_918 = _GEN_205[7:6] == 2'h1 ? tag_3_8 : _GEN_758; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_919 = _GEN_205[7:6] == 2'h1 ? tag_3_9 : _GEN_759; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_920 = _GEN_205[7:6] == 2'h1 ? tag_3_10 : _GEN_760; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_921 = _GEN_205[7:6] == 2'h1 ? tag_3_11 : _GEN_761; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_922 = _GEN_205[7:6] == 2'h1 ? tag_3_12 : _GEN_762; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_923 = _GEN_205[7:6] == 2'h1 ? tag_3_13 : _GEN_763; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_924 = _GEN_205[7:6] == 2'h1 ? tag_3_14 : _GEN_764; // @[i_cache.scala 115:52 26:24]
  wire [31:0] _GEN_925 = _GEN_205[7:6] == 2'h1 ? tag_3_15 : _GEN_765; // @[i_cache.scala 115:52 26:24]
  wire  _GEN_926 = _GEN_205[7:6] == 2'h1 ? valid_3_0 : _GEN_766; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_927 = _GEN_205[7:6] == 2'h1 ? valid_3_1 : _GEN_767; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_928 = _GEN_205[7:6] == 2'h1 ? valid_3_2 : _GEN_768; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_929 = _GEN_205[7:6] == 2'h1 ? valid_3_3 : _GEN_769; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_930 = _GEN_205[7:6] == 2'h1 ? valid_3_4 : _GEN_770; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_931 = _GEN_205[7:6] == 2'h1 ? valid_3_5 : _GEN_771; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_932 = _GEN_205[7:6] == 2'h1 ? valid_3_6 : _GEN_772; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_933 = _GEN_205[7:6] == 2'h1 ? valid_3_7 : _GEN_773; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_934 = _GEN_205[7:6] == 2'h1 ? valid_3_8 : _GEN_774; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_935 = _GEN_205[7:6] == 2'h1 ? valid_3_9 : _GEN_775; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_936 = _GEN_205[7:6] == 2'h1 ? valid_3_10 : _GEN_776; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_937 = _GEN_205[7:6] == 2'h1 ? valid_3_11 : _GEN_777; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_938 = _GEN_205[7:6] == 2'h1 ? valid_3_12 : _GEN_778; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_939 = _GEN_205[7:6] == 2'h1 ? valid_3_13 : _GEN_779; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_940 = _GEN_205[7:6] == 2'h1 ? valid_3_14 : _GEN_780; // @[i_cache.scala 115:52 30:26]
  wire  _GEN_941 = _GEN_205[7:6] == 2'h1 ? valid_3_15 : _GEN_781; // @[i_cache.scala 115:52 30:26]
  wire [127:0] _GEN_942 = _GEN_205[7:6] == 2'h0 ? _GEN_142 : ram_0_0; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_943 = _GEN_205[7:6] == 2'h0 ? _GEN_143 : ram_0_1; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_944 = _GEN_205[7:6] == 2'h0 ? _GEN_144 : ram_0_2; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_945 = _GEN_205[7:6] == 2'h0 ? _GEN_145 : ram_0_3; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_946 = _GEN_205[7:6] == 2'h0 ? _GEN_146 : ram_0_4; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_947 = _GEN_205[7:6] == 2'h0 ? _GEN_147 : ram_0_5; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_948 = _GEN_205[7:6] == 2'h0 ? _GEN_148 : ram_0_6; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_949 = _GEN_205[7:6] == 2'h0 ? _GEN_149 : ram_0_7; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_950 = _GEN_205[7:6] == 2'h0 ? _GEN_150 : ram_0_8; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_951 = _GEN_205[7:6] == 2'h0 ? _GEN_151 : ram_0_9; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_952 = _GEN_205[7:6] == 2'h0 ? _GEN_152 : ram_0_10; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_953 = _GEN_205[7:6] == 2'h0 ? _GEN_153 : ram_0_11; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_954 = _GEN_205[7:6] == 2'h0 ? _GEN_154 : ram_0_12; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_955 = _GEN_205[7:6] == 2'h0 ? _GEN_155 : ram_0_13; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_956 = _GEN_205[7:6] == 2'h0 ? _GEN_156 : ram_0_14; // @[i_cache.scala 110:46 19:24]
  wire [127:0] _GEN_957 = _GEN_205[7:6] == 2'h0 ? _GEN_157 : ram_0_15; // @[i_cache.scala 110:46 19:24]
  wire [31:0] _GEN_958 = _GEN_205[7:6] == 2'h0 ? _GEN_158 : tag_0_0; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_959 = _GEN_205[7:6] == 2'h0 ? _GEN_159 : tag_0_1; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_960 = _GEN_205[7:6] == 2'h0 ? _GEN_160 : tag_0_2; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_961 = _GEN_205[7:6] == 2'h0 ? _GEN_161 : tag_0_3; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_962 = _GEN_205[7:6] == 2'h0 ? _GEN_162 : tag_0_4; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_963 = _GEN_205[7:6] == 2'h0 ? _GEN_163 : tag_0_5; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_964 = _GEN_205[7:6] == 2'h0 ? _GEN_164 : tag_0_6; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_965 = _GEN_205[7:6] == 2'h0 ? _GEN_165 : tag_0_7; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_966 = _GEN_205[7:6] == 2'h0 ? _GEN_166 : tag_0_8; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_967 = _GEN_205[7:6] == 2'h0 ? _GEN_167 : tag_0_9; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_968 = _GEN_205[7:6] == 2'h0 ? _GEN_168 : tag_0_10; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_969 = _GEN_205[7:6] == 2'h0 ? _GEN_169 : tag_0_11; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_970 = _GEN_205[7:6] == 2'h0 ? _GEN_170 : tag_0_12; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_971 = _GEN_205[7:6] == 2'h0 ? _GEN_171 : tag_0_13; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_972 = _GEN_205[7:6] == 2'h0 ? _GEN_172 : tag_0_14; // @[i_cache.scala 110:46 23:24]
  wire [31:0] _GEN_973 = _GEN_205[7:6] == 2'h0 ? _GEN_173 : tag_0_15; // @[i_cache.scala 110:46 23:24]
  wire  _GEN_974 = _GEN_205[7:6] == 2'h0 ? _GEN_174 : valid_0_0; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_975 = _GEN_205[7:6] == 2'h0 ? _GEN_175 : valid_0_1; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_976 = _GEN_205[7:6] == 2'h0 ? _GEN_176 : valid_0_2; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_977 = _GEN_205[7:6] == 2'h0 ? _GEN_177 : valid_0_3; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_978 = _GEN_205[7:6] == 2'h0 ? _GEN_178 : valid_0_4; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_979 = _GEN_205[7:6] == 2'h0 ? _GEN_179 : valid_0_5; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_980 = _GEN_205[7:6] == 2'h0 ? _GEN_180 : valid_0_6; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_981 = _GEN_205[7:6] == 2'h0 ? _GEN_181 : valid_0_7; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_982 = _GEN_205[7:6] == 2'h0 ? _GEN_182 : valid_0_8; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_983 = _GEN_205[7:6] == 2'h0 ? _GEN_183 : valid_0_9; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_984 = _GEN_205[7:6] == 2'h0 ? _GEN_184 : valid_0_10; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_985 = _GEN_205[7:6] == 2'h0 ? _GEN_185 : valid_0_11; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_986 = _GEN_205[7:6] == 2'h0 ? _GEN_186 : valid_0_12; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_987 = _GEN_205[7:6] == 2'h0 ? _GEN_187 : valid_0_13; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_988 = _GEN_205[7:6] == 2'h0 ? _GEN_188 : valid_0_14; // @[i_cache.scala 110:46 27:26]
  wire  _GEN_989 = _GEN_205[7:6] == 2'h0 ? _GEN_189 : valid_0_15; // @[i_cache.scala 110:46 27:26]
  wire [7:0] _GEN_990 = _GEN_205[7:6] == 2'h0 ? _GEN_206 : _GEN_830; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_991 = _GEN_205[7:6] == 2'h0 ? _GEN_207 : _GEN_831; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_992 = _GEN_205[7:6] == 2'h0 ? _GEN_208 : _GEN_832; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_993 = _GEN_205[7:6] == 2'h0 ? _GEN_209 : _GEN_833; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_994 = _GEN_205[7:6] == 2'h0 ? _GEN_210 : _GEN_834; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_995 = _GEN_205[7:6] == 2'h0 ? _GEN_211 : _GEN_835; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_996 = _GEN_205[7:6] == 2'h0 ? _GEN_212 : _GEN_836; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_997 = _GEN_205[7:6] == 2'h0 ? _GEN_213 : _GEN_837; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_998 = _GEN_205[7:6] == 2'h0 ? _GEN_214 : _GEN_838; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_999 = _GEN_205[7:6] == 2'h0 ? _GEN_215 : _GEN_839; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_1000 = _GEN_205[7:6] == 2'h0 ? _GEN_216 : _GEN_840; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_1001 = _GEN_205[7:6] == 2'h0 ? _GEN_217 : _GEN_841; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_1002 = _GEN_205[7:6] == 2'h0 ? _GEN_218 : _GEN_842; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_1003 = _GEN_205[7:6] == 2'h0 ? _GEN_219 : _GEN_843; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_1004 = _GEN_205[7:6] == 2'h0 ? _GEN_220 : _GEN_844; // @[i_cache.scala 110:46]
  wire [7:0] _GEN_1005 = _GEN_205[7:6] == 2'h0 ? _GEN_221 : _GEN_845; // @[i_cache.scala 110:46]
  wire [127:0] _GEN_1006 = _GEN_205[7:6] == 2'h0 ? ram_1_0 : _GEN_782; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1007 = _GEN_205[7:6] == 2'h0 ? ram_1_1 : _GEN_783; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1008 = _GEN_205[7:6] == 2'h0 ? ram_1_2 : _GEN_784; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1009 = _GEN_205[7:6] == 2'h0 ? ram_1_3 : _GEN_785; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1010 = _GEN_205[7:6] == 2'h0 ? ram_1_4 : _GEN_786; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1011 = _GEN_205[7:6] == 2'h0 ? ram_1_5 : _GEN_787; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1012 = _GEN_205[7:6] == 2'h0 ? ram_1_6 : _GEN_788; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1013 = _GEN_205[7:6] == 2'h0 ? ram_1_7 : _GEN_789; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1014 = _GEN_205[7:6] == 2'h0 ? ram_1_8 : _GEN_790; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1015 = _GEN_205[7:6] == 2'h0 ? ram_1_9 : _GEN_791; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1016 = _GEN_205[7:6] == 2'h0 ? ram_1_10 : _GEN_792; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1017 = _GEN_205[7:6] == 2'h0 ? ram_1_11 : _GEN_793; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1018 = _GEN_205[7:6] == 2'h0 ? ram_1_12 : _GEN_794; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1019 = _GEN_205[7:6] == 2'h0 ? ram_1_13 : _GEN_795; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1020 = _GEN_205[7:6] == 2'h0 ? ram_1_14 : _GEN_796; // @[i_cache.scala 110:46 20:24]
  wire [127:0] _GEN_1021 = _GEN_205[7:6] == 2'h0 ? ram_1_15 : _GEN_797; // @[i_cache.scala 110:46 20:24]
  wire [31:0] _GEN_1022 = _GEN_205[7:6] == 2'h0 ? tag_1_0 : _GEN_798; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1023 = _GEN_205[7:6] == 2'h0 ? tag_1_1 : _GEN_799; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1024 = _GEN_205[7:6] == 2'h0 ? tag_1_2 : _GEN_800; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1025 = _GEN_205[7:6] == 2'h0 ? tag_1_3 : _GEN_801; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1026 = _GEN_205[7:6] == 2'h0 ? tag_1_4 : _GEN_802; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1027 = _GEN_205[7:6] == 2'h0 ? tag_1_5 : _GEN_803; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1028 = _GEN_205[7:6] == 2'h0 ? tag_1_6 : _GEN_804; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1029 = _GEN_205[7:6] == 2'h0 ? tag_1_7 : _GEN_805; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1030 = _GEN_205[7:6] == 2'h0 ? tag_1_8 : _GEN_806; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1031 = _GEN_205[7:6] == 2'h0 ? tag_1_9 : _GEN_807; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1032 = _GEN_205[7:6] == 2'h0 ? tag_1_10 : _GEN_808; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1033 = _GEN_205[7:6] == 2'h0 ? tag_1_11 : _GEN_809; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1034 = _GEN_205[7:6] == 2'h0 ? tag_1_12 : _GEN_810; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1035 = _GEN_205[7:6] == 2'h0 ? tag_1_13 : _GEN_811; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1036 = _GEN_205[7:6] == 2'h0 ? tag_1_14 : _GEN_812; // @[i_cache.scala 110:46 24:24]
  wire [31:0] _GEN_1037 = _GEN_205[7:6] == 2'h0 ? tag_1_15 : _GEN_813; // @[i_cache.scala 110:46 24:24]
  wire  _GEN_1038 = _GEN_205[7:6] == 2'h0 ? valid_1_0 : _GEN_814; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1039 = _GEN_205[7:6] == 2'h0 ? valid_1_1 : _GEN_815; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1040 = _GEN_205[7:6] == 2'h0 ? valid_1_2 : _GEN_816; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1041 = _GEN_205[7:6] == 2'h0 ? valid_1_3 : _GEN_817; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1042 = _GEN_205[7:6] == 2'h0 ? valid_1_4 : _GEN_818; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1043 = _GEN_205[7:6] == 2'h0 ? valid_1_5 : _GEN_819; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1044 = _GEN_205[7:6] == 2'h0 ? valid_1_6 : _GEN_820; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1045 = _GEN_205[7:6] == 2'h0 ? valid_1_7 : _GEN_821; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1046 = _GEN_205[7:6] == 2'h0 ? valid_1_8 : _GEN_822; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1047 = _GEN_205[7:6] == 2'h0 ? valid_1_9 : _GEN_823; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1048 = _GEN_205[7:6] == 2'h0 ? valid_1_10 : _GEN_824; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1049 = _GEN_205[7:6] == 2'h0 ? valid_1_11 : _GEN_825; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1050 = _GEN_205[7:6] == 2'h0 ? valid_1_12 : _GEN_826; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1051 = _GEN_205[7:6] == 2'h0 ? valid_1_13 : _GEN_827; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1052 = _GEN_205[7:6] == 2'h0 ? valid_1_14 : _GEN_828; // @[i_cache.scala 110:46 28:26]
  wire  _GEN_1053 = _GEN_205[7:6] == 2'h0 ? valid_1_15 : _GEN_829; // @[i_cache.scala 110:46 28:26]
  wire [127:0] _GEN_1054 = _GEN_205[7:6] == 2'h0 ? ram_2_0 : _GEN_846; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1055 = _GEN_205[7:6] == 2'h0 ? ram_2_1 : _GEN_847; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1056 = _GEN_205[7:6] == 2'h0 ? ram_2_2 : _GEN_848; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1057 = _GEN_205[7:6] == 2'h0 ? ram_2_3 : _GEN_849; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1058 = _GEN_205[7:6] == 2'h0 ? ram_2_4 : _GEN_850; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1059 = _GEN_205[7:6] == 2'h0 ? ram_2_5 : _GEN_851; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1060 = _GEN_205[7:6] == 2'h0 ? ram_2_6 : _GEN_852; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1061 = _GEN_205[7:6] == 2'h0 ? ram_2_7 : _GEN_853; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1062 = _GEN_205[7:6] == 2'h0 ? ram_2_8 : _GEN_854; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1063 = _GEN_205[7:6] == 2'h0 ? ram_2_9 : _GEN_855; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1064 = _GEN_205[7:6] == 2'h0 ? ram_2_10 : _GEN_856; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1065 = _GEN_205[7:6] == 2'h0 ? ram_2_11 : _GEN_857; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1066 = _GEN_205[7:6] == 2'h0 ? ram_2_12 : _GEN_858; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1067 = _GEN_205[7:6] == 2'h0 ? ram_2_13 : _GEN_859; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1068 = _GEN_205[7:6] == 2'h0 ? ram_2_14 : _GEN_860; // @[i_cache.scala 110:46 21:24]
  wire [127:0] _GEN_1069 = _GEN_205[7:6] == 2'h0 ? ram_2_15 : _GEN_861; // @[i_cache.scala 110:46 21:24]
  wire [31:0] _GEN_1070 = _GEN_205[7:6] == 2'h0 ? tag_2_0 : _GEN_862; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1071 = _GEN_205[7:6] == 2'h0 ? tag_2_1 : _GEN_863; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1072 = _GEN_205[7:6] == 2'h0 ? tag_2_2 : _GEN_864; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1073 = _GEN_205[7:6] == 2'h0 ? tag_2_3 : _GEN_865; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1074 = _GEN_205[7:6] == 2'h0 ? tag_2_4 : _GEN_866; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1075 = _GEN_205[7:6] == 2'h0 ? tag_2_5 : _GEN_867; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1076 = _GEN_205[7:6] == 2'h0 ? tag_2_6 : _GEN_868; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1077 = _GEN_205[7:6] == 2'h0 ? tag_2_7 : _GEN_869; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1078 = _GEN_205[7:6] == 2'h0 ? tag_2_8 : _GEN_870; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1079 = _GEN_205[7:6] == 2'h0 ? tag_2_9 : _GEN_871; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1080 = _GEN_205[7:6] == 2'h0 ? tag_2_10 : _GEN_872; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1081 = _GEN_205[7:6] == 2'h0 ? tag_2_11 : _GEN_873; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1082 = _GEN_205[7:6] == 2'h0 ? tag_2_12 : _GEN_874; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1083 = _GEN_205[7:6] == 2'h0 ? tag_2_13 : _GEN_875; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1084 = _GEN_205[7:6] == 2'h0 ? tag_2_14 : _GEN_876; // @[i_cache.scala 110:46 25:24]
  wire [31:0] _GEN_1085 = _GEN_205[7:6] == 2'h0 ? tag_2_15 : _GEN_877; // @[i_cache.scala 110:46 25:24]
  wire  _GEN_1086 = _GEN_205[7:6] == 2'h0 ? valid_2_0 : _GEN_878; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1087 = _GEN_205[7:6] == 2'h0 ? valid_2_1 : _GEN_879; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1088 = _GEN_205[7:6] == 2'h0 ? valid_2_2 : _GEN_880; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1089 = _GEN_205[7:6] == 2'h0 ? valid_2_3 : _GEN_881; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1090 = _GEN_205[7:6] == 2'h0 ? valid_2_4 : _GEN_882; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1091 = _GEN_205[7:6] == 2'h0 ? valid_2_5 : _GEN_883; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1092 = _GEN_205[7:6] == 2'h0 ? valid_2_6 : _GEN_884; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1093 = _GEN_205[7:6] == 2'h0 ? valid_2_7 : _GEN_885; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1094 = _GEN_205[7:6] == 2'h0 ? valid_2_8 : _GEN_886; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1095 = _GEN_205[7:6] == 2'h0 ? valid_2_9 : _GEN_887; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1096 = _GEN_205[7:6] == 2'h0 ? valid_2_10 : _GEN_888; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1097 = _GEN_205[7:6] == 2'h0 ? valid_2_11 : _GEN_889; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1098 = _GEN_205[7:6] == 2'h0 ? valid_2_12 : _GEN_890; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1099 = _GEN_205[7:6] == 2'h0 ? valid_2_13 : _GEN_891; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1100 = _GEN_205[7:6] == 2'h0 ? valid_2_14 : _GEN_892; // @[i_cache.scala 110:46 29:26]
  wire  _GEN_1101 = _GEN_205[7:6] == 2'h0 ? valid_2_15 : _GEN_893; // @[i_cache.scala 110:46 29:26]
  wire [127:0] _GEN_1102 = _GEN_205[7:6] == 2'h0 ? ram_3_0 : _GEN_894; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1103 = _GEN_205[7:6] == 2'h0 ? ram_3_1 : _GEN_895; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1104 = _GEN_205[7:6] == 2'h0 ? ram_3_2 : _GEN_896; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1105 = _GEN_205[7:6] == 2'h0 ? ram_3_3 : _GEN_897; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1106 = _GEN_205[7:6] == 2'h0 ? ram_3_4 : _GEN_898; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1107 = _GEN_205[7:6] == 2'h0 ? ram_3_5 : _GEN_899; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1108 = _GEN_205[7:6] == 2'h0 ? ram_3_6 : _GEN_900; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1109 = _GEN_205[7:6] == 2'h0 ? ram_3_7 : _GEN_901; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1110 = _GEN_205[7:6] == 2'h0 ? ram_3_8 : _GEN_902; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1111 = _GEN_205[7:6] == 2'h0 ? ram_3_9 : _GEN_903; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1112 = _GEN_205[7:6] == 2'h0 ? ram_3_10 : _GEN_904; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1113 = _GEN_205[7:6] == 2'h0 ? ram_3_11 : _GEN_905; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1114 = _GEN_205[7:6] == 2'h0 ? ram_3_12 : _GEN_906; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1115 = _GEN_205[7:6] == 2'h0 ? ram_3_13 : _GEN_907; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1116 = _GEN_205[7:6] == 2'h0 ? ram_3_14 : _GEN_908; // @[i_cache.scala 110:46 22:24]
  wire [127:0] _GEN_1117 = _GEN_205[7:6] == 2'h0 ? ram_3_15 : _GEN_909; // @[i_cache.scala 110:46 22:24]
  wire [31:0] _GEN_1118 = _GEN_205[7:6] == 2'h0 ? tag_3_0 : _GEN_910; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1119 = _GEN_205[7:6] == 2'h0 ? tag_3_1 : _GEN_911; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1120 = _GEN_205[7:6] == 2'h0 ? tag_3_2 : _GEN_912; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1121 = _GEN_205[7:6] == 2'h0 ? tag_3_3 : _GEN_913; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1122 = _GEN_205[7:6] == 2'h0 ? tag_3_4 : _GEN_914; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1123 = _GEN_205[7:6] == 2'h0 ? tag_3_5 : _GEN_915; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1124 = _GEN_205[7:6] == 2'h0 ? tag_3_6 : _GEN_916; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1125 = _GEN_205[7:6] == 2'h0 ? tag_3_7 : _GEN_917; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1126 = _GEN_205[7:6] == 2'h0 ? tag_3_8 : _GEN_918; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1127 = _GEN_205[7:6] == 2'h0 ? tag_3_9 : _GEN_919; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1128 = _GEN_205[7:6] == 2'h0 ? tag_3_10 : _GEN_920; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1129 = _GEN_205[7:6] == 2'h0 ? tag_3_11 : _GEN_921; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1130 = _GEN_205[7:6] == 2'h0 ? tag_3_12 : _GEN_922; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1131 = _GEN_205[7:6] == 2'h0 ? tag_3_13 : _GEN_923; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1132 = _GEN_205[7:6] == 2'h0 ? tag_3_14 : _GEN_924; // @[i_cache.scala 110:46 26:24]
  wire [31:0] _GEN_1133 = _GEN_205[7:6] == 2'h0 ? tag_3_15 : _GEN_925; // @[i_cache.scala 110:46 26:24]
  wire  _GEN_1134 = _GEN_205[7:6] == 2'h0 ? valid_3_0 : _GEN_926; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1135 = _GEN_205[7:6] == 2'h0 ? valid_3_1 : _GEN_927; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1136 = _GEN_205[7:6] == 2'h0 ? valid_3_2 : _GEN_928; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1137 = _GEN_205[7:6] == 2'h0 ? valid_3_3 : _GEN_929; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1138 = _GEN_205[7:6] == 2'h0 ? valid_3_4 : _GEN_930; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1139 = _GEN_205[7:6] == 2'h0 ? valid_3_5 : _GEN_931; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1140 = _GEN_205[7:6] == 2'h0 ? valid_3_6 : _GEN_932; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1141 = _GEN_205[7:6] == 2'h0 ? valid_3_7 : _GEN_933; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1142 = _GEN_205[7:6] == 2'h0 ? valid_3_8 : _GEN_934; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1143 = _GEN_205[7:6] == 2'h0 ? valid_3_9 : _GEN_935; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1144 = _GEN_205[7:6] == 2'h0 ? valid_3_10 : _GEN_936; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1145 = _GEN_205[7:6] == 2'h0 ? valid_3_11 : _GEN_937; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1146 = _GEN_205[7:6] == 2'h0 ? valid_3_12 : _GEN_938; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1147 = _GEN_205[7:6] == 2'h0 ? valid_3_13 : _GEN_939; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1148 = _GEN_205[7:6] == 2'h0 ? valid_3_14 : _GEN_940; // @[i_cache.scala 110:46 30:26]
  wire  _GEN_1149 = _GEN_205[7:6] == 2'h0 ? valid_3_15 : _GEN_941; // @[i_cache.scala 110:46 30:26]
  wire [127:0] _GEN_1150 = unuse_way == 3'h4 ? _GEN_350 : _GEN_1102; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1151 = unuse_way == 3'h4 ? _GEN_351 : _GEN_1103; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1152 = unuse_way == 3'h4 ? _GEN_352 : _GEN_1104; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1153 = unuse_way == 3'h4 ? _GEN_353 : _GEN_1105; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1154 = unuse_way == 3'h4 ? _GEN_354 : _GEN_1106; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1155 = unuse_way == 3'h4 ? _GEN_355 : _GEN_1107; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1156 = unuse_way == 3'h4 ? _GEN_356 : _GEN_1108; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1157 = unuse_way == 3'h4 ? _GEN_357 : _GEN_1109; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1158 = unuse_way == 3'h4 ? _GEN_358 : _GEN_1110; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1159 = unuse_way == 3'h4 ? _GEN_359 : _GEN_1111; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1160 = unuse_way == 3'h4 ? _GEN_360 : _GEN_1112; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1161 = unuse_way == 3'h4 ? _GEN_361 : _GEN_1113; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1162 = unuse_way == 3'h4 ? _GEN_362 : _GEN_1114; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1163 = unuse_way == 3'h4 ? _GEN_363 : _GEN_1115; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1164 = unuse_way == 3'h4 ? _GEN_364 : _GEN_1116; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1165 = unuse_way == 3'h4 ? _GEN_365 : _GEN_1117; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1166 = unuse_way == 3'h4 ? _GEN_366 : _GEN_1118; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1167 = unuse_way == 3'h4 ? _GEN_367 : _GEN_1119; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1168 = unuse_way == 3'h4 ? _GEN_368 : _GEN_1120; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1169 = unuse_way == 3'h4 ? _GEN_369 : _GEN_1121; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1170 = unuse_way == 3'h4 ? _GEN_370 : _GEN_1122; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1171 = unuse_way == 3'h4 ? _GEN_371 : _GEN_1123; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1172 = unuse_way == 3'h4 ? _GEN_372 : _GEN_1124; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1173 = unuse_way == 3'h4 ? _GEN_373 : _GEN_1125; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1174 = unuse_way == 3'h4 ? _GEN_374 : _GEN_1126; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1175 = unuse_way == 3'h4 ? _GEN_375 : _GEN_1127; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1176 = unuse_way == 3'h4 ? _GEN_376 : _GEN_1128; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1177 = unuse_way == 3'h4 ? _GEN_377 : _GEN_1129; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1178 = unuse_way == 3'h4 ? _GEN_378 : _GEN_1130; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1179 = unuse_way == 3'h4 ? _GEN_379 : _GEN_1131; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1180 = unuse_way == 3'h4 ? _GEN_380 : _GEN_1132; // @[i_cache.scala 104:40]
  wire [31:0] _GEN_1181 = unuse_way == 3'h4 ? _GEN_381 : _GEN_1133; // @[i_cache.scala 104:40]
  wire  _GEN_1182 = unuse_way == 3'h4 ? _GEN_382 : _GEN_1134; // @[i_cache.scala 104:40]
  wire  _GEN_1183 = unuse_way == 3'h4 ? _GEN_383 : _GEN_1135; // @[i_cache.scala 104:40]
  wire  _GEN_1184 = unuse_way == 3'h4 ? _GEN_384 : _GEN_1136; // @[i_cache.scala 104:40]
  wire  _GEN_1185 = unuse_way == 3'h4 ? _GEN_385 : _GEN_1137; // @[i_cache.scala 104:40]
  wire  _GEN_1186 = unuse_way == 3'h4 ? _GEN_386 : _GEN_1138; // @[i_cache.scala 104:40]
  wire  _GEN_1187 = unuse_way == 3'h4 ? _GEN_387 : _GEN_1139; // @[i_cache.scala 104:40]
  wire  _GEN_1188 = unuse_way == 3'h4 ? _GEN_388 : _GEN_1140; // @[i_cache.scala 104:40]
  wire  _GEN_1189 = unuse_way == 3'h4 ? _GEN_389 : _GEN_1141; // @[i_cache.scala 104:40]
  wire  _GEN_1190 = unuse_way == 3'h4 ? _GEN_390 : _GEN_1142; // @[i_cache.scala 104:40]
  wire  _GEN_1191 = unuse_way == 3'h4 ? _GEN_391 : _GEN_1143; // @[i_cache.scala 104:40]
  wire  _GEN_1192 = unuse_way == 3'h4 ? _GEN_392 : _GEN_1144; // @[i_cache.scala 104:40]
  wire  _GEN_1193 = unuse_way == 3'h4 ? _GEN_393 : _GEN_1145; // @[i_cache.scala 104:40]
  wire  _GEN_1194 = unuse_way == 3'h4 ? _GEN_394 : _GEN_1146; // @[i_cache.scala 104:40]
  wire  _GEN_1195 = unuse_way == 3'h4 ? _GEN_395 : _GEN_1147; // @[i_cache.scala 104:40]
  wire  _GEN_1196 = unuse_way == 3'h4 ? _GEN_396 : _GEN_1148; // @[i_cache.scala 104:40]
  wire  _GEN_1197 = unuse_way == 3'h4 ? _GEN_397 : _GEN_1149; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1198 = unuse_way == 3'h4 ? _GEN_398 : _GEN_990; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1199 = unuse_way == 3'h4 ? _GEN_399 : _GEN_991; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1200 = unuse_way == 3'h4 ? _GEN_400 : _GEN_992; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1201 = unuse_way == 3'h4 ? _GEN_401 : _GEN_993; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1202 = unuse_way == 3'h4 ? _GEN_402 : _GEN_994; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1203 = unuse_way == 3'h4 ? _GEN_403 : _GEN_995; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1204 = unuse_way == 3'h4 ? _GEN_404 : _GEN_996; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1205 = unuse_way == 3'h4 ? _GEN_405 : _GEN_997; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1206 = unuse_way == 3'h4 ? _GEN_406 : _GEN_998; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1207 = unuse_way == 3'h4 ? _GEN_407 : _GEN_999; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1208 = unuse_way == 3'h4 ? _GEN_408 : _GEN_1000; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1209 = unuse_way == 3'h4 ? _GEN_409 : _GEN_1001; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1210 = unuse_way == 3'h4 ? _GEN_410 : _GEN_1002; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1211 = unuse_way == 3'h4 ? _GEN_411 : _GEN_1003; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1212 = unuse_way == 3'h4 ? _GEN_412 : _GEN_1004; // @[i_cache.scala 104:40]
  wire [7:0] _GEN_1213 = unuse_way == 3'h4 ? _GEN_413 : _GEN_1005; // @[i_cache.scala 104:40]
  wire [127:0] _GEN_1214 = unuse_way == 3'h4 ? ram_0_0 : _GEN_942; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1215 = unuse_way == 3'h4 ? ram_0_1 : _GEN_943; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1216 = unuse_way == 3'h4 ? ram_0_2 : _GEN_944; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1217 = unuse_way == 3'h4 ? ram_0_3 : _GEN_945; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1218 = unuse_way == 3'h4 ? ram_0_4 : _GEN_946; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1219 = unuse_way == 3'h4 ? ram_0_5 : _GEN_947; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1220 = unuse_way == 3'h4 ? ram_0_6 : _GEN_948; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1221 = unuse_way == 3'h4 ? ram_0_7 : _GEN_949; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1222 = unuse_way == 3'h4 ? ram_0_8 : _GEN_950; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1223 = unuse_way == 3'h4 ? ram_0_9 : _GEN_951; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1224 = unuse_way == 3'h4 ? ram_0_10 : _GEN_952; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1225 = unuse_way == 3'h4 ? ram_0_11 : _GEN_953; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1226 = unuse_way == 3'h4 ? ram_0_12 : _GEN_954; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1227 = unuse_way == 3'h4 ? ram_0_13 : _GEN_955; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1228 = unuse_way == 3'h4 ? ram_0_14 : _GEN_956; // @[i_cache.scala 104:40 19:24]
  wire [127:0] _GEN_1229 = unuse_way == 3'h4 ? ram_0_15 : _GEN_957; // @[i_cache.scala 104:40 19:24]
  wire [31:0] _GEN_1230 = unuse_way == 3'h4 ? tag_0_0 : _GEN_958; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1231 = unuse_way == 3'h4 ? tag_0_1 : _GEN_959; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1232 = unuse_way == 3'h4 ? tag_0_2 : _GEN_960; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1233 = unuse_way == 3'h4 ? tag_0_3 : _GEN_961; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1234 = unuse_way == 3'h4 ? tag_0_4 : _GEN_962; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1235 = unuse_way == 3'h4 ? tag_0_5 : _GEN_963; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1236 = unuse_way == 3'h4 ? tag_0_6 : _GEN_964; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1237 = unuse_way == 3'h4 ? tag_0_7 : _GEN_965; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1238 = unuse_way == 3'h4 ? tag_0_8 : _GEN_966; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1239 = unuse_way == 3'h4 ? tag_0_9 : _GEN_967; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1240 = unuse_way == 3'h4 ? tag_0_10 : _GEN_968; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1241 = unuse_way == 3'h4 ? tag_0_11 : _GEN_969; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1242 = unuse_way == 3'h4 ? tag_0_12 : _GEN_970; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1243 = unuse_way == 3'h4 ? tag_0_13 : _GEN_971; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1244 = unuse_way == 3'h4 ? tag_0_14 : _GEN_972; // @[i_cache.scala 104:40 23:24]
  wire [31:0] _GEN_1245 = unuse_way == 3'h4 ? tag_0_15 : _GEN_973; // @[i_cache.scala 104:40 23:24]
  wire  _GEN_1246 = unuse_way == 3'h4 ? valid_0_0 : _GEN_974; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1247 = unuse_way == 3'h4 ? valid_0_1 : _GEN_975; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1248 = unuse_way == 3'h4 ? valid_0_2 : _GEN_976; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1249 = unuse_way == 3'h4 ? valid_0_3 : _GEN_977; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1250 = unuse_way == 3'h4 ? valid_0_4 : _GEN_978; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1251 = unuse_way == 3'h4 ? valid_0_5 : _GEN_979; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1252 = unuse_way == 3'h4 ? valid_0_6 : _GEN_980; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1253 = unuse_way == 3'h4 ? valid_0_7 : _GEN_981; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1254 = unuse_way == 3'h4 ? valid_0_8 : _GEN_982; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1255 = unuse_way == 3'h4 ? valid_0_9 : _GEN_983; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1256 = unuse_way == 3'h4 ? valid_0_10 : _GEN_984; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1257 = unuse_way == 3'h4 ? valid_0_11 : _GEN_985; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1258 = unuse_way == 3'h4 ? valid_0_12 : _GEN_986; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1259 = unuse_way == 3'h4 ? valid_0_13 : _GEN_987; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1260 = unuse_way == 3'h4 ? valid_0_14 : _GEN_988; // @[i_cache.scala 104:40 27:26]
  wire  _GEN_1261 = unuse_way == 3'h4 ? valid_0_15 : _GEN_989; // @[i_cache.scala 104:40 27:26]
  wire [127:0] _GEN_1262 = unuse_way == 3'h4 ? ram_1_0 : _GEN_1006; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1263 = unuse_way == 3'h4 ? ram_1_1 : _GEN_1007; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1264 = unuse_way == 3'h4 ? ram_1_2 : _GEN_1008; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1265 = unuse_way == 3'h4 ? ram_1_3 : _GEN_1009; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1266 = unuse_way == 3'h4 ? ram_1_4 : _GEN_1010; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1267 = unuse_way == 3'h4 ? ram_1_5 : _GEN_1011; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1268 = unuse_way == 3'h4 ? ram_1_6 : _GEN_1012; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1269 = unuse_way == 3'h4 ? ram_1_7 : _GEN_1013; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1270 = unuse_way == 3'h4 ? ram_1_8 : _GEN_1014; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1271 = unuse_way == 3'h4 ? ram_1_9 : _GEN_1015; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1272 = unuse_way == 3'h4 ? ram_1_10 : _GEN_1016; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1273 = unuse_way == 3'h4 ? ram_1_11 : _GEN_1017; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1274 = unuse_way == 3'h4 ? ram_1_12 : _GEN_1018; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1275 = unuse_way == 3'h4 ? ram_1_13 : _GEN_1019; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1276 = unuse_way == 3'h4 ? ram_1_14 : _GEN_1020; // @[i_cache.scala 104:40 20:24]
  wire [127:0] _GEN_1277 = unuse_way == 3'h4 ? ram_1_15 : _GEN_1021; // @[i_cache.scala 104:40 20:24]
  wire [31:0] _GEN_1278 = unuse_way == 3'h4 ? tag_1_0 : _GEN_1022; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1279 = unuse_way == 3'h4 ? tag_1_1 : _GEN_1023; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1280 = unuse_way == 3'h4 ? tag_1_2 : _GEN_1024; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1281 = unuse_way == 3'h4 ? tag_1_3 : _GEN_1025; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1282 = unuse_way == 3'h4 ? tag_1_4 : _GEN_1026; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1283 = unuse_way == 3'h4 ? tag_1_5 : _GEN_1027; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1284 = unuse_way == 3'h4 ? tag_1_6 : _GEN_1028; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1285 = unuse_way == 3'h4 ? tag_1_7 : _GEN_1029; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1286 = unuse_way == 3'h4 ? tag_1_8 : _GEN_1030; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1287 = unuse_way == 3'h4 ? tag_1_9 : _GEN_1031; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1288 = unuse_way == 3'h4 ? tag_1_10 : _GEN_1032; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1289 = unuse_way == 3'h4 ? tag_1_11 : _GEN_1033; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1290 = unuse_way == 3'h4 ? tag_1_12 : _GEN_1034; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1291 = unuse_way == 3'h4 ? tag_1_13 : _GEN_1035; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1292 = unuse_way == 3'h4 ? tag_1_14 : _GEN_1036; // @[i_cache.scala 104:40 24:24]
  wire [31:0] _GEN_1293 = unuse_way == 3'h4 ? tag_1_15 : _GEN_1037; // @[i_cache.scala 104:40 24:24]
  wire  _GEN_1294 = unuse_way == 3'h4 ? valid_1_0 : _GEN_1038; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1295 = unuse_way == 3'h4 ? valid_1_1 : _GEN_1039; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1296 = unuse_way == 3'h4 ? valid_1_2 : _GEN_1040; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1297 = unuse_way == 3'h4 ? valid_1_3 : _GEN_1041; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1298 = unuse_way == 3'h4 ? valid_1_4 : _GEN_1042; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1299 = unuse_way == 3'h4 ? valid_1_5 : _GEN_1043; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1300 = unuse_way == 3'h4 ? valid_1_6 : _GEN_1044; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1301 = unuse_way == 3'h4 ? valid_1_7 : _GEN_1045; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1302 = unuse_way == 3'h4 ? valid_1_8 : _GEN_1046; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1303 = unuse_way == 3'h4 ? valid_1_9 : _GEN_1047; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1304 = unuse_way == 3'h4 ? valid_1_10 : _GEN_1048; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1305 = unuse_way == 3'h4 ? valid_1_11 : _GEN_1049; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1306 = unuse_way == 3'h4 ? valid_1_12 : _GEN_1050; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1307 = unuse_way == 3'h4 ? valid_1_13 : _GEN_1051; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1308 = unuse_way == 3'h4 ? valid_1_14 : _GEN_1052; // @[i_cache.scala 104:40 28:26]
  wire  _GEN_1309 = unuse_way == 3'h4 ? valid_1_15 : _GEN_1053; // @[i_cache.scala 104:40 28:26]
  wire [127:0] _GEN_1310 = unuse_way == 3'h4 ? ram_2_0 : _GEN_1054; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1311 = unuse_way == 3'h4 ? ram_2_1 : _GEN_1055; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1312 = unuse_way == 3'h4 ? ram_2_2 : _GEN_1056; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1313 = unuse_way == 3'h4 ? ram_2_3 : _GEN_1057; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1314 = unuse_way == 3'h4 ? ram_2_4 : _GEN_1058; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1315 = unuse_way == 3'h4 ? ram_2_5 : _GEN_1059; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1316 = unuse_way == 3'h4 ? ram_2_6 : _GEN_1060; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1317 = unuse_way == 3'h4 ? ram_2_7 : _GEN_1061; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1318 = unuse_way == 3'h4 ? ram_2_8 : _GEN_1062; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1319 = unuse_way == 3'h4 ? ram_2_9 : _GEN_1063; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1320 = unuse_way == 3'h4 ? ram_2_10 : _GEN_1064; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1321 = unuse_way == 3'h4 ? ram_2_11 : _GEN_1065; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1322 = unuse_way == 3'h4 ? ram_2_12 : _GEN_1066; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1323 = unuse_way == 3'h4 ? ram_2_13 : _GEN_1067; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1324 = unuse_way == 3'h4 ? ram_2_14 : _GEN_1068; // @[i_cache.scala 104:40 21:24]
  wire [127:0] _GEN_1325 = unuse_way == 3'h4 ? ram_2_15 : _GEN_1069; // @[i_cache.scala 104:40 21:24]
  wire [31:0] _GEN_1326 = unuse_way == 3'h4 ? tag_2_0 : _GEN_1070; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1327 = unuse_way == 3'h4 ? tag_2_1 : _GEN_1071; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1328 = unuse_way == 3'h4 ? tag_2_2 : _GEN_1072; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1329 = unuse_way == 3'h4 ? tag_2_3 : _GEN_1073; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1330 = unuse_way == 3'h4 ? tag_2_4 : _GEN_1074; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1331 = unuse_way == 3'h4 ? tag_2_5 : _GEN_1075; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1332 = unuse_way == 3'h4 ? tag_2_6 : _GEN_1076; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1333 = unuse_way == 3'h4 ? tag_2_7 : _GEN_1077; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1334 = unuse_way == 3'h4 ? tag_2_8 : _GEN_1078; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1335 = unuse_way == 3'h4 ? tag_2_9 : _GEN_1079; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1336 = unuse_way == 3'h4 ? tag_2_10 : _GEN_1080; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1337 = unuse_way == 3'h4 ? tag_2_11 : _GEN_1081; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1338 = unuse_way == 3'h4 ? tag_2_12 : _GEN_1082; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1339 = unuse_way == 3'h4 ? tag_2_13 : _GEN_1083; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1340 = unuse_way == 3'h4 ? tag_2_14 : _GEN_1084; // @[i_cache.scala 104:40 25:24]
  wire [31:0] _GEN_1341 = unuse_way == 3'h4 ? tag_2_15 : _GEN_1085; // @[i_cache.scala 104:40 25:24]
  wire  _GEN_1342 = unuse_way == 3'h4 ? valid_2_0 : _GEN_1086; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1343 = unuse_way == 3'h4 ? valid_2_1 : _GEN_1087; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1344 = unuse_way == 3'h4 ? valid_2_2 : _GEN_1088; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1345 = unuse_way == 3'h4 ? valid_2_3 : _GEN_1089; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1346 = unuse_way == 3'h4 ? valid_2_4 : _GEN_1090; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1347 = unuse_way == 3'h4 ? valid_2_5 : _GEN_1091; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1348 = unuse_way == 3'h4 ? valid_2_6 : _GEN_1092; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1349 = unuse_way == 3'h4 ? valid_2_7 : _GEN_1093; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1350 = unuse_way == 3'h4 ? valid_2_8 : _GEN_1094; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1351 = unuse_way == 3'h4 ? valid_2_9 : _GEN_1095; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1352 = unuse_way == 3'h4 ? valid_2_10 : _GEN_1096; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1353 = unuse_way == 3'h4 ? valid_2_11 : _GEN_1097; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1354 = unuse_way == 3'h4 ? valid_2_12 : _GEN_1098; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1355 = unuse_way == 3'h4 ? valid_2_13 : _GEN_1099; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1356 = unuse_way == 3'h4 ? valid_2_14 : _GEN_1100; // @[i_cache.scala 104:40 29:26]
  wire  _GEN_1357 = unuse_way == 3'h4 ? valid_2_15 : _GEN_1101; // @[i_cache.scala 104:40 29:26]
  wire [127:0] _GEN_1358 = unuse_way == 3'h3 ? _GEN_286 : _GEN_1310; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1359 = unuse_way == 3'h3 ? _GEN_287 : _GEN_1311; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1360 = unuse_way == 3'h3 ? _GEN_288 : _GEN_1312; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1361 = unuse_way == 3'h3 ? _GEN_289 : _GEN_1313; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1362 = unuse_way == 3'h3 ? _GEN_290 : _GEN_1314; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1363 = unuse_way == 3'h3 ? _GEN_291 : _GEN_1315; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1364 = unuse_way == 3'h3 ? _GEN_292 : _GEN_1316; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1365 = unuse_way == 3'h3 ? _GEN_293 : _GEN_1317; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1366 = unuse_way == 3'h3 ? _GEN_294 : _GEN_1318; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1367 = unuse_way == 3'h3 ? _GEN_295 : _GEN_1319; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1368 = unuse_way == 3'h3 ? _GEN_296 : _GEN_1320; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1369 = unuse_way == 3'h3 ? _GEN_297 : _GEN_1321; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1370 = unuse_way == 3'h3 ? _GEN_298 : _GEN_1322; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1371 = unuse_way == 3'h3 ? _GEN_299 : _GEN_1323; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1372 = unuse_way == 3'h3 ? _GEN_300 : _GEN_1324; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1373 = unuse_way == 3'h3 ? _GEN_301 : _GEN_1325; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1374 = unuse_way == 3'h3 ? _GEN_302 : _GEN_1326; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1375 = unuse_way == 3'h3 ? _GEN_303 : _GEN_1327; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1376 = unuse_way == 3'h3 ? _GEN_304 : _GEN_1328; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1377 = unuse_way == 3'h3 ? _GEN_305 : _GEN_1329; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1378 = unuse_way == 3'h3 ? _GEN_306 : _GEN_1330; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1379 = unuse_way == 3'h3 ? _GEN_307 : _GEN_1331; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1380 = unuse_way == 3'h3 ? _GEN_308 : _GEN_1332; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1381 = unuse_way == 3'h3 ? _GEN_309 : _GEN_1333; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1382 = unuse_way == 3'h3 ? _GEN_310 : _GEN_1334; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1383 = unuse_way == 3'h3 ? _GEN_311 : _GEN_1335; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1384 = unuse_way == 3'h3 ? _GEN_312 : _GEN_1336; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1385 = unuse_way == 3'h3 ? _GEN_313 : _GEN_1337; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1386 = unuse_way == 3'h3 ? _GEN_314 : _GEN_1338; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1387 = unuse_way == 3'h3 ? _GEN_315 : _GEN_1339; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1388 = unuse_way == 3'h3 ? _GEN_316 : _GEN_1340; // @[i_cache.scala 99:40]
  wire [31:0] _GEN_1389 = unuse_way == 3'h3 ? _GEN_317 : _GEN_1341; // @[i_cache.scala 99:40]
  wire  _GEN_1390 = unuse_way == 3'h3 ? _GEN_318 : _GEN_1342; // @[i_cache.scala 99:40]
  wire  _GEN_1391 = unuse_way == 3'h3 ? _GEN_319 : _GEN_1343; // @[i_cache.scala 99:40]
  wire  _GEN_1392 = unuse_way == 3'h3 ? _GEN_320 : _GEN_1344; // @[i_cache.scala 99:40]
  wire  _GEN_1393 = unuse_way == 3'h3 ? _GEN_321 : _GEN_1345; // @[i_cache.scala 99:40]
  wire  _GEN_1394 = unuse_way == 3'h3 ? _GEN_322 : _GEN_1346; // @[i_cache.scala 99:40]
  wire  _GEN_1395 = unuse_way == 3'h3 ? _GEN_323 : _GEN_1347; // @[i_cache.scala 99:40]
  wire  _GEN_1396 = unuse_way == 3'h3 ? _GEN_324 : _GEN_1348; // @[i_cache.scala 99:40]
  wire  _GEN_1397 = unuse_way == 3'h3 ? _GEN_325 : _GEN_1349; // @[i_cache.scala 99:40]
  wire  _GEN_1398 = unuse_way == 3'h3 ? _GEN_326 : _GEN_1350; // @[i_cache.scala 99:40]
  wire  _GEN_1399 = unuse_way == 3'h3 ? _GEN_327 : _GEN_1351; // @[i_cache.scala 99:40]
  wire  _GEN_1400 = unuse_way == 3'h3 ? _GEN_328 : _GEN_1352; // @[i_cache.scala 99:40]
  wire  _GEN_1401 = unuse_way == 3'h3 ? _GEN_329 : _GEN_1353; // @[i_cache.scala 99:40]
  wire  _GEN_1402 = unuse_way == 3'h3 ? _GEN_330 : _GEN_1354; // @[i_cache.scala 99:40]
  wire  _GEN_1403 = unuse_way == 3'h3 ? _GEN_331 : _GEN_1355; // @[i_cache.scala 99:40]
  wire  _GEN_1404 = unuse_way == 3'h3 ? _GEN_332 : _GEN_1356; // @[i_cache.scala 99:40]
  wire  _GEN_1405 = unuse_way == 3'h3 ? _GEN_333 : _GEN_1357; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1406 = unuse_way == 3'h3 ? _GEN_334 : _GEN_1198; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1407 = unuse_way == 3'h3 ? _GEN_335 : _GEN_1199; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1408 = unuse_way == 3'h3 ? _GEN_336 : _GEN_1200; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1409 = unuse_way == 3'h3 ? _GEN_337 : _GEN_1201; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1410 = unuse_way == 3'h3 ? _GEN_338 : _GEN_1202; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1411 = unuse_way == 3'h3 ? _GEN_339 : _GEN_1203; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1412 = unuse_way == 3'h3 ? _GEN_340 : _GEN_1204; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1413 = unuse_way == 3'h3 ? _GEN_341 : _GEN_1205; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1414 = unuse_way == 3'h3 ? _GEN_342 : _GEN_1206; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1415 = unuse_way == 3'h3 ? _GEN_343 : _GEN_1207; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1416 = unuse_way == 3'h3 ? _GEN_344 : _GEN_1208; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1417 = unuse_way == 3'h3 ? _GEN_345 : _GEN_1209; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1418 = unuse_way == 3'h3 ? _GEN_346 : _GEN_1210; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1419 = unuse_way == 3'h3 ? _GEN_347 : _GEN_1211; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1420 = unuse_way == 3'h3 ? _GEN_348 : _GEN_1212; // @[i_cache.scala 99:40]
  wire [7:0] _GEN_1421 = unuse_way == 3'h3 ? _GEN_349 : _GEN_1213; // @[i_cache.scala 99:40]
  wire [127:0] _GEN_1422 = unuse_way == 3'h3 ? ram_3_0 : _GEN_1150; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1423 = unuse_way == 3'h3 ? ram_3_1 : _GEN_1151; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1424 = unuse_way == 3'h3 ? ram_3_2 : _GEN_1152; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1425 = unuse_way == 3'h3 ? ram_3_3 : _GEN_1153; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1426 = unuse_way == 3'h3 ? ram_3_4 : _GEN_1154; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1427 = unuse_way == 3'h3 ? ram_3_5 : _GEN_1155; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1428 = unuse_way == 3'h3 ? ram_3_6 : _GEN_1156; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1429 = unuse_way == 3'h3 ? ram_3_7 : _GEN_1157; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1430 = unuse_way == 3'h3 ? ram_3_8 : _GEN_1158; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1431 = unuse_way == 3'h3 ? ram_3_9 : _GEN_1159; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1432 = unuse_way == 3'h3 ? ram_3_10 : _GEN_1160; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1433 = unuse_way == 3'h3 ? ram_3_11 : _GEN_1161; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1434 = unuse_way == 3'h3 ? ram_3_12 : _GEN_1162; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1435 = unuse_way == 3'h3 ? ram_3_13 : _GEN_1163; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1436 = unuse_way == 3'h3 ? ram_3_14 : _GEN_1164; // @[i_cache.scala 22:24 99:40]
  wire [127:0] _GEN_1437 = unuse_way == 3'h3 ? ram_3_15 : _GEN_1165; // @[i_cache.scala 22:24 99:40]
  wire [31:0] _GEN_1438 = unuse_way == 3'h3 ? tag_3_0 : _GEN_1166; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1439 = unuse_way == 3'h3 ? tag_3_1 : _GEN_1167; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1440 = unuse_way == 3'h3 ? tag_3_2 : _GEN_1168; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1441 = unuse_way == 3'h3 ? tag_3_3 : _GEN_1169; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1442 = unuse_way == 3'h3 ? tag_3_4 : _GEN_1170; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1443 = unuse_way == 3'h3 ? tag_3_5 : _GEN_1171; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1444 = unuse_way == 3'h3 ? tag_3_6 : _GEN_1172; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1445 = unuse_way == 3'h3 ? tag_3_7 : _GEN_1173; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1446 = unuse_way == 3'h3 ? tag_3_8 : _GEN_1174; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1447 = unuse_way == 3'h3 ? tag_3_9 : _GEN_1175; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1448 = unuse_way == 3'h3 ? tag_3_10 : _GEN_1176; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1449 = unuse_way == 3'h3 ? tag_3_11 : _GEN_1177; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1450 = unuse_way == 3'h3 ? tag_3_12 : _GEN_1178; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1451 = unuse_way == 3'h3 ? tag_3_13 : _GEN_1179; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1452 = unuse_way == 3'h3 ? tag_3_14 : _GEN_1180; // @[i_cache.scala 26:24 99:40]
  wire [31:0] _GEN_1453 = unuse_way == 3'h3 ? tag_3_15 : _GEN_1181; // @[i_cache.scala 26:24 99:40]
  wire  _GEN_1454 = unuse_way == 3'h3 ? valid_3_0 : _GEN_1182; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1455 = unuse_way == 3'h3 ? valid_3_1 : _GEN_1183; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1456 = unuse_way == 3'h3 ? valid_3_2 : _GEN_1184; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1457 = unuse_way == 3'h3 ? valid_3_3 : _GEN_1185; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1458 = unuse_way == 3'h3 ? valid_3_4 : _GEN_1186; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1459 = unuse_way == 3'h3 ? valid_3_5 : _GEN_1187; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1460 = unuse_way == 3'h3 ? valid_3_6 : _GEN_1188; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1461 = unuse_way == 3'h3 ? valid_3_7 : _GEN_1189; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1462 = unuse_way == 3'h3 ? valid_3_8 : _GEN_1190; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1463 = unuse_way == 3'h3 ? valid_3_9 : _GEN_1191; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1464 = unuse_way == 3'h3 ? valid_3_10 : _GEN_1192; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1465 = unuse_way == 3'h3 ? valid_3_11 : _GEN_1193; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1466 = unuse_way == 3'h3 ? valid_3_12 : _GEN_1194; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1467 = unuse_way == 3'h3 ? valid_3_13 : _GEN_1195; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1468 = unuse_way == 3'h3 ? valid_3_14 : _GEN_1196; // @[i_cache.scala 30:26 99:40]
  wire  _GEN_1469 = unuse_way == 3'h3 ? valid_3_15 : _GEN_1197; // @[i_cache.scala 30:26 99:40]
  wire [127:0] _GEN_1470 = unuse_way == 3'h3 ? ram_0_0 : _GEN_1214; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1471 = unuse_way == 3'h3 ? ram_0_1 : _GEN_1215; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1472 = unuse_way == 3'h3 ? ram_0_2 : _GEN_1216; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1473 = unuse_way == 3'h3 ? ram_0_3 : _GEN_1217; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1474 = unuse_way == 3'h3 ? ram_0_4 : _GEN_1218; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1475 = unuse_way == 3'h3 ? ram_0_5 : _GEN_1219; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1476 = unuse_way == 3'h3 ? ram_0_6 : _GEN_1220; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1477 = unuse_way == 3'h3 ? ram_0_7 : _GEN_1221; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1478 = unuse_way == 3'h3 ? ram_0_8 : _GEN_1222; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1479 = unuse_way == 3'h3 ? ram_0_9 : _GEN_1223; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1480 = unuse_way == 3'h3 ? ram_0_10 : _GEN_1224; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1481 = unuse_way == 3'h3 ? ram_0_11 : _GEN_1225; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1482 = unuse_way == 3'h3 ? ram_0_12 : _GEN_1226; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1483 = unuse_way == 3'h3 ? ram_0_13 : _GEN_1227; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1484 = unuse_way == 3'h3 ? ram_0_14 : _GEN_1228; // @[i_cache.scala 19:24 99:40]
  wire [127:0] _GEN_1485 = unuse_way == 3'h3 ? ram_0_15 : _GEN_1229; // @[i_cache.scala 19:24 99:40]
  wire [31:0] _GEN_1486 = unuse_way == 3'h3 ? tag_0_0 : _GEN_1230; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1487 = unuse_way == 3'h3 ? tag_0_1 : _GEN_1231; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1488 = unuse_way == 3'h3 ? tag_0_2 : _GEN_1232; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1489 = unuse_way == 3'h3 ? tag_0_3 : _GEN_1233; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1490 = unuse_way == 3'h3 ? tag_0_4 : _GEN_1234; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1491 = unuse_way == 3'h3 ? tag_0_5 : _GEN_1235; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1492 = unuse_way == 3'h3 ? tag_0_6 : _GEN_1236; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1493 = unuse_way == 3'h3 ? tag_0_7 : _GEN_1237; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1494 = unuse_way == 3'h3 ? tag_0_8 : _GEN_1238; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1495 = unuse_way == 3'h3 ? tag_0_9 : _GEN_1239; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1496 = unuse_way == 3'h3 ? tag_0_10 : _GEN_1240; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1497 = unuse_way == 3'h3 ? tag_0_11 : _GEN_1241; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1498 = unuse_way == 3'h3 ? tag_0_12 : _GEN_1242; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1499 = unuse_way == 3'h3 ? tag_0_13 : _GEN_1243; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1500 = unuse_way == 3'h3 ? tag_0_14 : _GEN_1244; // @[i_cache.scala 23:24 99:40]
  wire [31:0] _GEN_1501 = unuse_way == 3'h3 ? tag_0_15 : _GEN_1245; // @[i_cache.scala 23:24 99:40]
  wire  _GEN_1502 = unuse_way == 3'h3 ? valid_0_0 : _GEN_1246; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1503 = unuse_way == 3'h3 ? valid_0_1 : _GEN_1247; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1504 = unuse_way == 3'h3 ? valid_0_2 : _GEN_1248; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1505 = unuse_way == 3'h3 ? valid_0_3 : _GEN_1249; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1506 = unuse_way == 3'h3 ? valid_0_4 : _GEN_1250; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1507 = unuse_way == 3'h3 ? valid_0_5 : _GEN_1251; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1508 = unuse_way == 3'h3 ? valid_0_6 : _GEN_1252; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1509 = unuse_way == 3'h3 ? valid_0_7 : _GEN_1253; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1510 = unuse_way == 3'h3 ? valid_0_8 : _GEN_1254; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1511 = unuse_way == 3'h3 ? valid_0_9 : _GEN_1255; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1512 = unuse_way == 3'h3 ? valid_0_10 : _GEN_1256; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1513 = unuse_way == 3'h3 ? valid_0_11 : _GEN_1257; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1514 = unuse_way == 3'h3 ? valid_0_12 : _GEN_1258; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1515 = unuse_way == 3'h3 ? valid_0_13 : _GEN_1259; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1516 = unuse_way == 3'h3 ? valid_0_14 : _GEN_1260; // @[i_cache.scala 27:26 99:40]
  wire  _GEN_1517 = unuse_way == 3'h3 ? valid_0_15 : _GEN_1261; // @[i_cache.scala 27:26 99:40]
  wire [127:0] _GEN_1518 = unuse_way == 3'h3 ? ram_1_0 : _GEN_1262; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1519 = unuse_way == 3'h3 ? ram_1_1 : _GEN_1263; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1520 = unuse_way == 3'h3 ? ram_1_2 : _GEN_1264; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1521 = unuse_way == 3'h3 ? ram_1_3 : _GEN_1265; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1522 = unuse_way == 3'h3 ? ram_1_4 : _GEN_1266; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1523 = unuse_way == 3'h3 ? ram_1_5 : _GEN_1267; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1524 = unuse_way == 3'h3 ? ram_1_6 : _GEN_1268; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1525 = unuse_way == 3'h3 ? ram_1_7 : _GEN_1269; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1526 = unuse_way == 3'h3 ? ram_1_8 : _GEN_1270; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1527 = unuse_way == 3'h3 ? ram_1_9 : _GEN_1271; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1528 = unuse_way == 3'h3 ? ram_1_10 : _GEN_1272; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1529 = unuse_way == 3'h3 ? ram_1_11 : _GEN_1273; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1530 = unuse_way == 3'h3 ? ram_1_12 : _GEN_1274; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1531 = unuse_way == 3'h3 ? ram_1_13 : _GEN_1275; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1532 = unuse_way == 3'h3 ? ram_1_14 : _GEN_1276; // @[i_cache.scala 20:24 99:40]
  wire [127:0] _GEN_1533 = unuse_way == 3'h3 ? ram_1_15 : _GEN_1277; // @[i_cache.scala 20:24 99:40]
  wire [31:0] _GEN_1534 = unuse_way == 3'h3 ? tag_1_0 : _GEN_1278; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1535 = unuse_way == 3'h3 ? tag_1_1 : _GEN_1279; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1536 = unuse_way == 3'h3 ? tag_1_2 : _GEN_1280; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1537 = unuse_way == 3'h3 ? tag_1_3 : _GEN_1281; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1538 = unuse_way == 3'h3 ? tag_1_4 : _GEN_1282; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1539 = unuse_way == 3'h3 ? tag_1_5 : _GEN_1283; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1540 = unuse_way == 3'h3 ? tag_1_6 : _GEN_1284; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1541 = unuse_way == 3'h3 ? tag_1_7 : _GEN_1285; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1542 = unuse_way == 3'h3 ? tag_1_8 : _GEN_1286; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1543 = unuse_way == 3'h3 ? tag_1_9 : _GEN_1287; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1544 = unuse_way == 3'h3 ? tag_1_10 : _GEN_1288; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1545 = unuse_way == 3'h3 ? tag_1_11 : _GEN_1289; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1546 = unuse_way == 3'h3 ? tag_1_12 : _GEN_1290; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1547 = unuse_way == 3'h3 ? tag_1_13 : _GEN_1291; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1548 = unuse_way == 3'h3 ? tag_1_14 : _GEN_1292; // @[i_cache.scala 24:24 99:40]
  wire [31:0] _GEN_1549 = unuse_way == 3'h3 ? tag_1_15 : _GEN_1293; // @[i_cache.scala 24:24 99:40]
  wire  _GEN_1550 = unuse_way == 3'h3 ? valid_1_0 : _GEN_1294; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1551 = unuse_way == 3'h3 ? valid_1_1 : _GEN_1295; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1552 = unuse_way == 3'h3 ? valid_1_2 : _GEN_1296; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1553 = unuse_way == 3'h3 ? valid_1_3 : _GEN_1297; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1554 = unuse_way == 3'h3 ? valid_1_4 : _GEN_1298; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1555 = unuse_way == 3'h3 ? valid_1_5 : _GEN_1299; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1556 = unuse_way == 3'h3 ? valid_1_6 : _GEN_1300; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1557 = unuse_way == 3'h3 ? valid_1_7 : _GEN_1301; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1558 = unuse_way == 3'h3 ? valid_1_8 : _GEN_1302; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1559 = unuse_way == 3'h3 ? valid_1_9 : _GEN_1303; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1560 = unuse_way == 3'h3 ? valid_1_10 : _GEN_1304; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1561 = unuse_way == 3'h3 ? valid_1_11 : _GEN_1305; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1562 = unuse_way == 3'h3 ? valid_1_12 : _GEN_1306; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1563 = unuse_way == 3'h3 ? valid_1_13 : _GEN_1307; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1564 = unuse_way == 3'h3 ? valid_1_14 : _GEN_1308; // @[i_cache.scala 28:26 99:40]
  wire  _GEN_1565 = unuse_way == 3'h3 ? valid_1_15 : _GEN_1309; // @[i_cache.scala 28:26 99:40]
  wire [127:0] _GEN_1566 = unuse_way == 3'h2 ? _GEN_222 : _GEN_1518; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1567 = unuse_way == 3'h2 ? _GEN_223 : _GEN_1519; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1568 = unuse_way == 3'h2 ? _GEN_224 : _GEN_1520; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1569 = unuse_way == 3'h2 ? _GEN_225 : _GEN_1521; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1570 = unuse_way == 3'h2 ? _GEN_226 : _GEN_1522; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1571 = unuse_way == 3'h2 ? _GEN_227 : _GEN_1523; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1572 = unuse_way == 3'h2 ? _GEN_228 : _GEN_1524; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1573 = unuse_way == 3'h2 ? _GEN_229 : _GEN_1525; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1574 = unuse_way == 3'h2 ? _GEN_230 : _GEN_1526; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1575 = unuse_way == 3'h2 ? _GEN_231 : _GEN_1527; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1576 = unuse_way == 3'h2 ? _GEN_232 : _GEN_1528; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1577 = unuse_way == 3'h2 ? _GEN_233 : _GEN_1529; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1578 = unuse_way == 3'h2 ? _GEN_234 : _GEN_1530; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1579 = unuse_way == 3'h2 ? _GEN_235 : _GEN_1531; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1580 = unuse_way == 3'h2 ? _GEN_236 : _GEN_1532; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1581 = unuse_way == 3'h2 ? _GEN_237 : _GEN_1533; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1582 = unuse_way == 3'h2 ? _GEN_238 : _GEN_1534; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1583 = unuse_way == 3'h2 ? _GEN_239 : _GEN_1535; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1584 = unuse_way == 3'h2 ? _GEN_240 : _GEN_1536; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1585 = unuse_way == 3'h2 ? _GEN_241 : _GEN_1537; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1586 = unuse_way == 3'h2 ? _GEN_242 : _GEN_1538; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1587 = unuse_way == 3'h2 ? _GEN_243 : _GEN_1539; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1588 = unuse_way == 3'h2 ? _GEN_244 : _GEN_1540; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1589 = unuse_way == 3'h2 ? _GEN_245 : _GEN_1541; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1590 = unuse_way == 3'h2 ? _GEN_246 : _GEN_1542; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1591 = unuse_way == 3'h2 ? _GEN_247 : _GEN_1543; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1592 = unuse_way == 3'h2 ? _GEN_248 : _GEN_1544; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1593 = unuse_way == 3'h2 ? _GEN_249 : _GEN_1545; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1594 = unuse_way == 3'h2 ? _GEN_250 : _GEN_1546; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1595 = unuse_way == 3'h2 ? _GEN_251 : _GEN_1547; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1596 = unuse_way == 3'h2 ? _GEN_252 : _GEN_1548; // @[i_cache.scala 94:40]
  wire [31:0] _GEN_1597 = unuse_way == 3'h2 ? _GEN_253 : _GEN_1549; // @[i_cache.scala 94:40]
  wire  _GEN_1598 = unuse_way == 3'h2 ? _GEN_254 : _GEN_1550; // @[i_cache.scala 94:40]
  wire  _GEN_1599 = unuse_way == 3'h2 ? _GEN_255 : _GEN_1551; // @[i_cache.scala 94:40]
  wire  _GEN_1600 = unuse_way == 3'h2 ? _GEN_256 : _GEN_1552; // @[i_cache.scala 94:40]
  wire  _GEN_1601 = unuse_way == 3'h2 ? _GEN_257 : _GEN_1553; // @[i_cache.scala 94:40]
  wire  _GEN_1602 = unuse_way == 3'h2 ? _GEN_258 : _GEN_1554; // @[i_cache.scala 94:40]
  wire  _GEN_1603 = unuse_way == 3'h2 ? _GEN_259 : _GEN_1555; // @[i_cache.scala 94:40]
  wire  _GEN_1604 = unuse_way == 3'h2 ? _GEN_260 : _GEN_1556; // @[i_cache.scala 94:40]
  wire  _GEN_1605 = unuse_way == 3'h2 ? _GEN_261 : _GEN_1557; // @[i_cache.scala 94:40]
  wire  _GEN_1606 = unuse_way == 3'h2 ? _GEN_262 : _GEN_1558; // @[i_cache.scala 94:40]
  wire  _GEN_1607 = unuse_way == 3'h2 ? _GEN_263 : _GEN_1559; // @[i_cache.scala 94:40]
  wire  _GEN_1608 = unuse_way == 3'h2 ? _GEN_264 : _GEN_1560; // @[i_cache.scala 94:40]
  wire  _GEN_1609 = unuse_way == 3'h2 ? _GEN_265 : _GEN_1561; // @[i_cache.scala 94:40]
  wire  _GEN_1610 = unuse_way == 3'h2 ? _GEN_266 : _GEN_1562; // @[i_cache.scala 94:40]
  wire  _GEN_1611 = unuse_way == 3'h2 ? _GEN_267 : _GEN_1563; // @[i_cache.scala 94:40]
  wire  _GEN_1612 = unuse_way == 3'h2 ? _GEN_268 : _GEN_1564; // @[i_cache.scala 94:40]
  wire  _GEN_1613 = unuse_way == 3'h2 ? _GEN_269 : _GEN_1565; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1614 = unuse_way == 3'h2 ? _GEN_270 : _GEN_1406; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1615 = unuse_way == 3'h2 ? _GEN_271 : _GEN_1407; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1616 = unuse_way == 3'h2 ? _GEN_272 : _GEN_1408; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1617 = unuse_way == 3'h2 ? _GEN_273 : _GEN_1409; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1618 = unuse_way == 3'h2 ? _GEN_274 : _GEN_1410; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1619 = unuse_way == 3'h2 ? _GEN_275 : _GEN_1411; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1620 = unuse_way == 3'h2 ? _GEN_276 : _GEN_1412; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1621 = unuse_way == 3'h2 ? _GEN_277 : _GEN_1413; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1622 = unuse_way == 3'h2 ? _GEN_278 : _GEN_1414; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1623 = unuse_way == 3'h2 ? _GEN_279 : _GEN_1415; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1624 = unuse_way == 3'h2 ? _GEN_280 : _GEN_1416; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1625 = unuse_way == 3'h2 ? _GEN_281 : _GEN_1417; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1626 = unuse_way == 3'h2 ? _GEN_282 : _GEN_1418; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1627 = unuse_way == 3'h2 ? _GEN_283 : _GEN_1419; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1628 = unuse_way == 3'h2 ? _GEN_284 : _GEN_1420; // @[i_cache.scala 94:40]
  wire [7:0] _GEN_1629 = unuse_way == 3'h2 ? _GEN_285 : _GEN_1421; // @[i_cache.scala 94:40]
  wire [127:0] _GEN_1630 = unuse_way == 3'h2 ? ram_2_0 : _GEN_1358; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1631 = unuse_way == 3'h2 ? ram_2_1 : _GEN_1359; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1632 = unuse_way == 3'h2 ? ram_2_2 : _GEN_1360; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1633 = unuse_way == 3'h2 ? ram_2_3 : _GEN_1361; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1634 = unuse_way == 3'h2 ? ram_2_4 : _GEN_1362; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1635 = unuse_way == 3'h2 ? ram_2_5 : _GEN_1363; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1636 = unuse_way == 3'h2 ? ram_2_6 : _GEN_1364; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1637 = unuse_way == 3'h2 ? ram_2_7 : _GEN_1365; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1638 = unuse_way == 3'h2 ? ram_2_8 : _GEN_1366; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1639 = unuse_way == 3'h2 ? ram_2_9 : _GEN_1367; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1640 = unuse_way == 3'h2 ? ram_2_10 : _GEN_1368; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1641 = unuse_way == 3'h2 ? ram_2_11 : _GEN_1369; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1642 = unuse_way == 3'h2 ? ram_2_12 : _GEN_1370; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1643 = unuse_way == 3'h2 ? ram_2_13 : _GEN_1371; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1644 = unuse_way == 3'h2 ? ram_2_14 : _GEN_1372; // @[i_cache.scala 21:24 94:40]
  wire [127:0] _GEN_1645 = unuse_way == 3'h2 ? ram_2_15 : _GEN_1373; // @[i_cache.scala 21:24 94:40]
  wire [31:0] _GEN_1646 = unuse_way == 3'h2 ? tag_2_0 : _GEN_1374; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1647 = unuse_way == 3'h2 ? tag_2_1 : _GEN_1375; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1648 = unuse_way == 3'h2 ? tag_2_2 : _GEN_1376; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1649 = unuse_way == 3'h2 ? tag_2_3 : _GEN_1377; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1650 = unuse_way == 3'h2 ? tag_2_4 : _GEN_1378; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1651 = unuse_way == 3'h2 ? tag_2_5 : _GEN_1379; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1652 = unuse_way == 3'h2 ? tag_2_6 : _GEN_1380; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1653 = unuse_way == 3'h2 ? tag_2_7 : _GEN_1381; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1654 = unuse_way == 3'h2 ? tag_2_8 : _GEN_1382; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1655 = unuse_way == 3'h2 ? tag_2_9 : _GEN_1383; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1656 = unuse_way == 3'h2 ? tag_2_10 : _GEN_1384; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1657 = unuse_way == 3'h2 ? tag_2_11 : _GEN_1385; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1658 = unuse_way == 3'h2 ? tag_2_12 : _GEN_1386; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1659 = unuse_way == 3'h2 ? tag_2_13 : _GEN_1387; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1660 = unuse_way == 3'h2 ? tag_2_14 : _GEN_1388; // @[i_cache.scala 25:24 94:40]
  wire [31:0] _GEN_1661 = unuse_way == 3'h2 ? tag_2_15 : _GEN_1389; // @[i_cache.scala 25:24 94:40]
  wire  _GEN_1662 = unuse_way == 3'h2 ? valid_2_0 : _GEN_1390; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1663 = unuse_way == 3'h2 ? valid_2_1 : _GEN_1391; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1664 = unuse_way == 3'h2 ? valid_2_2 : _GEN_1392; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1665 = unuse_way == 3'h2 ? valid_2_3 : _GEN_1393; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1666 = unuse_way == 3'h2 ? valid_2_4 : _GEN_1394; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1667 = unuse_way == 3'h2 ? valid_2_5 : _GEN_1395; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1668 = unuse_way == 3'h2 ? valid_2_6 : _GEN_1396; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1669 = unuse_way == 3'h2 ? valid_2_7 : _GEN_1397; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1670 = unuse_way == 3'h2 ? valid_2_8 : _GEN_1398; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1671 = unuse_way == 3'h2 ? valid_2_9 : _GEN_1399; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1672 = unuse_way == 3'h2 ? valid_2_10 : _GEN_1400; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1673 = unuse_way == 3'h2 ? valid_2_11 : _GEN_1401; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1674 = unuse_way == 3'h2 ? valid_2_12 : _GEN_1402; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1675 = unuse_way == 3'h2 ? valid_2_13 : _GEN_1403; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1676 = unuse_way == 3'h2 ? valid_2_14 : _GEN_1404; // @[i_cache.scala 29:26 94:40]
  wire  _GEN_1677 = unuse_way == 3'h2 ? valid_2_15 : _GEN_1405; // @[i_cache.scala 29:26 94:40]
  wire [127:0] _GEN_1678 = unuse_way == 3'h2 ? ram_3_0 : _GEN_1422; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1679 = unuse_way == 3'h2 ? ram_3_1 : _GEN_1423; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1680 = unuse_way == 3'h2 ? ram_3_2 : _GEN_1424; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1681 = unuse_way == 3'h2 ? ram_3_3 : _GEN_1425; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1682 = unuse_way == 3'h2 ? ram_3_4 : _GEN_1426; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1683 = unuse_way == 3'h2 ? ram_3_5 : _GEN_1427; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1684 = unuse_way == 3'h2 ? ram_3_6 : _GEN_1428; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1685 = unuse_way == 3'h2 ? ram_3_7 : _GEN_1429; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1686 = unuse_way == 3'h2 ? ram_3_8 : _GEN_1430; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1687 = unuse_way == 3'h2 ? ram_3_9 : _GEN_1431; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1688 = unuse_way == 3'h2 ? ram_3_10 : _GEN_1432; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1689 = unuse_way == 3'h2 ? ram_3_11 : _GEN_1433; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1690 = unuse_way == 3'h2 ? ram_3_12 : _GEN_1434; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1691 = unuse_way == 3'h2 ? ram_3_13 : _GEN_1435; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1692 = unuse_way == 3'h2 ? ram_3_14 : _GEN_1436; // @[i_cache.scala 22:24 94:40]
  wire [127:0] _GEN_1693 = unuse_way == 3'h2 ? ram_3_15 : _GEN_1437; // @[i_cache.scala 22:24 94:40]
  wire [31:0] _GEN_1694 = unuse_way == 3'h2 ? tag_3_0 : _GEN_1438; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1695 = unuse_way == 3'h2 ? tag_3_1 : _GEN_1439; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1696 = unuse_way == 3'h2 ? tag_3_2 : _GEN_1440; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1697 = unuse_way == 3'h2 ? tag_3_3 : _GEN_1441; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1698 = unuse_way == 3'h2 ? tag_3_4 : _GEN_1442; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1699 = unuse_way == 3'h2 ? tag_3_5 : _GEN_1443; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1700 = unuse_way == 3'h2 ? tag_3_6 : _GEN_1444; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1701 = unuse_way == 3'h2 ? tag_3_7 : _GEN_1445; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1702 = unuse_way == 3'h2 ? tag_3_8 : _GEN_1446; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1703 = unuse_way == 3'h2 ? tag_3_9 : _GEN_1447; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1704 = unuse_way == 3'h2 ? tag_3_10 : _GEN_1448; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1705 = unuse_way == 3'h2 ? tag_3_11 : _GEN_1449; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1706 = unuse_way == 3'h2 ? tag_3_12 : _GEN_1450; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1707 = unuse_way == 3'h2 ? tag_3_13 : _GEN_1451; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1708 = unuse_way == 3'h2 ? tag_3_14 : _GEN_1452; // @[i_cache.scala 26:24 94:40]
  wire [31:0] _GEN_1709 = unuse_way == 3'h2 ? tag_3_15 : _GEN_1453; // @[i_cache.scala 26:24 94:40]
  wire  _GEN_1710 = unuse_way == 3'h2 ? valid_3_0 : _GEN_1454; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1711 = unuse_way == 3'h2 ? valid_3_1 : _GEN_1455; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1712 = unuse_way == 3'h2 ? valid_3_2 : _GEN_1456; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1713 = unuse_way == 3'h2 ? valid_3_3 : _GEN_1457; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1714 = unuse_way == 3'h2 ? valid_3_4 : _GEN_1458; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1715 = unuse_way == 3'h2 ? valid_3_5 : _GEN_1459; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1716 = unuse_way == 3'h2 ? valid_3_6 : _GEN_1460; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1717 = unuse_way == 3'h2 ? valid_3_7 : _GEN_1461; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1718 = unuse_way == 3'h2 ? valid_3_8 : _GEN_1462; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1719 = unuse_way == 3'h2 ? valid_3_9 : _GEN_1463; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1720 = unuse_way == 3'h2 ? valid_3_10 : _GEN_1464; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1721 = unuse_way == 3'h2 ? valid_3_11 : _GEN_1465; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1722 = unuse_way == 3'h2 ? valid_3_12 : _GEN_1466; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1723 = unuse_way == 3'h2 ? valid_3_13 : _GEN_1467; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1724 = unuse_way == 3'h2 ? valid_3_14 : _GEN_1468; // @[i_cache.scala 30:26 94:40]
  wire  _GEN_1725 = unuse_way == 3'h2 ? valid_3_15 : _GEN_1469; // @[i_cache.scala 30:26 94:40]
  wire [127:0] _GEN_1726 = unuse_way == 3'h2 ? ram_0_0 : _GEN_1470; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1727 = unuse_way == 3'h2 ? ram_0_1 : _GEN_1471; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1728 = unuse_way == 3'h2 ? ram_0_2 : _GEN_1472; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1729 = unuse_way == 3'h2 ? ram_0_3 : _GEN_1473; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1730 = unuse_way == 3'h2 ? ram_0_4 : _GEN_1474; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1731 = unuse_way == 3'h2 ? ram_0_5 : _GEN_1475; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1732 = unuse_way == 3'h2 ? ram_0_6 : _GEN_1476; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1733 = unuse_way == 3'h2 ? ram_0_7 : _GEN_1477; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1734 = unuse_way == 3'h2 ? ram_0_8 : _GEN_1478; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1735 = unuse_way == 3'h2 ? ram_0_9 : _GEN_1479; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1736 = unuse_way == 3'h2 ? ram_0_10 : _GEN_1480; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1737 = unuse_way == 3'h2 ? ram_0_11 : _GEN_1481; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1738 = unuse_way == 3'h2 ? ram_0_12 : _GEN_1482; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1739 = unuse_way == 3'h2 ? ram_0_13 : _GEN_1483; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1740 = unuse_way == 3'h2 ? ram_0_14 : _GEN_1484; // @[i_cache.scala 19:24 94:40]
  wire [127:0] _GEN_1741 = unuse_way == 3'h2 ? ram_0_15 : _GEN_1485; // @[i_cache.scala 19:24 94:40]
  wire [31:0] _GEN_1742 = unuse_way == 3'h2 ? tag_0_0 : _GEN_1486; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1743 = unuse_way == 3'h2 ? tag_0_1 : _GEN_1487; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1744 = unuse_way == 3'h2 ? tag_0_2 : _GEN_1488; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1745 = unuse_way == 3'h2 ? tag_0_3 : _GEN_1489; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1746 = unuse_way == 3'h2 ? tag_0_4 : _GEN_1490; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1747 = unuse_way == 3'h2 ? tag_0_5 : _GEN_1491; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1748 = unuse_way == 3'h2 ? tag_0_6 : _GEN_1492; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1749 = unuse_way == 3'h2 ? tag_0_7 : _GEN_1493; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1750 = unuse_way == 3'h2 ? tag_0_8 : _GEN_1494; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1751 = unuse_way == 3'h2 ? tag_0_9 : _GEN_1495; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1752 = unuse_way == 3'h2 ? tag_0_10 : _GEN_1496; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1753 = unuse_way == 3'h2 ? tag_0_11 : _GEN_1497; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1754 = unuse_way == 3'h2 ? tag_0_12 : _GEN_1498; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1755 = unuse_way == 3'h2 ? tag_0_13 : _GEN_1499; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1756 = unuse_way == 3'h2 ? tag_0_14 : _GEN_1500; // @[i_cache.scala 23:24 94:40]
  wire [31:0] _GEN_1757 = unuse_way == 3'h2 ? tag_0_15 : _GEN_1501; // @[i_cache.scala 23:24 94:40]
  wire  _GEN_1758 = unuse_way == 3'h2 ? valid_0_0 : _GEN_1502; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1759 = unuse_way == 3'h2 ? valid_0_1 : _GEN_1503; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1760 = unuse_way == 3'h2 ? valid_0_2 : _GEN_1504; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1761 = unuse_way == 3'h2 ? valid_0_3 : _GEN_1505; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1762 = unuse_way == 3'h2 ? valid_0_4 : _GEN_1506; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1763 = unuse_way == 3'h2 ? valid_0_5 : _GEN_1507; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1764 = unuse_way == 3'h2 ? valid_0_6 : _GEN_1508; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1765 = unuse_way == 3'h2 ? valid_0_7 : _GEN_1509; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1766 = unuse_way == 3'h2 ? valid_0_8 : _GEN_1510; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1767 = unuse_way == 3'h2 ? valid_0_9 : _GEN_1511; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1768 = unuse_way == 3'h2 ? valid_0_10 : _GEN_1512; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1769 = unuse_way == 3'h2 ? valid_0_11 : _GEN_1513; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1770 = unuse_way == 3'h2 ? valid_0_12 : _GEN_1514; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1771 = unuse_way == 3'h2 ? valid_0_13 : _GEN_1515; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1772 = unuse_way == 3'h2 ? valid_0_14 : _GEN_1516; // @[i_cache.scala 27:26 94:40]
  wire  _GEN_1773 = unuse_way == 3'h2 ? valid_0_15 : _GEN_1517; // @[i_cache.scala 27:26 94:40]
  wire [127:0] _GEN_1774 = unuse_way == 3'h1 ? _GEN_142 : _GEN_1726; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1775 = unuse_way == 3'h1 ? _GEN_143 : _GEN_1727; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1776 = unuse_way == 3'h1 ? _GEN_144 : _GEN_1728; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1777 = unuse_way == 3'h1 ? _GEN_145 : _GEN_1729; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1778 = unuse_way == 3'h1 ? _GEN_146 : _GEN_1730; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1779 = unuse_way == 3'h1 ? _GEN_147 : _GEN_1731; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1780 = unuse_way == 3'h1 ? _GEN_148 : _GEN_1732; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1781 = unuse_way == 3'h1 ? _GEN_149 : _GEN_1733; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1782 = unuse_way == 3'h1 ? _GEN_150 : _GEN_1734; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1783 = unuse_way == 3'h1 ? _GEN_151 : _GEN_1735; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1784 = unuse_way == 3'h1 ? _GEN_152 : _GEN_1736; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1785 = unuse_way == 3'h1 ? _GEN_153 : _GEN_1737; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1786 = unuse_way == 3'h1 ? _GEN_154 : _GEN_1738; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1787 = unuse_way == 3'h1 ? _GEN_155 : _GEN_1739; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1788 = unuse_way == 3'h1 ? _GEN_156 : _GEN_1740; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1789 = unuse_way == 3'h1 ? _GEN_157 : _GEN_1741; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1790 = unuse_way == 3'h1 ? _GEN_158 : _GEN_1742; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1791 = unuse_way == 3'h1 ? _GEN_159 : _GEN_1743; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1792 = unuse_way == 3'h1 ? _GEN_160 : _GEN_1744; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1793 = unuse_way == 3'h1 ? _GEN_161 : _GEN_1745; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1794 = unuse_way == 3'h1 ? _GEN_162 : _GEN_1746; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1795 = unuse_way == 3'h1 ? _GEN_163 : _GEN_1747; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1796 = unuse_way == 3'h1 ? _GEN_164 : _GEN_1748; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1797 = unuse_way == 3'h1 ? _GEN_165 : _GEN_1749; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1798 = unuse_way == 3'h1 ? _GEN_166 : _GEN_1750; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1799 = unuse_way == 3'h1 ? _GEN_167 : _GEN_1751; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1800 = unuse_way == 3'h1 ? _GEN_168 : _GEN_1752; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1801 = unuse_way == 3'h1 ? _GEN_169 : _GEN_1753; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1802 = unuse_way == 3'h1 ? _GEN_170 : _GEN_1754; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1803 = unuse_way == 3'h1 ? _GEN_171 : _GEN_1755; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1804 = unuse_way == 3'h1 ? _GEN_172 : _GEN_1756; // @[i_cache.scala 89:34]
  wire [31:0] _GEN_1805 = unuse_way == 3'h1 ? _GEN_173 : _GEN_1757; // @[i_cache.scala 89:34]
  wire  _GEN_1806 = unuse_way == 3'h1 ? _GEN_174 : _GEN_1758; // @[i_cache.scala 89:34]
  wire  _GEN_1807 = unuse_way == 3'h1 ? _GEN_175 : _GEN_1759; // @[i_cache.scala 89:34]
  wire  _GEN_1808 = unuse_way == 3'h1 ? _GEN_176 : _GEN_1760; // @[i_cache.scala 89:34]
  wire  _GEN_1809 = unuse_way == 3'h1 ? _GEN_177 : _GEN_1761; // @[i_cache.scala 89:34]
  wire  _GEN_1810 = unuse_way == 3'h1 ? _GEN_178 : _GEN_1762; // @[i_cache.scala 89:34]
  wire  _GEN_1811 = unuse_way == 3'h1 ? _GEN_179 : _GEN_1763; // @[i_cache.scala 89:34]
  wire  _GEN_1812 = unuse_way == 3'h1 ? _GEN_180 : _GEN_1764; // @[i_cache.scala 89:34]
  wire  _GEN_1813 = unuse_way == 3'h1 ? _GEN_181 : _GEN_1765; // @[i_cache.scala 89:34]
  wire  _GEN_1814 = unuse_way == 3'h1 ? _GEN_182 : _GEN_1766; // @[i_cache.scala 89:34]
  wire  _GEN_1815 = unuse_way == 3'h1 ? _GEN_183 : _GEN_1767; // @[i_cache.scala 89:34]
  wire  _GEN_1816 = unuse_way == 3'h1 ? _GEN_184 : _GEN_1768; // @[i_cache.scala 89:34]
  wire  _GEN_1817 = unuse_way == 3'h1 ? _GEN_185 : _GEN_1769; // @[i_cache.scala 89:34]
  wire  _GEN_1818 = unuse_way == 3'h1 ? _GEN_186 : _GEN_1770; // @[i_cache.scala 89:34]
  wire  _GEN_1819 = unuse_way == 3'h1 ? _GEN_187 : _GEN_1771; // @[i_cache.scala 89:34]
  wire  _GEN_1820 = unuse_way == 3'h1 ? _GEN_188 : _GEN_1772; // @[i_cache.scala 89:34]
  wire  _GEN_1821 = unuse_way == 3'h1 ? _GEN_189 : _GEN_1773; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1822 = unuse_way == 3'h1 ? _GEN_206 : _GEN_1614; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1823 = unuse_way == 3'h1 ? _GEN_207 : _GEN_1615; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1824 = unuse_way == 3'h1 ? _GEN_208 : _GEN_1616; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1825 = unuse_way == 3'h1 ? _GEN_209 : _GEN_1617; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1826 = unuse_way == 3'h1 ? _GEN_210 : _GEN_1618; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1827 = unuse_way == 3'h1 ? _GEN_211 : _GEN_1619; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1828 = unuse_way == 3'h1 ? _GEN_212 : _GEN_1620; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1829 = unuse_way == 3'h1 ? _GEN_213 : _GEN_1621; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1830 = unuse_way == 3'h1 ? _GEN_214 : _GEN_1622; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1831 = unuse_way == 3'h1 ? _GEN_215 : _GEN_1623; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1832 = unuse_way == 3'h1 ? _GEN_216 : _GEN_1624; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1833 = unuse_way == 3'h1 ? _GEN_217 : _GEN_1625; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1834 = unuse_way == 3'h1 ? _GEN_218 : _GEN_1626; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1835 = unuse_way == 3'h1 ? _GEN_219 : _GEN_1627; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1836 = unuse_way == 3'h1 ? _GEN_220 : _GEN_1628; // @[i_cache.scala 89:34]
  wire [7:0] _GEN_1837 = unuse_way == 3'h1 ? _GEN_221 : _GEN_1629; // @[i_cache.scala 89:34]
  wire [127:0] _GEN_1838 = unuse_way == 3'h1 ? ram_1_0 : _GEN_1566; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1839 = unuse_way == 3'h1 ? ram_1_1 : _GEN_1567; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1840 = unuse_way == 3'h1 ? ram_1_2 : _GEN_1568; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1841 = unuse_way == 3'h1 ? ram_1_3 : _GEN_1569; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1842 = unuse_way == 3'h1 ? ram_1_4 : _GEN_1570; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1843 = unuse_way == 3'h1 ? ram_1_5 : _GEN_1571; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1844 = unuse_way == 3'h1 ? ram_1_6 : _GEN_1572; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1845 = unuse_way == 3'h1 ? ram_1_7 : _GEN_1573; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1846 = unuse_way == 3'h1 ? ram_1_8 : _GEN_1574; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1847 = unuse_way == 3'h1 ? ram_1_9 : _GEN_1575; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1848 = unuse_way == 3'h1 ? ram_1_10 : _GEN_1576; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1849 = unuse_way == 3'h1 ? ram_1_11 : _GEN_1577; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1850 = unuse_way == 3'h1 ? ram_1_12 : _GEN_1578; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1851 = unuse_way == 3'h1 ? ram_1_13 : _GEN_1579; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1852 = unuse_way == 3'h1 ? ram_1_14 : _GEN_1580; // @[i_cache.scala 20:24 89:34]
  wire [127:0] _GEN_1853 = unuse_way == 3'h1 ? ram_1_15 : _GEN_1581; // @[i_cache.scala 20:24 89:34]
  wire [31:0] _GEN_1854 = unuse_way == 3'h1 ? tag_1_0 : _GEN_1582; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1855 = unuse_way == 3'h1 ? tag_1_1 : _GEN_1583; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1856 = unuse_way == 3'h1 ? tag_1_2 : _GEN_1584; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1857 = unuse_way == 3'h1 ? tag_1_3 : _GEN_1585; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1858 = unuse_way == 3'h1 ? tag_1_4 : _GEN_1586; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1859 = unuse_way == 3'h1 ? tag_1_5 : _GEN_1587; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1860 = unuse_way == 3'h1 ? tag_1_6 : _GEN_1588; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1861 = unuse_way == 3'h1 ? tag_1_7 : _GEN_1589; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1862 = unuse_way == 3'h1 ? tag_1_8 : _GEN_1590; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1863 = unuse_way == 3'h1 ? tag_1_9 : _GEN_1591; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1864 = unuse_way == 3'h1 ? tag_1_10 : _GEN_1592; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1865 = unuse_way == 3'h1 ? tag_1_11 : _GEN_1593; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1866 = unuse_way == 3'h1 ? tag_1_12 : _GEN_1594; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1867 = unuse_way == 3'h1 ? tag_1_13 : _GEN_1595; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1868 = unuse_way == 3'h1 ? tag_1_14 : _GEN_1596; // @[i_cache.scala 24:24 89:34]
  wire [31:0] _GEN_1869 = unuse_way == 3'h1 ? tag_1_15 : _GEN_1597; // @[i_cache.scala 24:24 89:34]
  wire  _GEN_1870 = unuse_way == 3'h1 ? valid_1_0 : _GEN_1598; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1871 = unuse_way == 3'h1 ? valid_1_1 : _GEN_1599; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1872 = unuse_way == 3'h1 ? valid_1_2 : _GEN_1600; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1873 = unuse_way == 3'h1 ? valid_1_3 : _GEN_1601; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1874 = unuse_way == 3'h1 ? valid_1_4 : _GEN_1602; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1875 = unuse_way == 3'h1 ? valid_1_5 : _GEN_1603; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1876 = unuse_way == 3'h1 ? valid_1_6 : _GEN_1604; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1877 = unuse_way == 3'h1 ? valid_1_7 : _GEN_1605; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1878 = unuse_way == 3'h1 ? valid_1_8 : _GEN_1606; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1879 = unuse_way == 3'h1 ? valid_1_9 : _GEN_1607; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1880 = unuse_way == 3'h1 ? valid_1_10 : _GEN_1608; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1881 = unuse_way == 3'h1 ? valid_1_11 : _GEN_1609; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1882 = unuse_way == 3'h1 ? valid_1_12 : _GEN_1610; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1883 = unuse_way == 3'h1 ? valid_1_13 : _GEN_1611; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1884 = unuse_way == 3'h1 ? valid_1_14 : _GEN_1612; // @[i_cache.scala 28:26 89:34]
  wire  _GEN_1885 = unuse_way == 3'h1 ? valid_1_15 : _GEN_1613; // @[i_cache.scala 28:26 89:34]
  wire [127:0] _GEN_1886 = unuse_way == 3'h1 ? ram_2_0 : _GEN_1630; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1887 = unuse_way == 3'h1 ? ram_2_1 : _GEN_1631; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1888 = unuse_way == 3'h1 ? ram_2_2 : _GEN_1632; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1889 = unuse_way == 3'h1 ? ram_2_3 : _GEN_1633; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1890 = unuse_way == 3'h1 ? ram_2_4 : _GEN_1634; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1891 = unuse_way == 3'h1 ? ram_2_5 : _GEN_1635; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1892 = unuse_way == 3'h1 ? ram_2_6 : _GEN_1636; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1893 = unuse_way == 3'h1 ? ram_2_7 : _GEN_1637; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1894 = unuse_way == 3'h1 ? ram_2_8 : _GEN_1638; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1895 = unuse_way == 3'h1 ? ram_2_9 : _GEN_1639; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1896 = unuse_way == 3'h1 ? ram_2_10 : _GEN_1640; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1897 = unuse_way == 3'h1 ? ram_2_11 : _GEN_1641; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1898 = unuse_way == 3'h1 ? ram_2_12 : _GEN_1642; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1899 = unuse_way == 3'h1 ? ram_2_13 : _GEN_1643; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1900 = unuse_way == 3'h1 ? ram_2_14 : _GEN_1644; // @[i_cache.scala 21:24 89:34]
  wire [127:0] _GEN_1901 = unuse_way == 3'h1 ? ram_2_15 : _GEN_1645; // @[i_cache.scala 21:24 89:34]
  wire [31:0] _GEN_1902 = unuse_way == 3'h1 ? tag_2_0 : _GEN_1646; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1903 = unuse_way == 3'h1 ? tag_2_1 : _GEN_1647; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1904 = unuse_way == 3'h1 ? tag_2_2 : _GEN_1648; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1905 = unuse_way == 3'h1 ? tag_2_3 : _GEN_1649; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1906 = unuse_way == 3'h1 ? tag_2_4 : _GEN_1650; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1907 = unuse_way == 3'h1 ? tag_2_5 : _GEN_1651; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1908 = unuse_way == 3'h1 ? tag_2_6 : _GEN_1652; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1909 = unuse_way == 3'h1 ? tag_2_7 : _GEN_1653; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1910 = unuse_way == 3'h1 ? tag_2_8 : _GEN_1654; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1911 = unuse_way == 3'h1 ? tag_2_9 : _GEN_1655; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1912 = unuse_way == 3'h1 ? tag_2_10 : _GEN_1656; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1913 = unuse_way == 3'h1 ? tag_2_11 : _GEN_1657; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1914 = unuse_way == 3'h1 ? tag_2_12 : _GEN_1658; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1915 = unuse_way == 3'h1 ? tag_2_13 : _GEN_1659; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1916 = unuse_way == 3'h1 ? tag_2_14 : _GEN_1660; // @[i_cache.scala 25:24 89:34]
  wire [31:0] _GEN_1917 = unuse_way == 3'h1 ? tag_2_15 : _GEN_1661; // @[i_cache.scala 25:24 89:34]
  wire  _GEN_1918 = unuse_way == 3'h1 ? valid_2_0 : _GEN_1662; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1919 = unuse_way == 3'h1 ? valid_2_1 : _GEN_1663; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1920 = unuse_way == 3'h1 ? valid_2_2 : _GEN_1664; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1921 = unuse_way == 3'h1 ? valid_2_3 : _GEN_1665; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1922 = unuse_way == 3'h1 ? valid_2_4 : _GEN_1666; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1923 = unuse_way == 3'h1 ? valid_2_5 : _GEN_1667; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1924 = unuse_way == 3'h1 ? valid_2_6 : _GEN_1668; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1925 = unuse_way == 3'h1 ? valid_2_7 : _GEN_1669; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1926 = unuse_way == 3'h1 ? valid_2_8 : _GEN_1670; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1927 = unuse_way == 3'h1 ? valid_2_9 : _GEN_1671; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1928 = unuse_way == 3'h1 ? valid_2_10 : _GEN_1672; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1929 = unuse_way == 3'h1 ? valid_2_11 : _GEN_1673; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1930 = unuse_way == 3'h1 ? valid_2_12 : _GEN_1674; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1931 = unuse_way == 3'h1 ? valid_2_13 : _GEN_1675; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1932 = unuse_way == 3'h1 ? valid_2_14 : _GEN_1676; // @[i_cache.scala 29:26 89:34]
  wire  _GEN_1933 = unuse_way == 3'h1 ? valid_2_15 : _GEN_1677; // @[i_cache.scala 29:26 89:34]
  wire [127:0] _GEN_1934 = unuse_way == 3'h1 ? ram_3_0 : _GEN_1678; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1935 = unuse_way == 3'h1 ? ram_3_1 : _GEN_1679; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1936 = unuse_way == 3'h1 ? ram_3_2 : _GEN_1680; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1937 = unuse_way == 3'h1 ? ram_3_3 : _GEN_1681; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1938 = unuse_way == 3'h1 ? ram_3_4 : _GEN_1682; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1939 = unuse_way == 3'h1 ? ram_3_5 : _GEN_1683; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1940 = unuse_way == 3'h1 ? ram_3_6 : _GEN_1684; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1941 = unuse_way == 3'h1 ? ram_3_7 : _GEN_1685; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1942 = unuse_way == 3'h1 ? ram_3_8 : _GEN_1686; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1943 = unuse_way == 3'h1 ? ram_3_9 : _GEN_1687; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1944 = unuse_way == 3'h1 ? ram_3_10 : _GEN_1688; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1945 = unuse_way == 3'h1 ? ram_3_11 : _GEN_1689; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1946 = unuse_way == 3'h1 ? ram_3_12 : _GEN_1690; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1947 = unuse_way == 3'h1 ? ram_3_13 : _GEN_1691; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1948 = unuse_way == 3'h1 ? ram_3_14 : _GEN_1692; // @[i_cache.scala 22:24 89:34]
  wire [127:0] _GEN_1949 = unuse_way == 3'h1 ? ram_3_15 : _GEN_1693; // @[i_cache.scala 22:24 89:34]
  wire [31:0] _GEN_1950 = unuse_way == 3'h1 ? tag_3_0 : _GEN_1694; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1951 = unuse_way == 3'h1 ? tag_3_1 : _GEN_1695; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1952 = unuse_way == 3'h1 ? tag_3_2 : _GEN_1696; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1953 = unuse_way == 3'h1 ? tag_3_3 : _GEN_1697; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1954 = unuse_way == 3'h1 ? tag_3_4 : _GEN_1698; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1955 = unuse_way == 3'h1 ? tag_3_5 : _GEN_1699; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1956 = unuse_way == 3'h1 ? tag_3_6 : _GEN_1700; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1957 = unuse_way == 3'h1 ? tag_3_7 : _GEN_1701; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1958 = unuse_way == 3'h1 ? tag_3_8 : _GEN_1702; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1959 = unuse_way == 3'h1 ? tag_3_9 : _GEN_1703; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1960 = unuse_way == 3'h1 ? tag_3_10 : _GEN_1704; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1961 = unuse_way == 3'h1 ? tag_3_11 : _GEN_1705; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1962 = unuse_way == 3'h1 ? tag_3_12 : _GEN_1706; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1963 = unuse_way == 3'h1 ? tag_3_13 : _GEN_1707; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1964 = unuse_way == 3'h1 ? tag_3_14 : _GEN_1708; // @[i_cache.scala 26:24 89:34]
  wire [31:0] _GEN_1965 = unuse_way == 3'h1 ? tag_3_15 : _GEN_1709; // @[i_cache.scala 26:24 89:34]
  wire  _GEN_1966 = unuse_way == 3'h1 ? valid_3_0 : _GEN_1710; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1967 = unuse_way == 3'h1 ? valid_3_1 : _GEN_1711; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1968 = unuse_way == 3'h1 ? valid_3_2 : _GEN_1712; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1969 = unuse_way == 3'h1 ? valid_3_3 : _GEN_1713; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1970 = unuse_way == 3'h1 ? valid_3_4 : _GEN_1714; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1971 = unuse_way == 3'h1 ? valid_3_5 : _GEN_1715; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1972 = unuse_way == 3'h1 ? valid_3_6 : _GEN_1716; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1973 = unuse_way == 3'h1 ? valid_3_7 : _GEN_1717; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1974 = unuse_way == 3'h1 ? valid_3_8 : _GEN_1718; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1975 = unuse_way == 3'h1 ? valid_3_9 : _GEN_1719; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1976 = unuse_way == 3'h1 ? valid_3_10 : _GEN_1720; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1977 = unuse_way == 3'h1 ? valid_3_11 : _GEN_1721; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1978 = unuse_way == 3'h1 ? valid_3_12 : _GEN_1722; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1979 = unuse_way == 3'h1 ? valid_3_13 : _GEN_1723; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1980 = unuse_way == 3'h1 ? valid_3_14 : _GEN_1724; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1981 = unuse_way == 3'h1 ? valid_3_15 : _GEN_1725; // @[i_cache.scala 30:26 89:34]
  wire  _GEN_1982 = 3'h4 == state ? 1'h0 : valid_0_0; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1983 = 3'h4 == state ? 1'h0 : valid_0_1; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1984 = 3'h4 == state ? 1'h0 : valid_0_2; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1985 = 3'h4 == state ? 1'h0 : valid_0_3; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1986 = 3'h4 == state ? 1'h0 : valid_0_4; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1987 = 3'h4 == state ? 1'h0 : valid_0_5; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1988 = 3'h4 == state ? 1'h0 : valid_0_6; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1989 = 3'h4 == state ? 1'h0 : valid_0_7; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1990 = 3'h4 == state ? 1'h0 : valid_0_8; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1991 = 3'h4 == state ? 1'h0 : valid_0_9; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1992 = 3'h4 == state ? 1'h0 : valid_0_10; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1993 = 3'h4 == state ? 1'h0 : valid_0_11; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1994 = 3'h4 == state ? 1'h0 : valid_0_12; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1995 = 3'h4 == state ? 1'h0 : valid_0_13; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1996 = 3'h4 == state ? 1'h0 : valid_0_14; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1997 = 3'h4 == state ? 1'h0 : valid_0_15; // @[i_cache.scala 59:18 134:49 27:26]
  wire  _GEN_1998 = 3'h4 == state ? 1'h0 : valid_1_0; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_1999 = 3'h4 == state ? 1'h0 : valid_1_1; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2000 = 3'h4 == state ? 1'h0 : valid_1_2; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2001 = 3'h4 == state ? 1'h0 : valid_1_3; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2002 = 3'h4 == state ? 1'h0 : valid_1_4; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2003 = 3'h4 == state ? 1'h0 : valid_1_5; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2004 = 3'h4 == state ? 1'h0 : valid_1_6; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2005 = 3'h4 == state ? 1'h0 : valid_1_7; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2006 = 3'h4 == state ? 1'h0 : valid_1_8; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2007 = 3'h4 == state ? 1'h0 : valid_1_9; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2008 = 3'h4 == state ? 1'h0 : valid_1_10; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2009 = 3'h4 == state ? 1'h0 : valid_1_11; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2010 = 3'h4 == state ? 1'h0 : valid_1_12; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2011 = 3'h4 == state ? 1'h0 : valid_1_13; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2012 = 3'h4 == state ? 1'h0 : valid_1_14; // @[i_cache.scala 59:18 135:49 28:26]
  wire  _GEN_2013 = 3'h4 == state ? 1'h0 : valid_1_15; // @[i_cache.scala 59:18 135:49 28:26]
  wire [2:0] _GEN_2014 = 3'h4 == state ? 3'h0 : state; // @[i_cache.scala 136:18 59:18 56:24]
  wire [2:0] _GEN_2015 = 3'h3 == state ? 3'h1 : _GEN_2014; // @[i_cache.scala 59:18 88:19]
  wire [127:0] _GEN_2016 = 3'h3 == state ? _GEN_1774 : ram_0_0; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2017 = 3'h3 == state ? _GEN_1775 : ram_0_1; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2018 = 3'h3 == state ? _GEN_1776 : ram_0_2; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2019 = 3'h3 == state ? _GEN_1777 : ram_0_3; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2020 = 3'h3 == state ? _GEN_1778 : ram_0_4; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2021 = 3'h3 == state ? _GEN_1779 : ram_0_5; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2022 = 3'h3 == state ? _GEN_1780 : ram_0_6; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2023 = 3'h3 == state ? _GEN_1781 : ram_0_7; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2024 = 3'h3 == state ? _GEN_1782 : ram_0_8; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2025 = 3'h3 == state ? _GEN_1783 : ram_0_9; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2026 = 3'h3 == state ? _GEN_1784 : ram_0_10; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2027 = 3'h3 == state ? _GEN_1785 : ram_0_11; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2028 = 3'h3 == state ? _GEN_1786 : ram_0_12; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2029 = 3'h3 == state ? _GEN_1787 : ram_0_13; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2030 = 3'h3 == state ? _GEN_1788 : ram_0_14; // @[i_cache.scala 59:18 19:24]
  wire [127:0] _GEN_2031 = 3'h3 == state ? _GEN_1789 : ram_0_15; // @[i_cache.scala 59:18 19:24]
  wire [31:0] _GEN_2032 = 3'h3 == state ? _GEN_1790 : tag_0_0; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2033 = 3'h3 == state ? _GEN_1791 : tag_0_1; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2034 = 3'h3 == state ? _GEN_1792 : tag_0_2; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2035 = 3'h3 == state ? _GEN_1793 : tag_0_3; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2036 = 3'h3 == state ? _GEN_1794 : tag_0_4; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2037 = 3'h3 == state ? _GEN_1795 : tag_0_5; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2038 = 3'h3 == state ? _GEN_1796 : tag_0_6; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2039 = 3'h3 == state ? _GEN_1797 : tag_0_7; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2040 = 3'h3 == state ? _GEN_1798 : tag_0_8; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2041 = 3'h3 == state ? _GEN_1799 : tag_0_9; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2042 = 3'h3 == state ? _GEN_1800 : tag_0_10; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2043 = 3'h3 == state ? _GEN_1801 : tag_0_11; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2044 = 3'h3 == state ? _GEN_1802 : tag_0_12; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2045 = 3'h3 == state ? _GEN_1803 : tag_0_13; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2046 = 3'h3 == state ? _GEN_1804 : tag_0_14; // @[i_cache.scala 59:18 23:24]
  wire [31:0] _GEN_2047 = 3'h3 == state ? _GEN_1805 : tag_0_15; // @[i_cache.scala 59:18 23:24]
  wire  _GEN_2048 = 3'h3 == state ? _GEN_1806 : _GEN_1982; // @[i_cache.scala 59:18]
  wire  _GEN_2049 = 3'h3 == state ? _GEN_1807 : _GEN_1983; // @[i_cache.scala 59:18]
  wire  _GEN_2050 = 3'h3 == state ? _GEN_1808 : _GEN_1984; // @[i_cache.scala 59:18]
  wire  _GEN_2051 = 3'h3 == state ? _GEN_1809 : _GEN_1985; // @[i_cache.scala 59:18]
  wire  _GEN_2052 = 3'h3 == state ? _GEN_1810 : _GEN_1986; // @[i_cache.scala 59:18]
  wire  _GEN_2053 = 3'h3 == state ? _GEN_1811 : _GEN_1987; // @[i_cache.scala 59:18]
  wire  _GEN_2054 = 3'h3 == state ? _GEN_1812 : _GEN_1988; // @[i_cache.scala 59:18]
  wire  _GEN_2055 = 3'h3 == state ? _GEN_1813 : _GEN_1989; // @[i_cache.scala 59:18]
  wire  _GEN_2056 = 3'h3 == state ? _GEN_1814 : _GEN_1990; // @[i_cache.scala 59:18]
  wire  _GEN_2057 = 3'h3 == state ? _GEN_1815 : _GEN_1991; // @[i_cache.scala 59:18]
  wire  _GEN_2058 = 3'h3 == state ? _GEN_1816 : _GEN_1992; // @[i_cache.scala 59:18]
  wire  _GEN_2059 = 3'h3 == state ? _GEN_1817 : _GEN_1993; // @[i_cache.scala 59:18]
  wire  _GEN_2060 = 3'h3 == state ? _GEN_1818 : _GEN_1994; // @[i_cache.scala 59:18]
  wire  _GEN_2061 = 3'h3 == state ? _GEN_1819 : _GEN_1995; // @[i_cache.scala 59:18]
  wire  _GEN_2062 = 3'h3 == state ? _GEN_1820 : _GEN_1996; // @[i_cache.scala 59:18]
  wire  _GEN_2063 = 3'h3 == state ? _GEN_1821 : _GEN_1997; // @[i_cache.scala 59:18]
  wire [7:0] _GEN_2064 = 3'h3 == state ? _GEN_1822 : quene_0; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2065 = 3'h3 == state ? _GEN_1823 : quene_1; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2066 = 3'h3 == state ? _GEN_1824 : quene_2; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2067 = 3'h3 == state ? _GEN_1825 : quene_3; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2068 = 3'h3 == state ? _GEN_1826 : quene_4; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2069 = 3'h3 == state ? _GEN_1827 : quene_5; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2070 = 3'h3 == state ? _GEN_1828 : quene_6; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2071 = 3'h3 == state ? _GEN_1829 : quene_7; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2072 = 3'h3 == state ? _GEN_1830 : quene_8; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2073 = 3'h3 == state ? _GEN_1831 : quene_9; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2074 = 3'h3 == state ? _GEN_1832 : quene_10; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2075 = 3'h3 == state ? _GEN_1833 : quene_11; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2076 = 3'h3 == state ? _GEN_1834 : quene_12; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2077 = 3'h3 == state ? _GEN_1835 : quene_13; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2078 = 3'h3 == state ? _GEN_1836 : quene_14; // @[i_cache.scala 59:18 42:24]
  wire [7:0] _GEN_2079 = 3'h3 == state ? _GEN_1837 : quene_15; // @[i_cache.scala 59:18 42:24]
  wire [127:0] _GEN_2080 = 3'h3 == state ? _GEN_1838 : ram_1_0; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2081 = 3'h3 == state ? _GEN_1839 : ram_1_1; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2082 = 3'h3 == state ? _GEN_1840 : ram_1_2; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2083 = 3'h3 == state ? _GEN_1841 : ram_1_3; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2084 = 3'h3 == state ? _GEN_1842 : ram_1_4; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2085 = 3'h3 == state ? _GEN_1843 : ram_1_5; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2086 = 3'h3 == state ? _GEN_1844 : ram_1_6; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2087 = 3'h3 == state ? _GEN_1845 : ram_1_7; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2088 = 3'h3 == state ? _GEN_1846 : ram_1_8; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2089 = 3'h3 == state ? _GEN_1847 : ram_1_9; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2090 = 3'h3 == state ? _GEN_1848 : ram_1_10; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2091 = 3'h3 == state ? _GEN_1849 : ram_1_11; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2092 = 3'h3 == state ? _GEN_1850 : ram_1_12; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2093 = 3'h3 == state ? _GEN_1851 : ram_1_13; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2094 = 3'h3 == state ? _GEN_1852 : ram_1_14; // @[i_cache.scala 59:18 20:24]
  wire [127:0] _GEN_2095 = 3'h3 == state ? _GEN_1853 : ram_1_15; // @[i_cache.scala 59:18 20:24]
  wire [31:0] _GEN_2096 = 3'h3 == state ? _GEN_1854 : tag_1_0; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2097 = 3'h3 == state ? _GEN_1855 : tag_1_1; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2098 = 3'h3 == state ? _GEN_1856 : tag_1_2; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2099 = 3'h3 == state ? _GEN_1857 : tag_1_3; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2100 = 3'h3 == state ? _GEN_1858 : tag_1_4; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2101 = 3'h3 == state ? _GEN_1859 : tag_1_5; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2102 = 3'h3 == state ? _GEN_1860 : tag_1_6; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2103 = 3'h3 == state ? _GEN_1861 : tag_1_7; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2104 = 3'h3 == state ? _GEN_1862 : tag_1_8; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2105 = 3'h3 == state ? _GEN_1863 : tag_1_9; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2106 = 3'h3 == state ? _GEN_1864 : tag_1_10; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2107 = 3'h3 == state ? _GEN_1865 : tag_1_11; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2108 = 3'h3 == state ? _GEN_1866 : tag_1_12; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2109 = 3'h3 == state ? _GEN_1867 : tag_1_13; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2110 = 3'h3 == state ? _GEN_1868 : tag_1_14; // @[i_cache.scala 59:18 24:24]
  wire [31:0] _GEN_2111 = 3'h3 == state ? _GEN_1869 : tag_1_15; // @[i_cache.scala 59:18 24:24]
  wire  _GEN_2112 = 3'h3 == state ? _GEN_1870 : _GEN_1998; // @[i_cache.scala 59:18]
  wire  _GEN_2113 = 3'h3 == state ? _GEN_1871 : _GEN_1999; // @[i_cache.scala 59:18]
  wire  _GEN_2114 = 3'h3 == state ? _GEN_1872 : _GEN_2000; // @[i_cache.scala 59:18]
  wire  _GEN_2115 = 3'h3 == state ? _GEN_1873 : _GEN_2001; // @[i_cache.scala 59:18]
  wire  _GEN_2116 = 3'h3 == state ? _GEN_1874 : _GEN_2002; // @[i_cache.scala 59:18]
  wire  _GEN_2117 = 3'h3 == state ? _GEN_1875 : _GEN_2003; // @[i_cache.scala 59:18]
  wire  _GEN_2118 = 3'h3 == state ? _GEN_1876 : _GEN_2004; // @[i_cache.scala 59:18]
  wire  _GEN_2119 = 3'h3 == state ? _GEN_1877 : _GEN_2005; // @[i_cache.scala 59:18]
  wire  _GEN_2120 = 3'h3 == state ? _GEN_1878 : _GEN_2006; // @[i_cache.scala 59:18]
  wire  _GEN_2121 = 3'h3 == state ? _GEN_1879 : _GEN_2007; // @[i_cache.scala 59:18]
  wire  _GEN_2122 = 3'h3 == state ? _GEN_1880 : _GEN_2008; // @[i_cache.scala 59:18]
  wire  _GEN_2123 = 3'h3 == state ? _GEN_1881 : _GEN_2009; // @[i_cache.scala 59:18]
  wire  _GEN_2124 = 3'h3 == state ? _GEN_1882 : _GEN_2010; // @[i_cache.scala 59:18]
  wire  _GEN_2125 = 3'h3 == state ? _GEN_1883 : _GEN_2011; // @[i_cache.scala 59:18]
  wire  _GEN_2126 = 3'h3 == state ? _GEN_1884 : _GEN_2012; // @[i_cache.scala 59:18]
  wire  _GEN_2127 = 3'h3 == state ? _GEN_1885 : _GEN_2013; // @[i_cache.scala 59:18]
  wire [127:0] _GEN_2128 = 3'h3 == state ? _GEN_1886 : ram_2_0; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2129 = 3'h3 == state ? _GEN_1887 : ram_2_1; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2130 = 3'h3 == state ? _GEN_1888 : ram_2_2; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2131 = 3'h3 == state ? _GEN_1889 : ram_2_3; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2132 = 3'h3 == state ? _GEN_1890 : ram_2_4; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2133 = 3'h3 == state ? _GEN_1891 : ram_2_5; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2134 = 3'h3 == state ? _GEN_1892 : ram_2_6; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2135 = 3'h3 == state ? _GEN_1893 : ram_2_7; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2136 = 3'h3 == state ? _GEN_1894 : ram_2_8; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2137 = 3'h3 == state ? _GEN_1895 : ram_2_9; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2138 = 3'h3 == state ? _GEN_1896 : ram_2_10; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2139 = 3'h3 == state ? _GEN_1897 : ram_2_11; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2140 = 3'h3 == state ? _GEN_1898 : ram_2_12; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2141 = 3'h3 == state ? _GEN_1899 : ram_2_13; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2142 = 3'h3 == state ? _GEN_1900 : ram_2_14; // @[i_cache.scala 59:18 21:24]
  wire [127:0] _GEN_2143 = 3'h3 == state ? _GEN_1901 : ram_2_15; // @[i_cache.scala 59:18 21:24]
  wire [31:0] _GEN_2144 = 3'h3 == state ? _GEN_1902 : tag_2_0; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2145 = 3'h3 == state ? _GEN_1903 : tag_2_1; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2146 = 3'h3 == state ? _GEN_1904 : tag_2_2; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2147 = 3'h3 == state ? _GEN_1905 : tag_2_3; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2148 = 3'h3 == state ? _GEN_1906 : tag_2_4; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2149 = 3'h3 == state ? _GEN_1907 : tag_2_5; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2150 = 3'h3 == state ? _GEN_1908 : tag_2_6; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2151 = 3'h3 == state ? _GEN_1909 : tag_2_7; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2152 = 3'h3 == state ? _GEN_1910 : tag_2_8; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2153 = 3'h3 == state ? _GEN_1911 : tag_2_9; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2154 = 3'h3 == state ? _GEN_1912 : tag_2_10; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2155 = 3'h3 == state ? _GEN_1913 : tag_2_11; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2156 = 3'h3 == state ? _GEN_1914 : tag_2_12; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2157 = 3'h3 == state ? _GEN_1915 : tag_2_13; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2158 = 3'h3 == state ? _GEN_1916 : tag_2_14; // @[i_cache.scala 59:18 25:24]
  wire [31:0] _GEN_2159 = 3'h3 == state ? _GEN_1917 : tag_2_15; // @[i_cache.scala 59:18 25:24]
  wire  _GEN_2160 = 3'h3 == state ? _GEN_1918 : valid_2_0; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2161 = 3'h3 == state ? _GEN_1919 : valid_2_1; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2162 = 3'h3 == state ? _GEN_1920 : valid_2_2; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2163 = 3'h3 == state ? _GEN_1921 : valid_2_3; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2164 = 3'h3 == state ? _GEN_1922 : valid_2_4; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2165 = 3'h3 == state ? _GEN_1923 : valid_2_5; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2166 = 3'h3 == state ? _GEN_1924 : valid_2_6; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2167 = 3'h3 == state ? _GEN_1925 : valid_2_7; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2168 = 3'h3 == state ? _GEN_1926 : valid_2_8; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2169 = 3'h3 == state ? _GEN_1927 : valid_2_9; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2170 = 3'h3 == state ? _GEN_1928 : valid_2_10; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2171 = 3'h3 == state ? _GEN_1929 : valid_2_11; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2172 = 3'h3 == state ? _GEN_1930 : valid_2_12; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2173 = 3'h3 == state ? _GEN_1931 : valid_2_13; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2174 = 3'h3 == state ? _GEN_1932 : valid_2_14; // @[i_cache.scala 59:18 29:26]
  wire  _GEN_2175 = 3'h3 == state ? _GEN_1933 : valid_2_15; // @[i_cache.scala 59:18 29:26]
  wire [127:0] _GEN_2176 = 3'h3 == state ? _GEN_1934 : ram_3_0; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2177 = 3'h3 == state ? _GEN_1935 : ram_3_1; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2178 = 3'h3 == state ? _GEN_1936 : ram_3_2; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2179 = 3'h3 == state ? _GEN_1937 : ram_3_3; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2180 = 3'h3 == state ? _GEN_1938 : ram_3_4; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2181 = 3'h3 == state ? _GEN_1939 : ram_3_5; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2182 = 3'h3 == state ? _GEN_1940 : ram_3_6; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2183 = 3'h3 == state ? _GEN_1941 : ram_3_7; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2184 = 3'h3 == state ? _GEN_1942 : ram_3_8; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2185 = 3'h3 == state ? _GEN_1943 : ram_3_9; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2186 = 3'h3 == state ? _GEN_1944 : ram_3_10; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2187 = 3'h3 == state ? _GEN_1945 : ram_3_11; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2188 = 3'h3 == state ? _GEN_1946 : ram_3_12; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2189 = 3'h3 == state ? _GEN_1947 : ram_3_13; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2190 = 3'h3 == state ? _GEN_1948 : ram_3_14; // @[i_cache.scala 59:18 22:24]
  wire [127:0] _GEN_2191 = 3'h3 == state ? _GEN_1949 : ram_3_15; // @[i_cache.scala 59:18 22:24]
  wire [31:0] _GEN_2192 = 3'h3 == state ? _GEN_1950 : tag_3_0; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2193 = 3'h3 == state ? _GEN_1951 : tag_3_1; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2194 = 3'h3 == state ? _GEN_1952 : tag_3_2; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2195 = 3'h3 == state ? _GEN_1953 : tag_3_3; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2196 = 3'h3 == state ? _GEN_1954 : tag_3_4; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2197 = 3'h3 == state ? _GEN_1955 : tag_3_5; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2198 = 3'h3 == state ? _GEN_1956 : tag_3_6; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2199 = 3'h3 == state ? _GEN_1957 : tag_3_7; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2200 = 3'h3 == state ? _GEN_1958 : tag_3_8; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2201 = 3'h3 == state ? _GEN_1959 : tag_3_9; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2202 = 3'h3 == state ? _GEN_1960 : tag_3_10; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2203 = 3'h3 == state ? _GEN_1961 : tag_3_11; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2204 = 3'h3 == state ? _GEN_1962 : tag_3_12; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2205 = 3'h3 == state ? _GEN_1963 : tag_3_13; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2206 = 3'h3 == state ? _GEN_1964 : tag_3_14; // @[i_cache.scala 59:18 26:24]
  wire [31:0] _GEN_2207 = 3'h3 == state ? _GEN_1965 : tag_3_15; // @[i_cache.scala 59:18 26:24]
  wire  _GEN_2208 = 3'h3 == state ? _GEN_1966 : valid_3_0; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2209 = 3'h3 == state ? _GEN_1967 : valid_3_1; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2210 = 3'h3 == state ? _GEN_1968 : valid_3_2; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2211 = 3'h3 == state ? _GEN_1969 : valid_3_3; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2212 = 3'h3 == state ? _GEN_1970 : valid_3_4; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2213 = 3'h3 == state ? _GEN_1971 : valid_3_5; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2214 = 3'h3 == state ? _GEN_1972 : valid_3_6; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2215 = 3'h3 == state ? _GEN_1973 : valid_3_7; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2216 = 3'h3 == state ? _GEN_1974 : valid_3_8; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2217 = 3'h3 == state ? _GEN_1975 : valid_3_9; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2218 = 3'h3 == state ? _GEN_1976 : valid_3_10; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2219 = 3'h3 == state ? _GEN_1977 : valid_3_11; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2220 = 3'h3 == state ? _GEN_1978 : valid_3_12; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2221 = 3'h3 == state ? _GEN_1979 : valid_3_13; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2222 = 3'h3 == state ? _GEN_1980 : valid_3_14; // @[i_cache.scala 59:18 30:26]
  wire  _GEN_2223 = 3'h3 == state ? _GEN_1981 : valid_3_15; // @[i_cache.scala 59:18 30:26]
  wire [127:0] _GEN_2862 = 4'h1 == index ? ram_0_1 : ram_0_0; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2863 = 4'h2 == index ? ram_0_2 : _GEN_2862; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2864 = 4'h3 == index ? ram_0_3 : _GEN_2863; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2865 = 4'h4 == index ? ram_0_4 : _GEN_2864; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2866 = 4'h5 == index ? ram_0_5 : _GEN_2865; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2867 = 4'h6 == index ? ram_0_6 : _GEN_2866; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2868 = 4'h7 == index ? ram_0_7 : _GEN_2867; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2869 = 4'h8 == index ? ram_0_8 : _GEN_2868; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2870 = 4'h9 == index ? ram_0_9 : _GEN_2869; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2871 = 4'ha == index ? ram_0_10 : _GEN_2870; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2872 = 4'hb == index ? ram_0_11 : _GEN_2871; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2873 = 4'hc == index ? ram_0_12 : _GEN_2872; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2874 = 4'hd == index ? ram_0_13 : _GEN_2873; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2875 = 4'he == index ? ram_0_14 : _GEN_2874; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _GEN_2876 = 4'hf == index ? ram_0_15 : _GEN_2875; // @[i_cache.scala 157:{55,55}]
  wire [127:0] _io_to_ifu_rdata_T = _GEN_2876 >> shift_bit; // @[i_cache.scala 157:55]
  wire [127:0] _GEN_2878 = 4'h1 == index ? ram_1_1 : ram_1_0; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2879 = 4'h2 == index ? ram_1_2 : _GEN_2878; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2880 = 4'h3 == index ? ram_1_3 : _GEN_2879; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2881 = 4'h4 == index ? ram_1_4 : _GEN_2880; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2882 = 4'h5 == index ? ram_1_5 : _GEN_2881; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2883 = 4'h6 == index ? ram_1_6 : _GEN_2882; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2884 = 4'h7 == index ? ram_1_7 : _GEN_2883; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2885 = 4'h8 == index ? ram_1_8 : _GEN_2884; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2886 = 4'h9 == index ? ram_1_9 : _GEN_2885; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2887 = 4'ha == index ? ram_1_10 : _GEN_2886; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2888 = 4'hb == index ? ram_1_11 : _GEN_2887; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2889 = 4'hc == index ? ram_1_12 : _GEN_2888; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2890 = 4'hd == index ? ram_1_13 : _GEN_2889; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2891 = 4'he == index ? ram_1_14 : _GEN_2890; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _GEN_2892 = 4'hf == index ? ram_1_15 : _GEN_2891; // @[i_cache.scala 157:{95,95}]
  wire [127:0] _io_to_ifu_rdata_T_1 = _GEN_2892 >> shift_bit; // @[i_cache.scala 157:95]
  wire [127:0] _GEN_2894 = 4'h1 == index ? ram_2_1 : ram_2_0; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2895 = 4'h2 == index ? ram_2_2 : _GEN_2894; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2896 = 4'h3 == index ? ram_2_3 : _GEN_2895; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2897 = 4'h4 == index ? ram_2_4 : _GEN_2896; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2898 = 4'h5 == index ? ram_2_5 : _GEN_2897; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2899 = 4'h6 == index ? ram_2_6 : _GEN_2898; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2900 = 4'h7 == index ? ram_2_7 : _GEN_2899; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2901 = 4'h8 == index ? ram_2_8 : _GEN_2900; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2902 = 4'h9 == index ? ram_2_9 : _GEN_2901; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2903 = 4'ha == index ? ram_2_10 : _GEN_2902; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2904 = 4'hb == index ? ram_2_11 : _GEN_2903; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2905 = 4'hc == index ? ram_2_12 : _GEN_2904; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2906 = 4'hd == index ? ram_2_13 : _GEN_2905; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2907 = 4'he == index ? ram_2_14 : _GEN_2906; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _GEN_2908 = 4'hf == index ? ram_2_15 : _GEN_2907; // @[i_cache.scala 157:{135,135}]
  wire [127:0] _io_to_ifu_rdata_T_2 = _GEN_2908 >> shift_bit; // @[i_cache.scala 157:135]
  wire [127:0] _GEN_2910 = 4'h1 == index ? ram_3_1 : ram_3_0; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2911 = 4'h2 == index ? ram_3_2 : _GEN_2910; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2912 = 4'h3 == index ? ram_3_3 : _GEN_2911; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2913 = 4'h4 == index ? ram_3_4 : _GEN_2912; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2914 = 4'h5 == index ? ram_3_5 : _GEN_2913; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2915 = 4'h6 == index ? ram_3_6 : _GEN_2914; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2916 = 4'h7 == index ? ram_3_7 : _GEN_2915; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2917 = 4'h8 == index ? ram_3_8 : _GEN_2916; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2918 = 4'h9 == index ? ram_3_9 : _GEN_2917; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2919 = 4'ha == index ? ram_3_10 : _GEN_2918; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2920 = 4'hb == index ? ram_3_11 : _GEN_2919; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2921 = 4'hc == index ? ram_3_12 : _GEN_2920; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2922 = 4'hd == index ? ram_3_13 : _GEN_2921; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2923 = 4'he == index ? ram_3_14 : _GEN_2922; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _GEN_2924 = 4'hf == index ? ram_3_15 : _GEN_2923; // @[i_cache.scala 157:{162,162}]
  wire [127:0] _io_to_ifu_rdata_T_3 = _GEN_2924 >> shift_bit; // @[i_cache.scala 157:162]
  wire [127:0] _io_to_ifu_rdata_T_4 = way2_hit ? _io_to_ifu_rdata_T_2 : _io_to_ifu_rdata_T_3; // @[i_cache.scala 157:112]
  wire [127:0] _io_to_ifu_rdata_T_5 = way1_hit ? _io_to_ifu_rdata_T_1 : _io_to_ifu_rdata_T_4; // @[i_cache.scala 157:72]
  wire [127:0] _io_to_ifu_rdata_T_6 = way0_hit ? _io_to_ifu_rdata_T : _io_to_ifu_rdata_T_5; // @[i_cache.scala 157:32]
  wire  _T_20 = state == 3'h2; // @[i_cache.scala 164:21]
  wire [63:0] _GEN_3077 = {{32'd0}, addr}; // @[i_cache.scala 173:35]
  wire [63:0] _io_to_axi_araddr_T = _GEN_3077 & 64'hfffffffffffffff0; // @[i_cache.scala 173:35]
  wire  _GEN_2926 = state == 3'h2 ? 1'h0 : state == 3'h0; // @[i_cache.scala 164:29 166:27 190:27]
  wire [63:0] _GEN_2928 = state == 3'h2 ? _io_to_axi_araddr_T : {{32'd0}, addr}; // @[i_cache.scala 164:29 173:26 197:26]
  wire  _GEN_2930 = state == 3'h2 | io_from_ifu_rready; // @[i_cache.scala 164:29 177:26 198:26]
  wire  _GEN_2931 = state == 3'h1 ? 1'h0 : _T_20; // @[i_cache.scala 140:25 141:27]
  wire [63:0] _GEN_2932 = state == 3'h1 ? {{32'd0}, addr} : _GEN_2928; // @[i_cache.scala 140:25 142:26]
  wire [127:0] _GEN_2936 = state == 3'h1 ? _io_to_ifu_rdata_T_6 : 128'h0; // @[i_cache.scala 140:25 157:25]
  assign io_to_ifu_arready = state == 3'h1 ? 1'h0 : _GEN_2926; // @[i_cache.scala 140:25 158:27]
  assign io_to_ifu_rdata = _GEN_2936[63:0];
  assign io_to_ifu_rvalid = state == 3'h1 & _T_4; // @[i_cache.scala 140:25 159:26]
  assign io_to_axi_araddr = _GEN_2932[31:0];
  assign io_to_axi_arlen = {{7'd0}, _GEN_2931};
  assign io_to_axi_arvalid = state == 3'h1 ? 1'h0 : _T_20; // @[i_cache.scala 140:25 141:27]
  assign io_to_axi_rready = state == 3'h1 ? 1'h0 : _GEN_2930; // @[i_cache.scala 140:25 146:26]
  assign io_cache_init = state == 3'h4; // @[i_cache.scala 213:27]
  always @(posedge clock) begin
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_0 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_0 <= _GEN_2016;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_1 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_1 <= _GEN_2017;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_2 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_2 <= _GEN_2018;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_3 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_3 <= _GEN_2019;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_4 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_4 <= _GEN_2020;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_5 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_5 <= _GEN_2021;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_6 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_6 <= _GEN_2022;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_7 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_7 <= _GEN_2023;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_8 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_8 <= _GEN_2024;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_9 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_9 <= _GEN_2025;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_10 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_10 <= _GEN_2026;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_11 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_11 <= _GEN_2027;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_12 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_12 <= _GEN_2028;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_13 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_13 <= _GEN_2029;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_14 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_14 <= _GEN_2030;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 19:24]
      ram_0_15 <= 128'h0; // @[i_cache.scala 19:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_0_15 <= _GEN_2031;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_0 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_0 <= _GEN_2080;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_1 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_1 <= _GEN_2081;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_2 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_2 <= _GEN_2082;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_3 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_3 <= _GEN_2083;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_4 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_4 <= _GEN_2084;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_5 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_5 <= _GEN_2085;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_6 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_6 <= _GEN_2086;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_7 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_7 <= _GEN_2087;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_8 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_8 <= _GEN_2088;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_9 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_9 <= _GEN_2089;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_10 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_10 <= _GEN_2090;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_11 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_11 <= _GEN_2091;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_12 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_12 <= _GEN_2092;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_13 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_13 <= _GEN_2093;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_14 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_14 <= _GEN_2094;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 20:24]
      ram_1_15 <= 128'h0; // @[i_cache.scala 20:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_1_15 <= _GEN_2095;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_0 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_0 <= _GEN_2128;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_1 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_1 <= _GEN_2129;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_2 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_2 <= _GEN_2130;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_3 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_3 <= _GEN_2131;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_4 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_4 <= _GEN_2132;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_5 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_5 <= _GEN_2133;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_6 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_6 <= _GEN_2134;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_7 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_7 <= _GEN_2135;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_8 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_8 <= _GEN_2136;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_9 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_9 <= _GEN_2137;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_10 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_10 <= _GEN_2138;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_11 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_11 <= _GEN_2139;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_12 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_12 <= _GEN_2140;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_13 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_13 <= _GEN_2141;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_14 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_14 <= _GEN_2142;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 21:24]
      ram_2_15 <= 128'h0; // @[i_cache.scala 21:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_2_15 <= _GEN_2143;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_0 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_0 <= _GEN_2176;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_1 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_1 <= _GEN_2177;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_2 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_2 <= _GEN_2178;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_3 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_3 <= _GEN_2179;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_4 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_4 <= _GEN_2180;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_5 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_5 <= _GEN_2181;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_6 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_6 <= _GEN_2182;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_7 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_7 <= _GEN_2183;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_8 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_8 <= _GEN_2184;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_9 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_9 <= _GEN_2185;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_10 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_10 <= _GEN_2186;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_11 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_11 <= _GEN_2187;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_12 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_12 <= _GEN_2188;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_13 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_13 <= _GEN_2189;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_14 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_14 <= _GEN_2190;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 22:24]
      ram_3_15 <= 128'h0; // @[i_cache.scala 22:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          ram_3_15 <= _GEN_2191;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_0 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_0 <= _GEN_2032;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_1 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_1 <= _GEN_2033;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_2 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_2 <= _GEN_2034;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_3 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_3 <= _GEN_2035;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_4 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_4 <= _GEN_2036;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_5 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_5 <= _GEN_2037;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_6 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_6 <= _GEN_2038;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_7 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_7 <= _GEN_2039;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_8 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_8 <= _GEN_2040;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_9 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_9 <= _GEN_2041;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_10 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_10 <= _GEN_2042;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_11 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_11 <= _GEN_2043;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_12 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_12 <= _GEN_2044;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_13 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_13 <= _GEN_2045;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_14 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_14 <= _GEN_2046;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 23:24]
      tag_0_15 <= 32'h0; // @[i_cache.scala 23:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_0_15 <= _GEN_2047;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_0 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_0 <= _GEN_2096;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_1 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_1 <= _GEN_2097;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_2 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_2 <= _GEN_2098;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_3 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_3 <= _GEN_2099;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_4 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_4 <= _GEN_2100;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_5 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_5 <= _GEN_2101;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_6 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_6 <= _GEN_2102;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_7 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_7 <= _GEN_2103;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_8 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_8 <= _GEN_2104;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_9 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_9 <= _GEN_2105;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_10 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_10 <= _GEN_2106;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_11 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_11 <= _GEN_2107;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_12 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_12 <= _GEN_2108;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_13 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_13 <= _GEN_2109;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_14 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_14 <= _GEN_2110;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 24:24]
      tag_1_15 <= 32'h0; // @[i_cache.scala 24:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_1_15 <= _GEN_2111;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_0 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_0 <= _GEN_2144;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_1 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_1 <= _GEN_2145;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_2 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_2 <= _GEN_2146;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_3 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_3 <= _GEN_2147;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_4 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_4 <= _GEN_2148;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_5 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_5 <= _GEN_2149;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_6 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_6 <= _GEN_2150;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_7 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_7 <= _GEN_2151;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_8 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_8 <= _GEN_2152;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_9 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_9 <= _GEN_2153;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_10 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_10 <= _GEN_2154;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_11 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_11 <= _GEN_2155;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_12 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_12 <= _GEN_2156;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_13 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_13 <= _GEN_2157;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_14 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_14 <= _GEN_2158;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 25:24]
      tag_2_15 <= 32'h0; // @[i_cache.scala 25:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_2_15 <= _GEN_2159;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_0 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_0 <= _GEN_2192;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_1 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_1 <= _GEN_2193;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_2 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_2 <= _GEN_2194;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_3 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_3 <= _GEN_2195;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_4 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_4 <= _GEN_2196;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_5 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_5 <= _GEN_2197;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_6 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_6 <= _GEN_2198;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_7 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_7 <= _GEN_2199;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_8 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_8 <= _GEN_2200;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_9 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_9 <= _GEN_2201;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_10 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_10 <= _GEN_2202;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_11 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_11 <= _GEN_2203;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_12 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_12 <= _GEN_2204;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_13 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_13 <= _GEN_2205;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_14 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_14 <= _GEN_2206;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 26:24]
      tag_3_15 <= 32'h0; // @[i_cache.scala 26:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          tag_3_15 <= _GEN_2207;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_0 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_0 <= _GEN_2048;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_1 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_1 <= _GEN_2049;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_2 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_2 <= _GEN_2050;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_3 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_3 <= _GEN_2051;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_4 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_4 <= _GEN_2052;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_5 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_5 <= _GEN_2053;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_6 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_6 <= _GEN_2054;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_7 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_7 <= _GEN_2055;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_8 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_8 <= _GEN_2056;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_9 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_9 <= _GEN_2057;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_10 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_10 <= _GEN_2058;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_11 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_11 <= _GEN_2059;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_12 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_12 <= _GEN_2060;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_13 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_13 <= _GEN_2061;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_14 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_14 <= _GEN_2062;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 27:26]
      valid_0_15 <= 1'h0; // @[i_cache.scala 27:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_0_15 <= _GEN_2063;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_0 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_0 <= _GEN_2112;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_1 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_1 <= _GEN_2113;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_2 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_2 <= _GEN_2114;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_3 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_3 <= _GEN_2115;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_4 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_4 <= _GEN_2116;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_5 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_5 <= _GEN_2117;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_6 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_6 <= _GEN_2118;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_7 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_7 <= _GEN_2119;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_8 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_8 <= _GEN_2120;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_9 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_9 <= _GEN_2121;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_10 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_10 <= _GEN_2122;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_11 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_11 <= _GEN_2123;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_12 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_12 <= _GEN_2124;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_13 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_13 <= _GEN_2125;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_14 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_14 <= _GEN_2126;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 28:26]
      valid_1_15 <= 1'h0; // @[i_cache.scala 28:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_1_15 <= _GEN_2127;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_0 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_0 <= _GEN_2160;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_1 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_1 <= _GEN_2161;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_2 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_2 <= _GEN_2162;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_3 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_3 <= _GEN_2163;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_4 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_4 <= _GEN_2164;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_5 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_5 <= _GEN_2165;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_6 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_6 <= _GEN_2166;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_7 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_7 <= _GEN_2167;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_8 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_8 <= _GEN_2168;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_9 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_9 <= _GEN_2169;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_10 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_10 <= _GEN_2170;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_11 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_11 <= _GEN_2171;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_12 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_12 <= _GEN_2172;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_13 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_13 <= _GEN_2173;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_14 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_14 <= _GEN_2174;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 29:26]
      valid_2_15 <= 1'h0; // @[i_cache.scala 29:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_2_15 <= _GEN_2175;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_0 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_0 <= _GEN_2208;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_1 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_1 <= _GEN_2209;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_2 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_2 <= _GEN_2210;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_3 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_3 <= _GEN_2211;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_4 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_4 <= _GEN_2212;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_5 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_5 <= _GEN_2213;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_6 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_6 <= _GEN_2214;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_7 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_7 <= _GEN_2215;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_8 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_8 <= _GEN_2216;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_9 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_9 <= _GEN_2217;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_10 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_10 <= _GEN_2218;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_11 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_11 <= _GEN_2219;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_12 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_12 <= _GEN_2220;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_13 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_13 <= _GEN_2221;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_14 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_14 <= _GEN_2222;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 30:26]
      valid_3_15 <= 1'h0; // @[i_cache.scala 30:26]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          valid_3_15 <= _GEN_2223;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 32:23]
      addr <= 32'h0; // @[i_cache.scala 32:23]
    end else if (3'h0 == state) begin // @[i_cache.scala 59:18]
      if (!(io_clear_cache)) begin // @[i_cache.scala 61:33]
        if (io_from_ifu_arvalid) begin // @[i_cache.scala 63:44]
          addr <= io_from_ifu_araddr; // @[i_cache.scala 64:22]
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:31]
      receive_data_0 <= 64'h0; // @[i_cache.scala 40:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (3'h2 == state) begin // @[i_cache.scala 59:18]
          receive_data_0 <= _GEN_138;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 40:31]
      receive_data_1 <= 64'h0; // @[i_cache.scala 40:31]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (3'h2 == state) begin // @[i_cache.scala 59:18]
          receive_data_1 <= _GEN_139;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 41:30]
      receive_num <= 3'h0; // @[i_cache.scala 41:30]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (3'h1 == state) begin // @[i_cache.scala 59:18]
        if (!(way0_hit | way1_hit | way2_hit | way3_hit)) begin // @[i_cache.scala 69:57]
          receive_num <= 3'h0; // @[i_cache.scala 75:29]
        end
      end else if (3'h2 == state) begin // @[i_cache.scala 59:18]
        receive_num <= _GEN_140;
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_0 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_0 <= _GEN_2064;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_1 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_1 <= _GEN_2065;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_2 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_2 <= _GEN_2066;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_3 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_3 <= _GEN_2067;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_4 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_4 <= _GEN_2068;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_5 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_5 <= _GEN_2069;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_6 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_6 <= _GEN_2070;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_7 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_7 <= _GEN_2071;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_8 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_8 <= _GEN_2072;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_9 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_9 <= _GEN_2073;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_10 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_10 <= _GEN_2074;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_11 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_11 <= _GEN_2075;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_12 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_12 <= _GEN_2076;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_13 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_13 <= _GEN_2077;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_14 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_14 <= _GEN_2078;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 42:24]
      quene_15 <= 8'h0; // @[i_cache.scala 42:24]
    end else if (!(3'h0 == state)) begin // @[i_cache.scala 59:18]
      if (!(3'h1 == state)) begin // @[i_cache.scala 59:18]
        if (!(3'h2 == state)) begin // @[i_cache.scala 59:18]
          quene_15 <= _GEN_2079;
        end
      end
    end
    if (reset) begin // @[i_cache.scala 56:24]
      state <= 3'h0; // @[i_cache.scala 56:24]
    end else if (3'h0 == state) begin // @[i_cache.scala 59:18]
      if (io_clear_cache) begin // @[i_cache.scala 61:33]
        state <= 3'h4; // @[i_cache.scala 62:23]
      end else if (io_from_ifu_arvalid) begin // @[i_cache.scala 63:44]
        state <= 3'h1; // @[i_cache.scala 65:23]
      end
    end else if (3'h1 == state) begin // @[i_cache.scala 59:18]
      if (way0_hit | way1_hit | way2_hit | way3_hit) begin // @[i_cache.scala 69:57]
        state <= _GEN_132;
      end else begin
        state <= 3'h2; // @[i_cache.scala 74:23]
      end
    end else if (3'h2 == state) begin // @[i_cache.scala 59:18]
      state <= _GEN_141;
    end else begin
      state <= _GEN_2015;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  ram_0_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  ram_0_1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  ram_0_2 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  ram_0_3 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  ram_0_4 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  ram_0_5 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  ram_0_6 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  ram_0_7 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  ram_0_8 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  ram_0_9 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  ram_0_10 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  ram_0_11 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  ram_0_12 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  ram_0_13 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  ram_0_14 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  ram_0_15 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  ram_1_0 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  ram_1_1 = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  ram_1_2 = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  ram_1_3 = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  ram_1_4 = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  ram_1_5 = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  ram_1_6 = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  ram_1_7 = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  ram_1_8 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  ram_1_9 = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  ram_1_10 = _RAND_26[127:0];
  _RAND_27 = {4{`RANDOM}};
  ram_1_11 = _RAND_27[127:0];
  _RAND_28 = {4{`RANDOM}};
  ram_1_12 = _RAND_28[127:0];
  _RAND_29 = {4{`RANDOM}};
  ram_1_13 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  ram_1_14 = _RAND_30[127:0];
  _RAND_31 = {4{`RANDOM}};
  ram_1_15 = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  ram_2_0 = _RAND_32[127:0];
  _RAND_33 = {4{`RANDOM}};
  ram_2_1 = _RAND_33[127:0];
  _RAND_34 = {4{`RANDOM}};
  ram_2_2 = _RAND_34[127:0];
  _RAND_35 = {4{`RANDOM}};
  ram_2_3 = _RAND_35[127:0];
  _RAND_36 = {4{`RANDOM}};
  ram_2_4 = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  ram_2_5 = _RAND_37[127:0];
  _RAND_38 = {4{`RANDOM}};
  ram_2_6 = _RAND_38[127:0];
  _RAND_39 = {4{`RANDOM}};
  ram_2_7 = _RAND_39[127:0];
  _RAND_40 = {4{`RANDOM}};
  ram_2_8 = _RAND_40[127:0];
  _RAND_41 = {4{`RANDOM}};
  ram_2_9 = _RAND_41[127:0];
  _RAND_42 = {4{`RANDOM}};
  ram_2_10 = _RAND_42[127:0];
  _RAND_43 = {4{`RANDOM}};
  ram_2_11 = _RAND_43[127:0];
  _RAND_44 = {4{`RANDOM}};
  ram_2_12 = _RAND_44[127:0];
  _RAND_45 = {4{`RANDOM}};
  ram_2_13 = _RAND_45[127:0];
  _RAND_46 = {4{`RANDOM}};
  ram_2_14 = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  ram_2_15 = _RAND_47[127:0];
  _RAND_48 = {4{`RANDOM}};
  ram_3_0 = _RAND_48[127:0];
  _RAND_49 = {4{`RANDOM}};
  ram_3_1 = _RAND_49[127:0];
  _RAND_50 = {4{`RANDOM}};
  ram_3_2 = _RAND_50[127:0];
  _RAND_51 = {4{`RANDOM}};
  ram_3_3 = _RAND_51[127:0];
  _RAND_52 = {4{`RANDOM}};
  ram_3_4 = _RAND_52[127:0];
  _RAND_53 = {4{`RANDOM}};
  ram_3_5 = _RAND_53[127:0];
  _RAND_54 = {4{`RANDOM}};
  ram_3_6 = _RAND_54[127:0];
  _RAND_55 = {4{`RANDOM}};
  ram_3_7 = _RAND_55[127:0];
  _RAND_56 = {4{`RANDOM}};
  ram_3_8 = _RAND_56[127:0];
  _RAND_57 = {4{`RANDOM}};
  ram_3_9 = _RAND_57[127:0];
  _RAND_58 = {4{`RANDOM}};
  ram_3_10 = _RAND_58[127:0];
  _RAND_59 = {4{`RANDOM}};
  ram_3_11 = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  ram_3_12 = _RAND_60[127:0];
  _RAND_61 = {4{`RANDOM}};
  ram_3_13 = _RAND_61[127:0];
  _RAND_62 = {4{`RANDOM}};
  ram_3_14 = _RAND_62[127:0];
  _RAND_63 = {4{`RANDOM}};
  ram_3_15 = _RAND_63[127:0];
  _RAND_64 = {1{`RANDOM}};
  tag_0_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  tag_0_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  tag_0_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  tag_0_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  tag_0_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  tag_0_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  tag_0_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  tag_0_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  tag_0_8 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  tag_0_9 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  tag_0_10 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  tag_0_11 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  tag_0_12 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  tag_0_13 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  tag_0_14 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  tag_0_15 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  tag_1_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  tag_1_1 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  tag_1_2 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  tag_1_3 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  tag_1_4 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  tag_1_5 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  tag_1_6 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  tag_1_7 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  tag_1_8 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  tag_1_9 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  tag_1_10 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  tag_1_11 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  tag_1_12 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  tag_1_13 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  tag_1_14 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  tag_1_15 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  tag_2_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  tag_2_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  tag_2_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  tag_2_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  tag_2_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  tag_2_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  tag_2_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  tag_2_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  tag_2_8 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  tag_2_9 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  tag_2_10 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  tag_2_11 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  tag_2_12 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  tag_2_13 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  tag_2_14 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  tag_2_15 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  tag_3_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  tag_3_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  tag_3_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  tag_3_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  tag_3_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  tag_3_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  tag_3_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  tag_3_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  tag_3_8 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  tag_3_9 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  tag_3_10 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  tag_3_11 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  tag_3_12 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  tag_3_13 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  tag_3_14 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  tag_3_15 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_1_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_1_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_1_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_1_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_1_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_1_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_1_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_1_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_1_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_1_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_1_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_1_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_1_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_1_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_1_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_1_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_2_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_2_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_2_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_2_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_2_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_2_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_2_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_2_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_2_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_2_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_2_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_2_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_2_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_2_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_2_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_2_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_3_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_3_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_3_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_3_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_3_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_3_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_3_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_3_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_3_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_3_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_3_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_3_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_3_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_3_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_3_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_3_15 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  addr = _RAND_192[31:0];
  _RAND_193 = {2{`RANDOM}};
  receive_data_0 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  receive_data_1 = _RAND_194[63:0];
  _RAND_195 = {1{`RANDOM}};
  receive_num = _RAND_195[2:0];
  _RAND_196 = {1{`RANDOM}};
  quene_0 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  quene_1 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  quene_2 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  quene_3 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  quene_4 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  quene_5 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  quene_6 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  quene_7 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  quene_8 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  quene_9 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  quene_10 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  quene_11 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  quene_12 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  quene_13 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  quene_14 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  quene_15 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  state = _RAND_212[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [63:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_bvalid,
  output [31:0] io_to_axi_araddr,
  output [7:0]  io_to_axi_arlen,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output [7:0]  io_to_axi_awlen,
  output        io_to_axi_awvalid,
  output [63:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rlast,
  input         io_from_axi_rvalid,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [127:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] ram_0_0; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_1; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_2; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_3; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_4; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_5; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_6; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_7; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_8; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_9; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_10; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_11; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_12; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_13; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_14; // @[d_cache.scala 19:24]
  reg [127:0] ram_0_15; // @[d_cache.scala 19:24]
  reg [127:0] ram_1_0; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_1; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_2; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_3; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_4; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_5; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_6; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_7; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_8; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_9; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_10; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_11; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_12; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_13; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_14; // @[d_cache.scala 20:24]
  reg [127:0] ram_1_15; // @[d_cache.scala 20:24]
  reg [31:0] tag_0_0; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 22:24]
  reg [31:0] tag_1_0; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_1; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_2; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_3; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_4; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_5; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_6; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_7; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_8; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_9; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_10; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_11; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_12; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_13; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_14; // @[d_cache.scala 23:24]
  reg [31:0] tag_1_15; // @[d_cache.scala 23:24]
  reg  valid_0_0; // @[d_cache.scala 24:26]
  reg  valid_0_1; // @[d_cache.scala 24:26]
  reg  valid_0_2; // @[d_cache.scala 24:26]
  reg  valid_0_3; // @[d_cache.scala 24:26]
  reg  valid_0_4; // @[d_cache.scala 24:26]
  reg  valid_0_5; // @[d_cache.scala 24:26]
  reg  valid_0_6; // @[d_cache.scala 24:26]
  reg  valid_0_7; // @[d_cache.scala 24:26]
  reg  valid_0_8; // @[d_cache.scala 24:26]
  reg  valid_0_9; // @[d_cache.scala 24:26]
  reg  valid_0_10; // @[d_cache.scala 24:26]
  reg  valid_0_11; // @[d_cache.scala 24:26]
  reg  valid_0_12; // @[d_cache.scala 24:26]
  reg  valid_0_13; // @[d_cache.scala 24:26]
  reg  valid_0_14; // @[d_cache.scala 24:26]
  reg  valid_0_15; // @[d_cache.scala 24:26]
  reg  valid_1_0; // @[d_cache.scala 25:26]
  reg  valid_1_1; // @[d_cache.scala 25:26]
  reg  valid_1_2; // @[d_cache.scala 25:26]
  reg  valid_1_3; // @[d_cache.scala 25:26]
  reg  valid_1_4; // @[d_cache.scala 25:26]
  reg  valid_1_5; // @[d_cache.scala 25:26]
  reg  valid_1_6; // @[d_cache.scala 25:26]
  reg  valid_1_7; // @[d_cache.scala 25:26]
  reg  valid_1_8; // @[d_cache.scala 25:26]
  reg  valid_1_9; // @[d_cache.scala 25:26]
  reg  valid_1_10; // @[d_cache.scala 25:26]
  reg  valid_1_11; // @[d_cache.scala 25:26]
  reg  valid_1_12; // @[d_cache.scala 25:26]
  reg  valid_1_13; // @[d_cache.scala 25:26]
  reg  valid_1_14; // @[d_cache.scala 25:26]
  reg  valid_1_15; // @[d_cache.scala 25:26]
  reg  dirty_0_0; // @[d_cache.scala 26:26]
  reg  dirty_0_1; // @[d_cache.scala 26:26]
  reg  dirty_0_2; // @[d_cache.scala 26:26]
  reg  dirty_0_3; // @[d_cache.scala 26:26]
  reg  dirty_0_4; // @[d_cache.scala 26:26]
  reg  dirty_0_5; // @[d_cache.scala 26:26]
  reg  dirty_0_6; // @[d_cache.scala 26:26]
  reg  dirty_0_7; // @[d_cache.scala 26:26]
  reg  dirty_0_8; // @[d_cache.scala 26:26]
  reg  dirty_0_9; // @[d_cache.scala 26:26]
  reg  dirty_0_10; // @[d_cache.scala 26:26]
  reg  dirty_0_11; // @[d_cache.scala 26:26]
  reg  dirty_0_12; // @[d_cache.scala 26:26]
  reg  dirty_0_13; // @[d_cache.scala 26:26]
  reg  dirty_0_14; // @[d_cache.scala 26:26]
  reg  dirty_0_15; // @[d_cache.scala 26:26]
  reg  dirty_1_0; // @[d_cache.scala 27:26]
  reg  dirty_1_1; // @[d_cache.scala 27:26]
  reg  dirty_1_2; // @[d_cache.scala 27:26]
  reg  dirty_1_3; // @[d_cache.scala 27:26]
  reg  dirty_1_4; // @[d_cache.scala 27:26]
  reg  dirty_1_5; // @[d_cache.scala 27:26]
  reg  dirty_1_6; // @[d_cache.scala 27:26]
  reg  dirty_1_7; // @[d_cache.scala 27:26]
  reg  dirty_1_8; // @[d_cache.scala 27:26]
  reg  dirty_1_9; // @[d_cache.scala 27:26]
  reg  dirty_1_10; // @[d_cache.scala 27:26]
  reg  dirty_1_11; // @[d_cache.scala 27:26]
  reg  dirty_1_12; // @[d_cache.scala 27:26]
  reg  dirty_1_13; // @[d_cache.scala 27:26]
  reg  dirty_1_14; // @[d_cache.scala 27:26]
  reg  dirty_1_15; // @[d_cache.scala 27:26]
  reg [127:0] write_back_data; // @[d_cache.scala 31:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 32:34]
  reg [63:0] receive_data_0; // @[d_cache.scala 37:31]
  reg [63:0] receive_data_1; // @[d_cache.scala 37:31]
  reg [2:0] receive_num; // @[d_cache.scala 38:30]
  reg [1:0] quene_0; // @[d_cache.scala 39:24]
  reg [1:0] quene_1; // @[d_cache.scala 39:24]
  reg [1:0] quene_2; // @[d_cache.scala 39:24]
  reg [1:0] quene_3; // @[d_cache.scala 39:24]
  reg [1:0] quene_4; // @[d_cache.scala 39:24]
  reg [1:0] quene_5; // @[d_cache.scala 39:24]
  reg [1:0] quene_6; // @[d_cache.scala 39:24]
  reg [1:0] quene_7; // @[d_cache.scala 39:24]
  reg [1:0] quene_8; // @[d_cache.scala 39:24]
  reg [1:0] quene_9; // @[d_cache.scala 39:24]
  reg [1:0] quene_10; // @[d_cache.scala 39:24]
  reg [1:0] quene_11; // @[d_cache.scala 39:24]
  reg [1:0] quene_12; // @[d_cache.scala 39:24]
  reg [1:0] quene_13; // @[d_cache.scala 39:24]
  reg [1:0] quene_14; // @[d_cache.scala 39:24]
  reg [1:0] quene_15; // @[d_cache.scala 39:24]
  wire [3:0] offset = io_from_lsu_araddr[3:0]; // @[d_cache.scala 41:36]
  wire [3:0] index = io_from_lsu_araddr[7:4]; // @[d_cache.scala 42:35]
  wire [23:0] tag = io_from_lsu_araddr[31:8]; // @[d_cache.scala 43:33]
  wire [6:0] shift_bit = {offset, 3'h0}; // @[d_cache.scala 45:28]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 51:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 50:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 49:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 48:20]
  wire [31:0] _GEN_1 = 4'h1 == index ? tag_0_1 : tag_0_0; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_2 = 4'h2 == index ? tag_0_2 : _GEN_1; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_3 = 4'h3 == index ? tag_0_3 : _GEN_2; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_4 = 4'h4 == index ? tag_0_4 : _GEN_3; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_5 = 4'h5 == index ? tag_0_5 : _GEN_4; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_6 = 4'h6 == index ? tag_0_6 : _GEN_5; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_7 = 4'h7 == index ? tag_0_7 : _GEN_6; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_8 = 4'h8 == index ? tag_0_8 : _GEN_7; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_9 = 4'h9 == index ? tag_0_9 : _GEN_8; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_10 = 4'ha == index ? tag_0_10 : _GEN_9; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_11 = 4'hb == index ? tag_0_11 : _GEN_10; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_12 = 4'hc == index ? tag_0_12 : _GEN_11; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_13 = 4'hd == index ? tag_0_13 : _GEN_12; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_14 = 4'he == index ? tag_0_14 : _GEN_13; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_15 = 4'hf == index ? tag_0_15 : _GEN_14; // @[d_cache.scala 53:{31,31}]
  wire [31:0] _GEN_2254 = {{8'd0}, tag}; // @[d_cache.scala 53:31]
  wire  _GEN_17 = 4'h1 == index ? valid_0_1 : valid_0_0; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_18 = 4'h2 == index ? valid_0_2 : _GEN_17; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_19 = 4'h3 == index ? valid_0_3 : _GEN_18; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_20 = 4'h4 == index ? valid_0_4 : _GEN_19; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_21 = 4'h5 == index ? valid_0_5 : _GEN_20; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_22 = 4'h6 == index ? valid_0_6 : _GEN_21; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_23 = 4'h7 == index ? valid_0_7 : _GEN_22; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_24 = 4'h8 == index ? valid_0_8 : _GEN_23; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_25 = 4'h9 == index ? valid_0_9 : _GEN_24; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_26 = 4'ha == index ? valid_0_10 : _GEN_25; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_27 = 4'hb == index ? valid_0_11 : _GEN_26; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_28 = 4'hc == index ? valid_0_12 : _GEN_27; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_29 = 4'hd == index ? valid_0_13 : _GEN_28; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_30 = 4'he == index ? valid_0_14 : _GEN_29; // @[d_cache.scala 53:{57,57}]
  wire  _GEN_31 = 4'hf == index ? valid_0_15 : _GEN_30; // @[d_cache.scala 53:{57,57}]
  wire  way0_hit = _GEN_15 == _GEN_2254 & _GEN_31; // @[d_cache.scala 53:40]
  wire [31:0] _GEN_33 = 4'h1 == index ? tag_1_1 : tag_1_0; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_34 = 4'h2 == index ? tag_1_2 : _GEN_33; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_35 = 4'h3 == index ? tag_1_3 : _GEN_34; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_36 = 4'h4 == index ? tag_1_4 : _GEN_35; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_37 = 4'h5 == index ? tag_1_5 : _GEN_36; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_38 = 4'h6 == index ? tag_1_6 : _GEN_37; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_39 = 4'h7 == index ? tag_1_7 : _GEN_38; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_40 = 4'h8 == index ? tag_1_8 : _GEN_39; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_41 = 4'h9 == index ? tag_1_9 : _GEN_40; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_42 = 4'ha == index ? tag_1_10 : _GEN_41; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_43 = 4'hb == index ? tag_1_11 : _GEN_42; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_44 = 4'hc == index ? tag_1_12 : _GEN_43; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_45 = 4'hd == index ? tag_1_13 : _GEN_44; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_46 = 4'he == index ? tag_1_14 : _GEN_45; // @[d_cache.scala 55:{31,31}]
  wire [31:0] _GEN_47 = 4'hf == index ? tag_1_15 : _GEN_46; // @[d_cache.scala 55:{31,31}]
  wire  _GEN_49 = 4'h1 == index ? valid_1_1 : valid_1_0; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_50 = 4'h2 == index ? valid_1_2 : _GEN_49; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_51 = 4'h3 == index ? valid_1_3 : _GEN_50; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_52 = 4'h4 == index ? valid_1_4 : _GEN_51; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_53 = 4'h5 == index ? valid_1_5 : _GEN_52; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_54 = 4'h6 == index ? valid_1_6 : _GEN_53; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_55 = 4'h7 == index ? valid_1_7 : _GEN_54; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_56 = 4'h8 == index ? valid_1_8 : _GEN_55; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_57 = 4'h9 == index ? valid_1_9 : _GEN_56; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_58 = 4'ha == index ? valid_1_10 : _GEN_57; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_59 = 4'hb == index ? valid_1_11 : _GEN_58; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_60 = 4'hc == index ? valid_1_12 : _GEN_59; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_61 = 4'hd == index ? valid_1_13 : _GEN_60; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_62 = 4'he == index ? valid_1_14 : _GEN_61; // @[d_cache.scala 55:{57,57}]
  wire  _GEN_63 = 4'hf == index ? valid_1_15 : _GEN_62; // @[d_cache.scala 55:{57,57}]
  wire  way1_hit = _GEN_47 == _GEN_2254 & _GEN_63; // @[d_cache.scala 55:40]
  wire [1:0] _unuse_way_T_2 = ~_GEN_63 ? 2'h2 : 2'h0; // @[d_cache.scala 58:50]
  wire [1:0] unuse_way = ~_GEN_31 ? 2'h1 : _unuse_way_T_2; // @[d_cache.scala 58:21]
  reg [3:0] state; // @[d_cache.scala 60:24]
  wire  _T_3 = (io_from_lsu_arvalid | io_from_lsu_awvalid) & io_from_lsu_araddr >= 32'ha0000000; // @[d_cache.scala 67:60]
  wire [3:0] _GEN_64 = io_from_lsu_awvalid ? 4'h2 : state; // @[d_cache.scala 71:44 72:23 60:24]
  wire [3:0] _GEN_68 = way1_hit ? 4'h0 : 4'h3; // @[d_cache.scala 82:33 88:23]
  wire [2:0] _GEN_69 = way1_hit ? receive_num : 3'h0; // @[d_cache.scala 38:30 82:33 89:29]
  wire [63:0] _ram_0_T = io_from_lsu_wdata & wmask; // @[d_cache.scala 97:53]
  wire [190:0] _GEN_2487 = {{127'd0}, _ram_0_T}; // @[d_cache.scala 97:62]
  wire [190:0] _ram_0_T_1 = _GEN_2487 << shift_bit; // @[d_cache.scala 97:62]
  wire [190:0] _GEN_2488 = {{127'd0}, wmask}; // @[d_cache.scala 97:102]
  wire [190:0] _ram_0_T_2 = _GEN_2488 << shift_bit; // @[d_cache.scala 97:102]
  wire [190:0] _ram_0_T_3 = ~_ram_0_T_2; // @[d_cache.scala 97:94]
  wire [127:0] _GEN_74 = 4'h1 == index ? ram_0_1 : ram_0_0; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_75 = 4'h2 == index ? ram_0_2 : _GEN_74; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_76 = 4'h3 == index ? ram_0_3 : _GEN_75; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_77 = 4'h4 == index ? ram_0_4 : _GEN_76; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_78 = 4'h5 == index ? ram_0_5 : _GEN_77; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_79 = 4'h6 == index ? ram_0_6 : _GEN_78; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_80 = 4'h7 == index ? ram_0_7 : _GEN_79; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_81 = 4'h8 == index ? ram_0_8 : _GEN_80; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_82 = 4'h9 == index ? ram_0_9 : _GEN_81; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_83 = 4'ha == index ? ram_0_10 : _GEN_82; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_84 = 4'hb == index ? ram_0_11 : _GEN_83; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_85 = 4'hc == index ? ram_0_12 : _GEN_84; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_86 = 4'hd == index ? ram_0_13 : _GEN_85; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_87 = 4'he == index ? ram_0_14 : _GEN_86; // @[d_cache.scala 97:{92,92}]
  wire [127:0] _GEN_88 = 4'hf == index ? ram_0_15 : _GEN_87; // @[d_cache.scala 97:{92,92}]
  wire [190:0] _GEN_2258 = {{63'd0}, _GEN_88}; // @[d_cache.scala 97:92]
  wire [190:0] _ram_0_T_4 = _GEN_2258 & _ram_0_T_3; // @[d_cache.scala 97:92]
  wire [190:0] _ram_0_T_5 = _ram_0_T_1 | _ram_0_T_4; // @[d_cache.scala 97:76]
  wire [127:0] _GEN_89 = 4'h0 == index ? _ram_0_T_5[127:0] : ram_0_0; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_90 = 4'h1 == index ? _ram_0_T_5[127:0] : ram_0_1; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_91 = 4'h2 == index ? _ram_0_T_5[127:0] : ram_0_2; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_92 = 4'h3 == index ? _ram_0_T_5[127:0] : ram_0_3; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_93 = 4'h4 == index ? _ram_0_T_5[127:0] : ram_0_4; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_94 = 4'h5 == index ? _ram_0_T_5[127:0] : ram_0_5; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_95 = 4'h6 == index ? _ram_0_T_5[127:0] : ram_0_6; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_96 = 4'h7 == index ? _ram_0_T_5[127:0] : ram_0_7; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_97 = 4'h8 == index ? _ram_0_T_5[127:0] : ram_0_8; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_98 = 4'h9 == index ? _ram_0_T_5[127:0] : ram_0_9; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_99 = 4'ha == index ? _ram_0_T_5[127:0] : ram_0_10; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_100 = 4'hb == index ? _ram_0_T_5[127:0] : ram_0_11; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_101 = 4'hc == index ? _ram_0_T_5[127:0] : ram_0_12; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_102 = 4'hd == index ? _ram_0_T_5[127:0] : ram_0_13; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_103 = 4'he == index ? _ram_0_T_5[127:0] : ram_0_14; // @[d_cache.scala 19:24 97:{30,30}]
  wire [127:0] _GEN_104 = 4'hf == index ? _ram_0_T_5[127:0] : ram_0_15; // @[d_cache.scala 19:24 97:{30,30}]
  wire  _GEN_2259 = 4'h0 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_105 = 4'h0 == index | dirty_0_0; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2263 = 4'h1 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_106 = 4'h1 == index | dirty_0_1; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2264 = 4'h2 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_107 = 4'h2 == index | dirty_0_2; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2269 = 4'h3 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_108 = 4'h3 == index | dirty_0_3; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2270 = 4'h4 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_109 = 4'h4 == index | dirty_0_4; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2274 = 4'h5 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_110 = 4'h5 == index | dirty_0_5; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2277 = 4'h6 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_111 = 4'h6 == index | dirty_0_6; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2279 = 4'h7 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_112 = 4'h7 == index | dirty_0_7; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2281 = 4'h8 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_113 = 4'h8 == index | dirty_0_8; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2282 = 4'h9 == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_114 = 4'h9 == index | dirty_0_9; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2286 = 4'ha == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_115 = 4'ha == index | dirty_0_10; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2287 = 4'hb == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_116 = 4'hb == index | dirty_0_11; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2292 = 4'hc == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_117 = 4'hc == index | dirty_0_12; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2293 = 4'hd == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_118 = 4'hd == index | dirty_0_13; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2297 = 4'he == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_119 = 4'he == index | dirty_0_14; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_2301 = 4'hf == index; // @[d_cache.scala 26:26 98:{32,32}]
  wire  _GEN_120 = 4'hf == index | dirty_0_15; // @[d_cache.scala 26:26 98:{32,32}]
  wire [127:0] _GEN_122 = 4'h1 == index ? ram_1_1 : ram_1_0; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_123 = 4'h2 == index ? ram_1_2 : _GEN_122; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_124 = 4'h3 == index ? ram_1_3 : _GEN_123; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_125 = 4'h4 == index ? ram_1_4 : _GEN_124; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_126 = 4'h5 == index ? ram_1_5 : _GEN_125; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_127 = 4'h6 == index ? ram_1_6 : _GEN_126; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_128 = 4'h7 == index ? ram_1_7 : _GEN_127; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_129 = 4'h8 == index ? ram_1_8 : _GEN_128; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_130 = 4'h9 == index ? ram_1_9 : _GEN_129; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_131 = 4'ha == index ? ram_1_10 : _GEN_130; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_132 = 4'hb == index ? ram_1_11 : _GEN_131; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_133 = 4'hc == index ? ram_1_12 : _GEN_132; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_134 = 4'hd == index ? ram_1_13 : _GEN_133; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_135 = 4'he == index ? ram_1_14 : _GEN_134; // @[d_cache.scala 105:{92,92}]
  wire [127:0] _GEN_136 = 4'hf == index ? ram_1_15 : _GEN_135; // @[d_cache.scala 105:{92,92}]
  wire [190:0] _GEN_2303 = {{63'd0}, _GEN_136}; // @[d_cache.scala 105:92]
  wire [190:0] _ram_1_T_4 = _GEN_2303 & _ram_0_T_3; // @[d_cache.scala 105:92]
  wire [190:0] _ram_1_T_5 = _ram_0_T_1 | _ram_1_T_4; // @[d_cache.scala 105:76]
  wire [127:0] _GEN_137 = 4'h0 == index ? _ram_1_T_5[127:0] : ram_1_0; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_138 = 4'h1 == index ? _ram_1_T_5[127:0] : ram_1_1; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_139 = 4'h2 == index ? _ram_1_T_5[127:0] : ram_1_2; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_140 = 4'h3 == index ? _ram_1_T_5[127:0] : ram_1_3; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_141 = 4'h4 == index ? _ram_1_T_5[127:0] : ram_1_4; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_142 = 4'h5 == index ? _ram_1_T_5[127:0] : ram_1_5; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_143 = 4'h6 == index ? _ram_1_T_5[127:0] : ram_1_6; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_144 = 4'h7 == index ? _ram_1_T_5[127:0] : ram_1_7; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_145 = 4'h8 == index ? _ram_1_T_5[127:0] : ram_1_8; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_146 = 4'h9 == index ? _ram_1_T_5[127:0] : ram_1_9; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_147 = 4'ha == index ? _ram_1_T_5[127:0] : ram_1_10; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_148 = 4'hb == index ? _ram_1_T_5[127:0] : ram_1_11; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_149 = 4'hc == index ? _ram_1_T_5[127:0] : ram_1_12; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_150 = 4'hd == index ? _ram_1_T_5[127:0] : ram_1_13; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_151 = 4'he == index ? _ram_1_T_5[127:0] : ram_1_14; // @[d_cache.scala 105:{30,30} 20:24]
  wire [127:0] _GEN_152 = 4'hf == index ? _ram_1_T_5[127:0] : ram_1_15; // @[d_cache.scala 105:{30,30} 20:24]
  wire  _GEN_153 = _GEN_2259 | dirty_1_0; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_154 = _GEN_2263 | dirty_1_1; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_155 = _GEN_2264 | dirty_1_2; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_156 = _GEN_2269 | dirty_1_3; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_157 = _GEN_2270 | dirty_1_4; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_158 = _GEN_2274 | dirty_1_5; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_159 = _GEN_2277 | dirty_1_6; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_160 = _GEN_2279 | dirty_1_7; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_161 = _GEN_2281 | dirty_1_8; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_162 = _GEN_2282 | dirty_1_9; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_163 = _GEN_2286 | dirty_1_10; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_164 = _GEN_2287 | dirty_1_11; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_165 = _GEN_2292 | dirty_1_12; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_166 = _GEN_2293 | dirty_1_13; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_167 = _GEN_2297 | dirty_1_14; // @[d_cache.scala 106:{32,32} 27:26]
  wire  _GEN_168 = _GEN_2301 | dirty_1_15; // @[d_cache.scala 106:{32,32} 27:26]
  wire [3:0] _GEN_169 = way1_hit ? 4'h0 : 4'h4; // @[d_cache.scala 100:33 108:23]
  wire [127:0] _GEN_170 = way1_hit ? _GEN_137 : ram_1_0; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_171 = way1_hit ? _GEN_138 : ram_1_1; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_172 = way1_hit ? _GEN_139 : ram_1_2; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_173 = way1_hit ? _GEN_140 : ram_1_3; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_174 = way1_hit ? _GEN_141 : ram_1_4; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_175 = way1_hit ? _GEN_142 : ram_1_5; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_176 = way1_hit ? _GEN_143 : ram_1_6; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_177 = way1_hit ? _GEN_144 : ram_1_7; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_178 = way1_hit ? _GEN_145 : ram_1_8; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_179 = way1_hit ? _GEN_146 : ram_1_9; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_180 = way1_hit ? _GEN_147 : ram_1_10; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_181 = way1_hit ? _GEN_148 : ram_1_11; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_182 = way1_hit ? _GEN_149 : ram_1_12; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_183 = way1_hit ? _GEN_150 : ram_1_13; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_184 = way1_hit ? _GEN_151 : ram_1_14; // @[d_cache.scala 100:33 20:24]
  wire [127:0] _GEN_185 = way1_hit ? _GEN_152 : ram_1_15; // @[d_cache.scala 100:33 20:24]
  wire  _GEN_186 = way1_hit ? _GEN_153 : dirty_1_0; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_187 = way1_hit ? _GEN_154 : dirty_1_1; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_188 = way1_hit ? _GEN_155 : dirty_1_2; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_189 = way1_hit ? _GEN_156 : dirty_1_3; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_190 = way1_hit ? _GEN_157 : dirty_1_4; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_191 = way1_hit ? _GEN_158 : dirty_1_5; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_192 = way1_hit ? _GEN_159 : dirty_1_6; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_193 = way1_hit ? _GEN_160 : dirty_1_7; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_194 = way1_hit ? _GEN_161 : dirty_1_8; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_195 = way1_hit ? _GEN_162 : dirty_1_9; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_196 = way1_hit ? _GEN_163 : dirty_1_10; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_197 = way1_hit ? _GEN_164 : dirty_1_11; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_198 = way1_hit ? _GEN_165 : dirty_1_12; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_199 = way1_hit ? _GEN_166 : dirty_1_13; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_200 = way1_hit ? _GEN_167 : dirty_1_14; // @[d_cache.scala 100:33 27:26]
  wire  _GEN_201 = way1_hit ? _GEN_168 : dirty_1_15; // @[d_cache.scala 100:33 27:26]
  wire [3:0] _GEN_202 = way0_hit ? 4'h0 : _GEN_169; // @[d_cache.scala 93:27]
  wire [127:0] _GEN_203 = way0_hit ? _GEN_89 : ram_0_0; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_204 = way0_hit ? _GEN_90 : ram_0_1; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_205 = way0_hit ? _GEN_91 : ram_0_2; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_206 = way0_hit ? _GEN_92 : ram_0_3; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_207 = way0_hit ? _GEN_93 : ram_0_4; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_208 = way0_hit ? _GEN_94 : ram_0_5; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_209 = way0_hit ? _GEN_95 : ram_0_6; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_210 = way0_hit ? _GEN_96 : ram_0_7; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_211 = way0_hit ? _GEN_97 : ram_0_8; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_212 = way0_hit ? _GEN_98 : ram_0_9; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_213 = way0_hit ? _GEN_99 : ram_0_10; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_214 = way0_hit ? _GEN_100 : ram_0_11; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_215 = way0_hit ? _GEN_101 : ram_0_12; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_216 = way0_hit ? _GEN_102 : ram_0_13; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_217 = way0_hit ? _GEN_103 : ram_0_14; // @[d_cache.scala 19:24 93:27]
  wire [127:0] _GEN_218 = way0_hit ? _GEN_104 : ram_0_15; // @[d_cache.scala 19:24 93:27]
  wire  _GEN_219 = way0_hit ? _GEN_105 : dirty_0_0; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_220 = way0_hit ? _GEN_106 : dirty_0_1; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_221 = way0_hit ? _GEN_107 : dirty_0_2; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_222 = way0_hit ? _GEN_108 : dirty_0_3; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_223 = way0_hit ? _GEN_109 : dirty_0_4; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_224 = way0_hit ? _GEN_110 : dirty_0_5; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_225 = way0_hit ? _GEN_111 : dirty_0_6; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_226 = way0_hit ? _GEN_112 : dirty_0_7; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_227 = way0_hit ? _GEN_113 : dirty_0_8; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_228 = way0_hit ? _GEN_114 : dirty_0_9; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_229 = way0_hit ? _GEN_115 : dirty_0_10; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_230 = way0_hit ? _GEN_116 : dirty_0_11; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_231 = way0_hit ? _GEN_117 : dirty_0_12; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_232 = way0_hit ? _GEN_118 : dirty_0_13; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_233 = way0_hit ? _GEN_119 : dirty_0_14; // @[d_cache.scala 26:26 93:27]
  wire  _GEN_234 = way0_hit ? _GEN_120 : dirty_0_15; // @[d_cache.scala 26:26 93:27]
  wire [127:0] _GEN_235 = way0_hit ? ram_1_0 : _GEN_170; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_236 = way0_hit ? ram_1_1 : _GEN_171; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_237 = way0_hit ? ram_1_2 : _GEN_172; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_238 = way0_hit ? ram_1_3 : _GEN_173; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_239 = way0_hit ? ram_1_4 : _GEN_174; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_240 = way0_hit ? ram_1_5 : _GEN_175; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_241 = way0_hit ? ram_1_6 : _GEN_176; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_242 = way0_hit ? ram_1_7 : _GEN_177; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_243 = way0_hit ? ram_1_8 : _GEN_178; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_244 = way0_hit ? ram_1_9 : _GEN_179; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_245 = way0_hit ? ram_1_10 : _GEN_180; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_246 = way0_hit ? ram_1_11 : _GEN_181; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_247 = way0_hit ? ram_1_12 : _GEN_182; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_248 = way0_hit ? ram_1_13 : _GEN_183; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_249 = way0_hit ? ram_1_14 : _GEN_184; // @[d_cache.scala 20:24 93:27]
  wire [127:0] _GEN_250 = way0_hit ? ram_1_15 : _GEN_185; // @[d_cache.scala 20:24 93:27]
  wire  _GEN_251 = way0_hit ? dirty_1_0 : _GEN_186; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_252 = way0_hit ? dirty_1_1 : _GEN_187; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_253 = way0_hit ? dirty_1_2 : _GEN_188; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_254 = way0_hit ? dirty_1_3 : _GEN_189; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_255 = way0_hit ? dirty_1_4 : _GEN_190; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_256 = way0_hit ? dirty_1_5 : _GEN_191; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_257 = way0_hit ? dirty_1_6 : _GEN_192; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_258 = way0_hit ? dirty_1_7 : _GEN_193; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_259 = way0_hit ? dirty_1_8 : _GEN_194; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_260 = way0_hit ? dirty_1_9 : _GEN_195; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_261 = way0_hit ? dirty_1_10 : _GEN_196; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_262 = way0_hit ? dirty_1_11 : _GEN_197; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_263 = way0_hit ? dirty_1_12 : _GEN_198; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_264 = way0_hit ? dirty_1_13 : _GEN_199; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_265 = way0_hit ? dirty_1_14 : _GEN_200; // @[d_cache.scala 27:26 93:27]
  wire  _GEN_266 = way0_hit ? dirty_1_15 : _GEN_201; // @[d_cache.scala 27:26 93:27]
  wire [63:0] _GEN_267 = ~receive_num[0] ? io_from_axi_rdata : receive_data_0; // @[d_cache.scala 113:{43,43} 37:31]
  wire [63:0] _GEN_268 = receive_num[0] ? io_from_axi_rdata : receive_data_1; // @[d_cache.scala 113:{43,43} 37:31]
  wire [2:0] _receive_num_T_1 = receive_num + 3'h1; // @[d_cache.scala 114:44]
  wire [3:0] _GEN_269 = io_from_axi_rlast ? 4'h5 : state; // @[d_cache.scala 115:40 116:27 60:24]
  wire [63:0] _GEN_270 = io_from_axi_rvalid ? _GEN_267 : receive_data_0; // @[d_cache.scala 112:37 37:31]
  wire [63:0] _GEN_271 = io_from_axi_rvalid ? _GEN_268 : receive_data_1; // @[d_cache.scala 112:37 37:31]
  wire [2:0] _GEN_272 = io_from_axi_rvalid ? _receive_num_T_1 : receive_num; // @[d_cache.scala 112:37 114:29 38:30]
  wire [3:0] _GEN_273 = io_from_axi_rvalid ? _GEN_269 : state; // @[d_cache.scala 112:37 60:24]
  wire [3:0] _GEN_274 = io_from_axi_bvalid ? 4'h0 : state; // @[d_cache.scala 121:59 122:23 60:24]
  wire [127:0] _ram_0_T_6 = {receive_data_1,receive_data_0}; // @[Cat.scala 31:58]
  wire [127:0] _GEN_275 = 4'h0 == index ? _ram_0_T_6 : ram_0_0; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_276 = 4'h1 == index ? _ram_0_T_6 : ram_0_1; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_277 = 4'h2 == index ? _ram_0_T_6 : ram_0_2; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_278 = 4'h3 == index ? _ram_0_T_6 : ram_0_3; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_279 = 4'h4 == index ? _ram_0_T_6 : ram_0_4; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_280 = 4'h5 == index ? _ram_0_T_6 : ram_0_5; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_281 = 4'h6 == index ? _ram_0_T_6 : ram_0_6; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_282 = 4'h7 == index ? _ram_0_T_6 : ram_0_7; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_283 = 4'h8 == index ? _ram_0_T_6 : ram_0_8; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_284 = 4'h9 == index ? _ram_0_T_6 : ram_0_9; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_285 = 4'ha == index ? _ram_0_T_6 : ram_0_10; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_286 = 4'hb == index ? _ram_0_T_6 : ram_0_11; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_287 = 4'hc == index ? _ram_0_T_6 : ram_0_12; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_288 = 4'hd == index ? _ram_0_T_6 : ram_0_13; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_289 = 4'he == index ? _ram_0_T_6 : ram_0_14; // @[d_cache.scala 128:{30,30} 19:24]
  wire [127:0] _GEN_290 = 4'hf == index ? _ram_0_T_6 : ram_0_15; // @[d_cache.scala 128:{30,30} 19:24]
  wire [31:0] _GEN_291 = 4'h0 == index ? _GEN_2254 : tag_0_0; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_292 = 4'h1 == index ? _GEN_2254 : tag_0_1; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_293 = 4'h2 == index ? _GEN_2254 : tag_0_2; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_294 = 4'h3 == index ? _GEN_2254 : tag_0_3; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_295 = 4'h4 == index ? _GEN_2254 : tag_0_4; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_296 = 4'h5 == index ? _GEN_2254 : tag_0_5; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_297 = 4'h6 == index ? _GEN_2254 : tag_0_6; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_298 = 4'h7 == index ? _GEN_2254 : tag_0_7; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_299 = 4'h8 == index ? _GEN_2254 : tag_0_8; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_300 = 4'h9 == index ? _GEN_2254 : tag_0_9; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_301 = 4'ha == index ? _GEN_2254 : tag_0_10; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_302 = 4'hb == index ? _GEN_2254 : tag_0_11; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_303 = 4'hc == index ? _GEN_2254 : tag_0_12; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_304 = 4'hd == index ? _GEN_2254 : tag_0_13; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_305 = 4'he == index ? _GEN_2254 : tag_0_14; // @[d_cache.scala 129:{30,30} 22:24]
  wire [31:0] _GEN_306 = 4'hf == index ? _GEN_2254 : tag_0_15; // @[d_cache.scala 129:{30,30} 22:24]
  wire  _GEN_307 = _GEN_2259 | valid_0_0; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_308 = _GEN_2263 | valid_0_1; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_309 = _GEN_2264 | valid_0_2; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_310 = _GEN_2269 | valid_0_3; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_311 = _GEN_2270 | valid_0_4; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_312 = _GEN_2274 | valid_0_5; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_313 = _GEN_2277 | valid_0_6; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_314 = _GEN_2279 | valid_0_7; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_315 = _GEN_2281 | valid_0_8; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_316 = _GEN_2282 | valid_0_9; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_317 = _GEN_2286 | valid_0_10; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_318 = _GEN_2287 | valid_0_11; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_319 = _GEN_2292 | valid_0_12; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_320 = _GEN_2293 | valid_0_13; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_321 = _GEN_2297 | valid_0_14; // @[d_cache.scala 130:{32,32} 24:26]
  wire  _GEN_322 = _GEN_2301 | valid_0_15; // @[d_cache.scala 130:{32,32} 24:26]
  wire [1:0] _GEN_324 = 4'h1 == index ? quene_1 : quene_0; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_325 = 4'h2 == index ? quene_2 : _GEN_324; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_326 = 4'h3 == index ? quene_3 : _GEN_325; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_327 = 4'h4 == index ? quene_4 : _GEN_326; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_328 = 4'h5 == index ? quene_5 : _GEN_327; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_329 = 4'h6 == index ? quene_6 : _GEN_328; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_330 = 4'h7 == index ? quene_7 : _GEN_329; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_331 = 4'h8 == index ? quene_8 : _GEN_330; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_332 = 4'h9 == index ? quene_9 : _GEN_331; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_333 = 4'ha == index ? quene_10 : _GEN_332; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_334 = 4'hb == index ? quene_11 : _GEN_333; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_335 = 4'hc == index ? quene_12 : _GEN_334; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_336 = 4'hd == index ? quene_13 : _GEN_335; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_337 = 4'he == index ? quene_14 : _GEN_336; // @[d_cache.scala 131:{46,46}]
  wire [1:0] _GEN_338 = 4'hf == index ? quene_15 : _GEN_337; // @[d_cache.scala 131:{46,46}]
  wire [2:0] _quene_T = {_GEN_338, 1'h0}; // @[d_cache.scala 131:46]
  wire [1:0] _GEN_339 = 4'h0 == index ? _quene_T[1:0] : quene_0; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_340 = 4'h1 == index ? _quene_T[1:0] : quene_1; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_341 = 4'h2 == index ? _quene_T[1:0] : quene_2; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_342 = 4'h3 == index ? _quene_T[1:0] : quene_3; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_343 = 4'h4 == index ? _quene_T[1:0] : quene_4; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_344 = 4'h5 == index ? _quene_T[1:0] : quene_5; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_345 = 4'h6 == index ? _quene_T[1:0] : quene_6; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_346 = 4'h7 == index ? _quene_T[1:0] : quene_7; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_347 = 4'h8 == index ? _quene_T[1:0] : quene_8; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_348 = 4'h9 == index ? _quene_T[1:0] : quene_9; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_349 = 4'ha == index ? _quene_T[1:0] : quene_10; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_350 = 4'hb == index ? _quene_T[1:0] : quene_11; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_351 = 4'hc == index ? _quene_T[1:0] : quene_12; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_352 = 4'hd == index ? _quene_T[1:0] : quene_13; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_353 = 4'he == index ? _quene_T[1:0] : quene_14; // @[d_cache.scala 131:{30,30} 39:24]
  wire [1:0] _GEN_354 = 4'hf == index ? _quene_T[1:0] : quene_15; // @[d_cache.scala 131:{30,30} 39:24]
  wire [127:0] _GEN_355 = 4'h0 == index ? _ram_0_T_6 : ram_1_0; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_356 = 4'h1 == index ? _ram_0_T_6 : ram_1_1; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_357 = 4'h2 == index ? _ram_0_T_6 : ram_1_2; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_358 = 4'h3 == index ? _ram_0_T_6 : ram_1_3; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_359 = 4'h4 == index ? _ram_0_T_6 : ram_1_4; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_360 = 4'h5 == index ? _ram_0_T_6 : ram_1_5; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_361 = 4'h6 == index ? _ram_0_T_6 : ram_1_6; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_362 = 4'h7 == index ? _ram_0_T_6 : ram_1_7; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_363 = 4'h8 == index ? _ram_0_T_6 : ram_1_8; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_364 = 4'h9 == index ? _ram_0_T_6 : ram_1_9; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_365 = 4'ha == index ? _ram_0_T_6 : ram_1_10; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_366 = 4'hb == index ? _ram_0_T_6 : ram_1_11; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_367 = 4'hc == index ? _ram_0_T_6 : ram_1_12; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_368 = 4'hd == index ? _ram_0_T_6 : ram_1_13; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_369 = 4'he == index ? _ram_0_T_6 : ram_1_14; // @[d_cache.scala 134:{30,30} 20:24]
  wire [127:0] _GEN_370 = 4'hf == index ? _ram_0_T_6 : ram_1_15; // @[d_cache.scala 134:{30,30} 20:24]
  wire [31:0] _GEN_371 = 4'h0 == index ? _GEN_2254 : tag_1_0; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_372 = 4'h1 == index ? _GEN_2254 : tag_1_1; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_373 = 4'h2 == index ? _GEN_2254 : tag_1_2; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_374 = 4'h3 == index ? _GEN_2254 : tag_1_3; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_375 = 4'h4 == index ? _GEN_2254 : tag_1_4; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_376 = 4'h5 == index ? _GEN_2254 : tag_1_5; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_377 = 4'h6 == index ? _GEN_2254 : tag_1_6; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_378 = 4'h7 == index ? _GEN_2254 : tag_1_7; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_379 = 4'h8 == index ? _GEN_2254 : tag_1_8; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_380 = 4'h9 == index ? _GEN_2254 : tag_1_9; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_381 = 4'ha == index ? _GEN_2254 : tag_1_10; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_382 = 4'hb == index ? _GEN_2254 : tag_1_11; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_383 = 4'hc == index ? _GEN_2254 : tag_1_12; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_384 = 4'hd == index ? _GEN_2254 : tag_1_13; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_385 = 4'he == index ? _GEN_2254 : tag_1_14; // @[d_cache.scala 135:{30,30} 23:24]
  wire [31:0] _GEN_386 = 4'hf == index ? _GEN_2254 : tag_1_15; // @[d_cache.scala 135:{30,30} 23:24]
  wire  _GEN_387 = _GEN_2259 | valid_1_0; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_388 = _GEN_2263 | valid_1_1; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_389 = _GEN_2264 | valid_1_2; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_390 = _GEN_2269 | valid_1_3; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_391 = _GEN_2270 | valid_1_4; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_392 = _GEN_2274 | valid_1_5; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_393 = _GEN_2277 | valid_1_6; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_394 = _GEN_2279 | valid_1_7; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_395 = _GEN_2281 | valid_1_8; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_396 = _GEN_2282 | valid_1_9; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_397 = _GEN_2286 | valid_1_10; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_398 = _GEN_2287 | valid_1_11; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_399 = _GEN_2292 | valid_1_12; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_400 = _GEN_2293 | valid_1_13; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_401 = _GEN_2297 | valid_1_14; // @[d_cache.scala 136:{32,32} 25:26]
  wire  _GEN_402 = _GEN_2301 | valid_1_15; // @[d_cache.scala 136:{32,32} 25:26]
  wire [2:0] _quene_T_2 = _quene_T | 3'h1; // @[d_cache.scala 137:55]
  wire [1:0] _GEN_403 = 4'h0 == index ? _quene_T_2[1:0] : quene_0; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_404 = 4'h1 == index ? _quene_T_2[1:0] : quene_1; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_405 = 4'h2 == index ? _quene_T_2[1:0] : quene_2; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_406 = 4'h3 == index ? _quene_T_2[1:0] : quene_3; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_407 = 4'h4 == index ? _quene_T_2[1:0] : quene_4; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_408 = 4'h5 == index ? _quene_T_2[1:0] : quene_5; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_409 = 4'h6 == index ? _quene_T_2[1:0] : quene_6; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_410 = 4'h7 == index ? _quene_T_2[1:0] : quene_7; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_411 = 4'h8 == index ? _quene_T_2[1:0] : quene_8; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_412 = 4'h9 == index ? _quene_T_2[1:0] : quene_9; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_413 = 4'ha == index ? _quene_T_2[1:0] : quene_10; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_414 = 4'hb == index ? _quene_T_2[1:0] : quene_11; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_415 = 4'hc == index ? _quene_T_2[1:0] : quene_12; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_416 = 4'hd == index ? _quene_T_2[1:0] : quene_13; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_417 = 4'he == index ? _quene_T_2[1:0] : quene_14; // @[d_cache.scala 137:{30,30} 39:24]
  wire [1:0] _GEN_418 = 4'hf == index ? _quene_T_2[1:0] : quene_15; // @[d_cache.scala 137:{30,30} 39:24]
  wire  _GEN_420 = 4'h1 == index ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_421 = 4'h2 == index ? dirty_0_2 : _GEN_420; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_422 = 4'h3 == index ? dirty_0_3 : _GEN_421; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_423 = 4'h4 == index ? dirty_0_4 : _GEN_422; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_424 = 4'h5 == index ? dirty_0_5 : _GEN_423; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_425 = 4'h6 == index ? dirty_0_6 : _GEN_424; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_426 = 4'h7 == index ? dirty_0_7 : _GEN_425; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_427 = 4'h8 == index ? dirty_0_8 : _GEN_426; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_428 = 4'h9 == index ? dirty_0_9 : _GEN_427; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_429 = 4'ha == index ? dirty_0_10 : _GEN_428; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_430 = 4'hb == index ? dirty_0_11 : _GEN_429; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_431 = 4'hc == index ? dirty_0_12 : _GEN_430; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_432 = 4'hd == index ? dirty_0_13 : _GEN_431; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_433 = 4'he == index ? dirty_0_14 : _GEN_432; // @[d_cache.scala 141:{40,40}]
  wire  _GEN_434 = 4'hf == index ? dirty_0_15 : _GEN_433; // @[d_cache.scala 141:{40,40}]
  wire [39:0] _write_back_addr_T_1 = {_GEN_15,index,4'h0}; // @[Cat.scala 31:58]
  wire  _GEN_467 = 4'h0 == index ? 1'h0 : dirty_0_0; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_468 = 4'h1 == index ? 1'h0 : dirty_0_1; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_469 = 4'h2 == index ? 1'h0 : dirty_0_2; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_470 = 4'h3 == index ? 1'h0 : dirty_0_3; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_471 = 4'h4 == index ? 1'h0 : dirty_0_4; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_472 = 4'h5 == index ? 1'h0 : dirty_0_5; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_473 = 4'h6 == index ? 1'h0 : dirty_0_6; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_474 = 4'h7 == index ? 1'h0 : dirty_0_7; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_475 = 4'h8 == index ? 1'h0 : dirty_0_8; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_476 = 4'h9 == index ? 1'h0 : dirty_0_9; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_477 = 4'ha == index ? 1'h0 : dirty_0_10; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_478 = 4'hb == index ? 1'h0 : dirty_0_11; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_479 = 4'hc == index ? 1'h0 : dirty_0_12; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_480 = 4'hd == index ? 1'h0 : dirty_0_13; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_481 = 4'he == index ? 1'h0 : dirty_0_14; // @[d_cache.scala 146:{40,40} 26:26]
  wire  _GEN_482 = 4'hf == index ? 1'h0 : dirty_0_15; // @[d_cache.scala 146:{40,40} 26:26]
  wire [127:0] _GEN_579 = _GEN_434 ? _GEN_88 : write_back_data; // @[d_cache.scala 141:47 142:41 31:34]
  wire [39:0] _GEN_580 = _GEN_434 ? _write_back_addr_T_1 : {{8'd0}, write_back_addr}; // @[d_cache.scala 141:47 143:41 32:34]
  wire [127:0] _GEN_581 = _GEN_434 ? _GEN_275 : _GEN_275; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_582 = _GEN_434 ? _GEN_276 : _GEN_276; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_583 = _GEN_434 ? _GEN_277 : _GEN_277; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_584 = _GEN_434 ? _GEN_278 : _GEN_278; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_585 = _GEN_434 ? _GEN_279 : _GEN_279; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_586 = _GEN_434 ? _GEN_280 : _GEN_280; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_587 = _GEN_434 ? _GEN_281 : _GEN_281; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_588 = _GEN_434 ? _GEN_282 : _GEN_282; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_589 = _GEN_434 ? _GEN_283 : _GEN_283; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_590 = _GEN_434 ? _GEN_284 : _GEN_284; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_591 = _GEN_434 ? _GEN_285 : _GEN_285; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_592 = _GEN_434 ? _GEN_286 : _GEN_286; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_593 = _GEN_434 ? _GEN_287 : _GEN_287; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_594 = _GEN_434 ? _GEN_288 : _GEN_288; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_595 = _GEN_434 ? _GEN_289 : _GEN_289; // @[d_cache.scala 141:47]
  wire [127:0] _GEN_596 = _GEN_434 ? _GEN_290 : _GEN_290; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_597 = _GEN_434 ? _GEN_291 : _GEN_291; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_598 = _GEN_434 ? _GEN_292 : _GEN_292; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_599 = _GEN_434 ? _GEN_293 : _GEN_293; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_600 = _GEN_434 ? _GEN_294 : _GEN_294; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_601 = _GEN_434 ? _GEN_295 : _GEN_295; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_602 = _GEN_434 ? _GEN_296 : _GEN_296; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_603 = _GEN_434 ? _GEN_297 : _GEN_297; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_604 = _GEN_434 ? _GEN_298 : _GEN_298; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_605 = _GEN_434 ? _GEN_299 : _GEN_299; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_606 = _GEN_434 ? _GEN_300 : _GEN_300; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_607 = _GEN_434 ? _GEN_301 : _GEN_301; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_608 = _GEN_434 ? _GEN_302 : _GEN_302; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_609 = _GEN_434 ? _GEN_303 : _GEN_303; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_610 = _GEN_434 ? _GEN_304 : _GEN_304; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_611 = _GEN_434 ? _GEN_305 : _GEN_305; // @[d_cache.scala 141:47]
  wire [31:0] _GEN_612 = _GEN_434 ? _GEN_306 : _GEN_306; // @[d_cache.scala 141:47]
  wire  _GEN_613 = _GEN_434 ? _GEN_467 : dirty_0_0; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_614 = _GEN_434 ? _GEN_468 : dirty_0_1; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_615 = _GEN_434 ? _GEN_469 : dirty_0_2; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_616 = _GEN_434 ? _GEN_470 : dirty_0_3; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_617 = _GEN_434 ? _GEN_471 : dirty_0_4; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_618 = _GEN_434 ? _GEN_472 : dirty_0_5; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_619 = _GEN_434 ? _GEN_473 : dirty_0_6; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_620 = _GEN_434 ? _GEN_474 : dirty_0_7; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_621 = _GEN_434 ? _GEN_475 : dirty_0_8; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_622 = _GEN_434 ? _GEN_476 : dirty_0_9; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_623 = _GEN_434 ? _GEN_477 : dirty_0_10; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_624 = _GEN_434 ? _GEN_478 : dirty_0_11; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_625 = _GEN_434 ? _GEN_479 : dirty_0_12; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_626 = _GEN_434 ? _GEN_480 : dirty_0_13; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_627 = _GEN_434 ? _GEN_481 : dirty_0_14; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_628 = _GEN_434 ? _GEN_482 : dirty_0_15; // @[d_cache.scala 141:47 26:26]
  wire  _GEN_629 = _GEN_434 ? _GEN_307 : _GEN_307; // @[d_cache.scala 141:47]
  wire  _GEN_630 = _GEN_434 ? _GEN_308 : _GEN_308; // @[d_cache.scala 141:47]
  wire  _GEN_631 = _GEN_434 ? _GEN_309 : _GEN_309; // @[d_cache.scala 141:47]
  wire  _GEN_632 = _GEN_434 ? _GEN_310 : _GEN_310; // @[d_cache.scala 141:47]
  wire  _GEN_633 = _GEN_434 ? _GEN_311 : _GEN_311; // @[d_cache.scala 141:47]
  wire  _GEN_634 = _GEN_434 ? _GEN_312 : _GEN_312; // @[d_cache.scala 141:47]
  wire  _GEN_635 = _GEN_434 ? _GEN_313 : _GEN_313; // @[d_cache.scala 141:47]
  wire  _GEN_636 = _GEN_434 ? _GEN_314 : _GEN_314; // @[d_cache.scala 141:47]
  wire  _GEN_637 = _GEN_434 ? _GEN_315 : _GEN_315; // @[d_cache.scala 141:47]
  wire  _GEN_638 = _GEN_434 ? _GEN_316 : _GEN_316; // @[d_cache.scala 141:47]
  wire  _GEN_639 = _GEN_434 ? _GEN_317 : _GEN_317; // @[d_cache.scala 141:47]
  wire  _GEN_640 = _GEN_434 ? _GEN_318 : _GEN_318; // @[d_cache.scala 141:47]
  wire  _GEN_641 = _GEN_434 ? _GEN_319 : _GEN_319; // @[d_cache.scala 141:47]
  wire  _GEN_642 = _GEN_434 ? _GEN_320 : _GEN_320; // @[d_cache.scala 141:47]
  wire  _GEN_643 = _GEN_434 ? _GEN_321 : _GEN_321; // @[d_cache.scala 141:47]
  wire  _GEN_644 = _GEN_434 ? _GEN_322 : _GEN_322; // @[d_cache.scala 141:47]
  wire [3:0] _GEN_645 = _GEN_434 ? 4'h6 : 4'h1; // @[d_cache.scala 141:47 148:31 151:31]
  wire [1:0] _GEN_646 = _GEN_434 ? _GEN_339 : _GEN_339; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_647 = _GEN_434 ? _GEN_340 : _GEN_340; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_648 = _GEN_434 ? _GEN_341 : _GEN_341; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_649 = _GEN_434 ? _GEN_342 : _GEN_342; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_650 = _GEN_434 ? _GEN_343 : _GEN_343; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_651 = _GEN_434 ? _GEN_344 : _GEN_344; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_652 = _GEN_434 ? _GEN_345 : _GEN_345; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_653 = _GEN_434 ? _GEN_346 : _GEN_346; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_654 = _GEN_434 ? _GEN_347 : _GEN_347; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_655 = _GEN_434 ? _GEN_348 : _GEN_348; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_656 = _GEN_434 ? _GEN_349 : _GEN_349; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_657 = _GEN_434 ? _GEN_350 : _GEN_350; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_658 = _GEN_434 ? _GEN_351 : _GEN_351; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_659 = _GEN_434 ? _GEN_352 : _GEN_352; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_660 = _GEN_434 ? _GEN_353 : _GEN_353; // @[d_cache.scala 141:47]
  wire [1:0] _GEN_661 = _GEN_434 ? _GEN_354 : _GEN_354; // @[d_cache.scala 141:47]
  wire  _GEN_663 = 4'h1 == index ? dirty_1_1 : dirty_1_0; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_664 = 4'h2 == index ? dirty_1_2 : _GEN_663; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_665 = 4'h3 == index ? dirty_1_3 : _GEN_664; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_666 = 4'h4 == index ? dirty_1_4 : _GEN_665; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_667 = 4'h5 == index ? dirty_1_5 : _GEN_666; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_668 = 4'h6 == index ? dirty_1_6 : _GEN_667; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_669 = 4'h7 == index ? dirty_1_7 : _GEN_668; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_670 = 4'h8 == index ? dirty_1_8 : _GEN_669; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_671 = 4'h9 == index ? dirty_1_9 : _GEN_670; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_672 = 4'ha == index ? dirty_1_10 : _GEN_671; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_673 = 4'hb == index ? dirty_1_11 : _GEN_672; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_674 = 4'hc == index ? dirty_1_12 : _GEN_673; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_675 = 4'hd == index ? dirty_1_13 : _GEN_674; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_676 = 4'he == index ? dirty_1_14 : _GEN_675; // @[d_cache.scala 158:{40,40}]
  wire  _GEN_677 = 4'hf == index ? dirty_1_15 : _GEN_676; // @[d_cache.scala 158:{40,40}]
  wire [39:0] _write_back_addr_T_3 = {_GEN_47,index,4'h0}; // @[Cat.scala 31:58]
  wire  _GEN_710 = 4'h0 == index ? 1'h0 : dirty_1_0; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_711 = 4'h1 == index ? 1'h0 : dirty_1_1; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_712 = 4'h2 == index ? 1'h0 : dirty_1_2; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_713 = 4'h3 == index ? 1'h0 : dirty_1_3; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_714 = 4'h4 == index ? 1'h0 : dirty_1_4; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_715 = 4'h5 == index ? 1'h0 : dirty_1_5; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_716 = 4'h6 == index ? 1'h0 : dirty_1_6; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_717 = 4'h7 == index ? 1'h0 : dirty_1_7; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_718 = 4'h8 == index ? 1'h0 : dirty_1_8; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_719 = 4'h9 == index ? 1'h0 : dirty_1_9; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_720 = 4'ha == index ? 1'h0 : dirty_1_10; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_721 = 4'hb == index ? 1'h0 : dirty_1_11; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_722 = 4'hc == index ? 1'h0 : dirty_1_12; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_723 = 4'hd == index ? 1'h0 : dirty_1_13; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_724 = 4'he == index ? 1'h0 : dirty_1_14; // @[d_cache.scala 163:{40,40} 27:26]
  wire  _GEN_725 = 4'hf == index ? 1'h0 : dirty_1_15; // @[d_cache.scala 163:{40,40} 27:26]
  wire [127:0] _GEN_822 = _GEN_677 ? _GEN_136 : write_back_data; // @[d_cache.scala 158:47 159:41 31:34]
  wire [39:0] _GEN_823 = _GEN_677 ? _write_back_addr_T_3 : {{8'd0}, write_back_addr}; // @[d_cache.scala 158:47 160:41 32:34]
  wire [127:0] _GEN_824 = _GEN_677 ? _GEN_355 : _GEN_355; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_825 = _GEN_677 ? _GEN_356 : _GEN_356; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_826 = _GEN_677 ? _GEN_357 : _GEN_357; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_827 = _GEN_677 ? _GEN_358 : _GEN_358; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_828 = _GEN_677 ? _GEN_359 : _GEN_359; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_829 = _GEN_677 ? _GEN_360 : _GEN_360; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_830 = _GEN_677 ? _GEN_361 : _GEN_361; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_831 = _GEN_677 ? _GEN_362 : _GEN_362; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_832 = _GEN_677 ? _GEN_363 : _GEN_363; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_833 = _GEN_677 ? _GEN_364 : _GEN_364; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_834 = _GEN_677 ? _GEN_365 : _GEN_365; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_835 = _GEN_677 ? _GEN_366 : _GEN_366; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_836 = _GEN_677 ? _GEN_367 : _GEN_367; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_837 = _GEN_677 ? _GEN_368 : _GEN_368; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_838 = _GEN_677 ? _GEN_369 : _GEN_369; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_839 = _GEN_677 ? _GEN_370 : _GEN_370; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_840 = _GEN_677 ? _GEN_371 : _GEN_371; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_841 = _GEN_677 ? _GEN_372 : _GEN_372; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_842 = _GEN_677 ? _GEN_373 : _GEN_373; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_843 = _GEN_677 ? _GEN_374 : _GEN_374; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_844 = _GEN_677 ? _GEN_375 : _GEN_375; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_845 = _GEN_677 ? _GEN_376 : _GEN_376; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_846 = _GEN_677 ? _GEN_377 : _GEN_377; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_847 = _GEN_677 ? _GEN_378 : _GEN_378; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_848 = _GEN_677 ? _GEN_379 : _GEN_379; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_849 = _GEN_677 ? _GEN_380 : _GEN_380; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_850 = _GEN_677 ? _GEN_381 : _GEN_381; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_851 = _GEN_677 ? _GEN_382 : _GEN_382; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_852 = _GEN_677 ? _GEN_383 : _GEN_383; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_853 = _GEN_677 ? _GEN_384 : _GEN_384; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_854 = _GEN_677 ? _GEN_385 : _GEN_385; // @[d_cache.scala 158:47]
  wire [31:0] _GEN_855 = _GEN_677 ? _GEN_386 : _GEN_386; // @[d_cache.scala 158:47]
  wire  _GEN_856 = _GEN_677 ? _GEN_710 : dirty_1_0; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_857 = _GEN_677 ? _GEN_711 : dirty_1_1; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_858 = _GEN_677 ? _GEN_712 : dirty_1_2; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_859 = _GEN_677 ? _GEN_713 : dirty_1_3; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_860 = _GEN_677 ? _GEN_714 : dirty_1_4; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_861 = _GEN_677 ? _GEN_715 : dirty_1_5; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_862 = _GEN_677 ? _GEN_716 : dirty_1_6; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_863 = _GEN_677 ? _GEN_717 : dirty_1_7; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_864 = _GEN_677 ? _GEN_718 : dirty_1_8; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_865 = _GEN_677 ? _GEN_719 : dirty_1_9; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_866 = _GEN_677 ? _GEN_720 : dirty_1_10; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_867 = _GEN_677 ? _GEN_721 : dirty_1_11; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_868 = _GEN_677 ? _GEN_722 : dirty_1_12; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_869 = _GEN_677 ? _GEN_723 : dirty_1_13; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_870 = _GEN_677 ? _GEN_724 : dirty_1_14; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_871 = _GEN_677 ? _GEN_725 : dirty_1_15; // @[d_cache.scala 158:47 27:26]
  wire  _GEN_872 = _GEN_677 ? _GEN_387 : _GEN_387; // @[d_cache.scala 158:47]
  wire  _GEN_873 = _GEN_677 ? _GEN_388 : _GEN_388; // @[d_cache.scala 158:47]
  wire  _GEN_874 = _GEN_677 ? _GEN_389 : _GEN_389; // @[d_cache.scala 158:47]
  wire  _GEN_875 = _GEN_677 ? _GEN_390 : _GEN_390; // @[d_cache.scala 158:47]
  wire  _GEN_876 = _GEN_677 ? _GEN_391 : _GEN_391; // @[d_cache.scala 158:47]
  wire  _GEN_877 = _GEN_677 ? _GEN_392 : _GEN_392; // @[d_cache.scala 158:47]
  wire  _GEN_878 = _GEN_677 ? _GEN_393 : _GEN_393; // @[d_cache.scala 158:47]
  wire  _GEN_879 = _GEN_677 ? _GEN_394 : _GEN_394; // @[d_cache.scala 158:47]
  wire  _GEN_880 = _GEN_677 ? _GEN_395 : _GEN_395; // @[d_cache.scala 158:47]
  wire  _GEN_881 = _GEN_677 ? _GEN_396 : _GEN_396; // @[d_cache.scala 158:47]
  wire  _GEN_882 = _GEN_677 ? _GEN_397 : _GEN_397; // @[d_cache.scala 158:47]
  wire  _GEN_883 = _GEN_677 ? _GEN_398 : _GEN_398; // @[d_cache.scala 158:47]
  wire  _GEN_884 = _GEN_677 ? _GEN_399 : _GEN_399; // @[d_cache.scala 158:47]
  wire  _GEN_885 = _GEN_677 ? _GEN_400 : _GEN_400; // @[d_cache.scala 158:47]
  wire  _GEN_886 = _GEN_677 ? _GEN_401 : _GEN_401; // @[d_cache.scala 158:47]
  wire  _GEN_887 = _GEN_677 ? _GEN_402 : _GEN_402; // @[d_cache.scala 158:47]
  wire [3:0] _GEN_888 = _GEN_677 ? 4'h6 : 4'h1; // @[d_cache.scala 158:47 165:31 168:31]
  wire [1:0] _GEN_889 = _GEN_677 ? _GEN_403 : _GEN_403; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_890 = _GEN_677 ? _GEN_404 : _GEN_404; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_891 = _GEN_677 ? _GEN_405 : _GEN_405; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_892 = _GEN_677 ? _GEN_406 : _GEN_406; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_893 = _GEN_677 ? _GEN_407 : _GEN_407; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_894 = _GEN_677 ? _GEN_408 : _GEN_408; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_895 = _GEN_677 ? _GEN_409 : _GEN_409; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_896 = _GEN_677 ? _GEN_410 : _GEN_410; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_897 = _GEN_677 ? _GEN_411 : _GEN_411; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_898 = _GEN_677 ? _GEN_412 : _GEN_412; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_899 = _GEN_677 ? _GEN_413 : _GEN_413; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_900 = _GEN_677 ? _GEN_414 : _GEN_414; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_901 = _GEN_677 ? _GEN_415 : _GEN_415; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_902 = _GEN_677 ? _GEN_416 : _GEN_416; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_903 = _GEN_677 ? _GEN_417 : _GEN_417; // @[d_cache.scala 158:47]
  wire [1:0] _GEN_904 = _GEN_677 ? _GEN_418 : _GEN_418; // @[d_cache.scala 158:47]
  wire [127:0] _GEN_905 = ~_GEN_338[1] ? _GEN_579 : _GEN_822; // @[d_cache.scala 139:44]
  wire [39:0] _GEN_906 = ~_GEN_338[1] ? _GEN_580 : _GEN_823; // @[d_cache.scala 139:44]
  wire [127:0] _GEN_907 = ~_GEN_338[1] ? _GEN_581 : ram_0_0; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_908 = ~_GEN_338[1] ? _GEN_582 : ram_0_1; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_909 = ~_GEN_338[1] ? _GEN_583 : ram_0_2; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_910 = ~_GEN_338[1] ? _GEN_584 : ram_0_3; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_911 = ~_GEN_338[1] ? _GEN_585 : ram_0_4; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_912 = ~_GEN_338[1] ? _GEN_586 : ram_0_5; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_913 = ~_GEN_338[1] ? _GEN_587 : ram_0_6; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_914 = ~_GEN_338[1] ? _GEN_588 : ram_0_7; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_915 = ~_GEN_338[1] ? _GEN_589 : ram_0_8; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_916 = ~_GEN_338[1] ? _GEN_590 : ram_0_9; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_917 = ~_GEN_338[1] ? _GEN_591 : ram_0_10; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_918 = ~_GEN_338[1] ? _GEN_592 : ram_0_11; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_919 = ~_GEN_338[1] ? _GEN_593 : ram_0_12; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_920 = ~_GEN_338[1] ? _GEN_594 : ram_0_13; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_921 = ~_GEN_338[1] ? _GEN_595 : ram_0_14; // @[d_cache.scala 139:44 19:24]
  wire [127:0] _GEN_922 = ~_GEN_338[1] ? _GEN_596 : ram_0_15; // @[d_cache.scala 139:44 19:24]
  wire [31:0] _GEN_923 = ~_GEN_338[1] ? _GEN_597 : tag_0_0; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_924 = ~_GEN_338[1] ? _GEN_598 : tag_0_1; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_925 = ~_GEN_338[1] ? _GEN_599 : tag_0_2; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_926 = ~_GEN_338[1] ? _GEN_600 : tag_0_3; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_927 = ~_GEN_338[1] ? _GEN_601 : tag_0_4; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_928 = ~_GEN_338[1] ? _GEN_602 : tag_0_5; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_929 = ~_GEN_338[1] ? _GEN_603 : tag_0_6; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_930 = ~_GEN_338[1] ? _GEN_604 : tag_0_7; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_931 = ~_GEN_338[1] ? _GEN_605 : tag_0_8; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_932 = ~_GEN_338[1] ? _GEN_606 : tag_0_9; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_933 = ~_GEN_338[1] ? _GEN_607 : tag_0_10; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_934 = ~_GEN_338[1] ? _GEN_608 : tag_0_11; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_935 = ~_GEN_338[1] ? _GEN_609 : tag_0_12; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_936 = ~_GEN_338[1] ? _GEN_610 : tag_0_13; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_937 = ~_GEN_338[1] ? _GEN_611 : tag_0_14; // @[d_cache.scala 139:44 22:24]
  wire [31:0] _GEN_938 = ~_GEN_338[1] ? _GEN_612 : tag_0_15; // @[d_cache.scala 139:44 22:24]
  wire  _GEN_939 = ~_GEN_338[1] ? _GEN_613 : dirty_0_0; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_940 = ~_GEN_338[1] ? _GEN_614 : dirty_0_1; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_941 = ~_GEN_338[1] ? _GEN_615 : dirty_0_2; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_942 = ~_GEN_338[1] ? _GEN_616 : dirty_0_3; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_943 = ~_GEN_338[1] ? _GEN_617 : dirty_0_4; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_944 = ~_GEN_338[1] ? _GEN_618 : dirty_0_5; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_945 = ~_GEN_338[1] ? _GEN_619 : dirty_0_6; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_946 = ~_GEN_338[1] ? _GEN_620 : dirty_0_7; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_947 = ~_GEN_338[1] ? _GEN_621 : dirty_0_8; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_948 = ~_GEN_338[1] ? _GEN_622 : dirty_0_9; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_949 = ~_GEN_338[1] ? _GEN_623 : dirty_0_10; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_950 = ~_GEN_338[1] ? _GEN_624 : dirty_0_11; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_951 = ~_GEN_338[1] ? _GEN_625 : dirty_0_12; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_952 = ~_GEN_338[1] ? _GEN_626 : dirty_0_13; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_953 = ~_GEN_338[1] ? _GEN_627 : dirty_0_14; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_954 = ~_GEN_338[1] ? _GEN_628 : dirty_0_15; // @[d_cache.scala 139:44 26:26]
  wire  _GEN_955 = ~_GEN_338[1] ? _GEN_629 : valid_0_0; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_956 = ~_GEN_338[1] ? _GEN_630 : valid_0_1; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_957 = ~_GEN_338[1] ? _GEN_631 : valid_0_2; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_958 = ~_GEN_338[1] ? _GEN_632 : valid_0_3; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_959 = ~_GEN_338[1] ? _GEN_633 : valid_0_4; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_960 = ~_GEN_338[1] ? _GEN_634 : valid_0_5; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_961 = ~_GEN_338[1] ? _GEN_635 : valid_0_6; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_962 = ~_GEN_338[1] ? _GEN_636 : valid_0_7; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_963 = ~_GEN_338[1] ? _GEN_637 : valid_0_8; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_964 = ~_GEN_338[1] ? _GEN_638 : valid_0_9; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_965 = ~_GEN_338[1] ? _GEN_639 : valid_0_10; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_966 = ~_GEN_338[1] ? _GEN_640 : valid_0_11; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_967 = ~_GEN_338[1] ? _GEN_641 : valid_0_12; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_968 = ~_GEN_338[1] ? _GEN_642 : valid_0_13; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_969 = ~_GEN_338[1] ? _GEN_643 : valid_0_14; // @[d_cache.scala 139:44 24:26]
  wire  _GEN_970 = ~_GEN_338[1] ? _GEN_644 : valid_0_15; // @[d_cache.scala 139:44 24:26]
  wire [3:0] _GEN_971 = ~_GEN_338[1] ? _GEN_645 : _GEN_888; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_972 = ~_GEN_338[1] ? _GEN_646 : _GEN_889; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_973 = ~_GEN_338[1] ? _GEN_647 : _GEN_890; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_974 = ~_GEN_338[1] ? _GEN_648 : _GEN_891; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_975 = ~_GEN_338[1] ? _GEN_649 : _GEN_892; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_976 = ~_GEN_338[1] ? _GEN_650 : _GEN_893; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_977 = ~_GEN_338[1] ? _GEN_651 : _GEN_894; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_978 = ~_GEN_338[1] ? _GEN_652 : _GEN_895; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_979 = ~_GEN_338[1] ? _GEN_653 : _GEN_896; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_980 = ~_GEN_338[1] ? _GEN_654 : _GEN_897; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_981 = ~_GEN_338[1] ? _GEN_655 : _GEN_898; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_982 = ~_GEN_338[1] ? _GEN_656 : _GEN_899; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_983 = ~_GEN_338[1] ? _GEN_657 : _GEN_900; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_984 = ~_GEN_338[1] ? _GEN_658 : _GEN_901; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_985 = ~_GEN_338[1] ? _GEN_659 : _GEN_902; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_986 = ~_GEN_338[1] ? _GEN_660 : _GEN_903; // @[d_cache.scala 139:44]
  wire [1:0] _GEN_987 = ~_GEN_338[1] ? _GEN_661 : _GEN_904; // @[d_cache.scala 139:44]
  wire [127:0] _GEN_988 = ~_GEN_338[1] ? ram_1_0 : _GEN_824; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_989 = ~_GEN_338[1] ? ram_1_1 : _GEN_825; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_990 = ~_GEN_338[1] ? ram_1_2 : _GEN_826; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_991 = ~_GEN_338[1] ? ram_1_3 : _GEN_827; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_992 = ~_GEN_338[1] ? ram_1_4 : _GEN_828; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_993 = ~_GEN_338[1] ? ram_1_5 : _GEN_829; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_994 = ~_GEN_338[1] ? ram_1_6 : _GEN_830; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_995 = ~_GEN_338[1] ? ram_1_7 : _GEN_831; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_996 = ~_GEN_338[1] ? ram_1_8 : _GEN_832; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_997 = ~_GEN_338[1] ? ram_1_9 : _GEN_833; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_998 = ~_GEN_338[1] ? ram_1_10 : _GEN_834; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_999 = ~_GEN_338[1] ? ram_1_11 : _GEN_835; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_1000 = ~_GEN_338[1] ? ram_1_12 : _GEN_836; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_1001 = ~_GEN_338[1] ? ram_1_13 : _GEN_837; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_1002 = ~_GEN_338[1] ? ram_1_14 : _GEN_838; // @[d_cache.scala 139:44 20:24]
  wire [127:0] _GEN_1003 = ~_GEN_338[1] ? ram_1_15 : _GEN_839; // @[d_cache.scala 139:44 20:24]
  wire [31:0] _GEN_1004 = ~_GEN_338[1] ? tag_1_0 : _GEN_840; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1005 = ~_GEN_338[1] ? tag_1_1 : _GEN_841; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1006 = ~_GEN_338[1] ? tag_1_2 : _GEN_842; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1007 = ~_GEN_338[1] ? tag_1_3 : _GEN_843; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1008 = ~_GEN_338[1] ? tag_1_4 : _GEN_844; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1009 = ~_GEN_338[1] ? tag_1_5 : _GEN_845; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1010 = ~_GEN_338[1] ? tag_1_6 : _GEN_846; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1011 = ~_GEN_338[1] ? tag_1_7 : _GEN_847; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1012 = ~_GEN_338[1] ? tag_1_8 : _GEN_848; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1013 = ~_GEN_338[1] ? tag_1_9 : _GEN_849; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1014 = ~_GEN_338[1] ? tag_1_10 : _GEN_850; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1015 = ~_GEN_338[1] ? tag_1_11 : _GEN_851; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1016 = ~_GEN_338[1] ? tag_1_12 : _GEN_852; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1017 = ~_GEN_338[1] ? tag_1_13 : _GEN_853; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1018 = ~_GEN_338[1] ? tag_1_14 : _GEN_854; // @[d_cache.scala 139:44 23:24]
  wire [31:0] _GEN_1019 = ~_GEN_338[1] ? tag_1_15 : _GEN_855; // @[d_cache.scala 139:44 23:24]
  wire  _GEN_1020 = ~_GEN_338[1] ? dirty_1_0 : _GEN_856; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1021 = ~_GEN_338[1] ? dirty_1_1 : _GEN_857; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1022 = ~_GEN_338[1] ? dirty_1_2 : _GEN_858; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1023 = ~_GEN_338[1] ? dirty_1_3 : _GEN_859; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1024 = ~_GEN_338[1] ? dirty_1_4 : _GEN_860; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1025 = ~_GEN_338[1] ? dirty_1_5 : _GEN_861; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1026 = ~_GEN_338[1] ? dirty_1_6 : _GEN_862; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1027 = ~_GEN_338[1] ? dirty_1_7 : _GEN_863; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1028 = ~_GEN_338[1] ? dirty_1_8 : _GEN_864; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1029 = ~_GEN_338[1] ? dirty_1_9 : _GEN_865; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1030 = ~_GEN_338[1] ? dirty_1_10 : _GEN_866; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1031 = ~_GEN_338[1] ? dirty_1_11 : _GEN_867; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1032 = ~_GEN_338[1] ? dirty_1_12 : _GEN_868; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1033 = ~_GEN_338[1] ? dirty_1_13 : _GEN_869; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1034 = ~_GEN_338[1] ? dirty_1_14 : _GEN_870; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1035 = ~_GEN_338[1] ? dirty_1_15 : _GEN_871; // @[d_cache.scala 139:44 27:26]
  wire  _GEN_1036 = ~_GEN_338[1] ? valid_1_0 : _GEN_872; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1037 = ~_GEN_338[1] ? valid_1_1 : _GEN_873; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1038 = ~_GEN_338[1] ? valid_1_2 : _GEN_874; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1039 = ~_GEN_338[1] ? valid_1_3 : _GEN_875; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1040 = ~_GEN_338[1] ? valid_1_4 : _GEN_876; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1041 = ~_GEN_338[1] ? valid_1_5 : _GEN_877; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1042 = ~_GEN_338[1] ? valid_1_6 : _GEN_878; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1043 = ~_GEN_338[1] ? valid_1_7 : _GEN_879; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1044 = ~_GEN_338[1] ? valid_1_8 : _GEN_880; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1045 = ~_GEN_338[1] ? valid_1_9 : _GEN_881; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1046 = ~_GEN_338[1] ? valid_1_10 : _GEN_882; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1047 = ~_GEN_338[1] ? valid_1_11 : _GEN_883; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1048 = ~_GEN_338[1] ? valid_1_12 : _GEN_884; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1049 = ~_GEN_338[1] ? valid_1_13 : _GEN_885; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1050 = ~_GEN_338[1] ? valid_1_14 : _GEN_886; // @[d_cache.scala 139:44 25:26]
  wire  _GEN_1051 = ~_GEN_338[1] ? valid_1_15 : _GEN_887; // @[d_cache.scala 139:44 25:26]
  wire [3:0] _GEN_1052 = unuse_way == 2'h2 ? 4'h1 : _GEN_971; // @[d_cache.scala 132:40 133:23]
  wire [127:0] _GEN_1053 = unuse_way == 2'h2 ? _GEN_355 : _GEN_988; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1054 = unuse_way == 2'h2 ? _GEN_356 : _GEN_989; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1055 = unuse_way == 2'h2 ? _GEN_357 : _GEN_990; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1056 = unuse_way == 2'h2 ? _GEN_358 : _GEN_991; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1057 = unuse_way == 2'h2 ? _GEN_359 : _GEN_992; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1058 = unuse_way == 2'h2 ? _GEN_360 : _GEN_993; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1059 = unuse_way == 2'h2 ? _GEN_361 : _GEN_994; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1060 = unuse_way == 2'h2 ? _GEN_362 : _GEN_995; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1061 = unuse_way == 2'h2 ? _GEN_363 : _GEN_996; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1062 = unuse_way == 2'h2 ? _GEN_364 : _GEN_997; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1063 = unuse_way == 2'h2 ? _GEN_365 : _GEN_998; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1064 = unuse_way == 2'h2 ? _GEN_366 : _GEN_999; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1065 = unuse_way == 2'h2 ? _GEN_367 : _GEN_1000; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1066 = unuse_way == 2'h2 ? _GEN_368 : _GEN_1001; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1067 = unuse_way == 2'h2 ? _GEN_369 : _GEN_1002; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1068 = unuse_way == 2'h2 ? _GEN_370 : _GEN_1003; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1069 = unuse_way == 2'h2 ? _GEN_371 : _GEN_1004; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1070 = unuse_way == 2'h2 ? _GEN_372 : _GEN_1005; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1071 = unuse_way == 2'h2 ? _GEN_373 : _GEN_1006; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1072 = unuse_way == 2'h2 ? _GEN_374 : _GEN_1007; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1073 = unuse_way == 2'h2 ? _GEN_375 : _GEN_1008; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1074 = unuse_way == 2'h2 ? _GEN_376 : _GEN_1009; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1075 = unuse_way == 2'h2 ? _GEN_377 : _GEN_1010; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1076 = unuse_way == 2'h2 ? _GEN_378 : _GEN_1011; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1077 = unuse_way == 2'h2 ? _GEN_379 : _GEN_1012; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1078 = unuse_way == 2'h2 ? _GEN_380 : _GEN_1013; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1079 = unuse_way == 2'h2 ? _GEN_381 : _GEN_1014; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1080 = unuse_way == 2'h2 ? _GEN_382 : _GEN_1015; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1081 = unuse_way == 2'h2 ? _GEN_383 : _GEN_1016; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1082 = unuse_way == 2'h2 ? _GEN_384 : _GEN_1017; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1083 = unuse_way == 2'h2 ? _GEN_385 : _GEN_1018; // @[d_cache.scala 132:40]
  wire [31:0] _GEN_1084 = unuse_way == 2'h2 ? _GEN_386 : _GEN_1019; // @[d_cache.scala 132:40]
  wire  _GEN_1085 = unuse_way == 2'h2 ? _GEN_387 : _GEN_1036; // @[d_cache.scala 132:40]
  wire  _GEN_1086 = unuse_way == 2'h2 ? _GEN_388 : _GEN_1037; // @[d_cache.scala 132:40]
  wire  _GEN_1087 = unuse_way == 2'h2 ? _GEN_389 : _GEN_1038; // @[d_cache.scala 132:40]
  wire  _GEN_1088 = unuse_way == 2'h2 ? _GEN_390 : _GEN_1039; // @[d_cache.scala 132:40]
  wire  _GEN_1089 = unuse_way == 2'h2 ? _GEN_391 : _GEN_1040; // @[d_cache.scala 132:40]
  wire  _GEN_1090 = unuse_way == 2'h2 ? _GEN_392 : _GEN_1041; // @[d_cache.scala 132:40]
  wire  _GEN_1091 = unuse_way == 2'h2 ? _GEN_393 : _GEN_1042; // @[d_cache.scala 132:40]
  wire  _GEN_1092 = unuse_way == 2'h2 ? _GEN_394 : _GEN_1043; // @[d_cache.scala 132:40]
  wire  _GEN_1093 = unuse_way == 2'h2 ? _GEN_395 : _GEN_1044; // @[d_cache.scala 132:40]
  wire  _GEN_1094 = unuse_way == 2'h2 ? _GEN_396 : _GEN_1045; // @[d_cache.scala 132:40]
  wire  _GEN_1095 = unuse_way == 2'h2 ? _GEN_397 : _GEN_1046; // @[d_cache.scala 132:40]
  wire  _GEN_1096 = unuse_way == 2'h2 ? _GEN_398 : _GEN_1047; // @[d_cache.scala 132:40]
  wire  _GEN_1097 = unuse_way == 2'h2 ? _GEN_399 : _GEN_1048; // @[d_cache.scala 132:40]
  wire  _GEN_1098 = unuse_way == 2'h2 ? _GEN_400 : _GEN_1049; // @[d_cache.scala 132:40]
  wire  _GEN_1099 = unuse_way == 2'h2 ? _GEN_401 : _GEN_1050; // @[d_cache.scala 132:40]
  wire  _GEN_1100 = unuse_way == 2'h2 ? _GEN_402 : _GEN_1051; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1101 = unuse_way == 2'h2 ? _GEN_403 : _GEN_972; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1102 = unuse_way == 2'h2 ? _GEN_404 : _GEN_973; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1103 = unuse_way == 2'h2 ? _GEN_405 : _GEN_974; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1104 = unuse_way == 2'h2 ? _GEN_406 : _GEN_975; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1105 = unuse_way == 2'h2 ? _GEN_407 : _GEN_976; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1106 = unuse_way == 2'h2 ? _GEN_408 : _GEN_977; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1107 = unuse_way == 2'h2 ? _GEN_409 : _GEN_978; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1108 = unuse_way == 2'h2 ? _GEN_410 : _GEN_979; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1109 = unuse_way == 2'h2 ? _GEN_411 : _GEN_980; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1110 = unuse_way == 2'h2 ? _GEN_412 : _GEN_981; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1111 = unuse_way == 2'h2 ? _GEN_413 : _GEN_982; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1112 = unuse_way == 2'h2 ? _GEN_414 : _GEN_983; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1113 = unuse_way == 2'h2 ? _GEN_415 : _GEN_984; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1114 = unuse_way == 2'h2 ? _GEN_416 : _GEN_985; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1115 = unuse_way == 2'h2 ? _GEN_417 : _GEN_986; // @[d_cache.scala 132:40]
  wire [1:0] _GEN_1116 = unuse_way == 2'h2 ? _GEN_418 : _GEN_987; // @[d_cache.scala 132:40]
  wire [127:0] _GEN_1117 = unuse_way == 2'h2 ? write_back_data : _GEN_905; // @[d_cache.scala 132:40 31:34]
  wire [39:0] _GEN_1118 = unuse_way == 2'h2 ? {{8'd0}, write_back_addr} : _GEN_906; // @[d_cache.scala 132:40 32:34]
  wire [127:0] _GEN_1119 = unuse_way == 2'h2 ? ram_0_0 : _GEN_907; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1120 = unuse_way == 2'h2 ? ram_0_1 : _GEN_908; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1121 = unuse_way == 2'h2 ? ram_0_2 : _GEN_909; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1122 = unuse_way == 2'h2 ? ram_0_3 : _GEN_910; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1123 = unuse_way == 2'h2 ? ram_0_4 : _GEN_911; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1124 = unuse_way == 2'h2 ? ram_0_5 : _GEN_912; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1125 = unuse_way == 2'h2 ? ram_0_6 : _GEN_913; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1126 = unuse_way == 2'h2 ? ram_0_7 : _GEN_914; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1127 = unuse_way == 2'h2 ? ram_0_8 : _GEN_915; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1128 = unuse_way == 2'h2 ? ram_0_9 : _GEN_916; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1129 = unuse_way == 2'h2 ? ram_0_10 : _GEN_917; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1130 = unuse_way == 2'h2 ? ram_0_11 : _GEN_918; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1131 = unuse_way == 2'h2 ? ram_0_12 : _GEN_919; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1132 = unuse_way == 2'h2 ? ram_0_13 : _GEN_920; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1133 = unuse_way == 2'h2 ? ram_0_14 : _GEN_921; // @[d_cache.scala 132:40 19:24]
  wire [127:0] _GEN_1134 = unuse_way == 2'h2 ? ram_0_15 : _GEN_922; // @[d_cache.scala 132:40 19:24]
  wire [31:0] _GEN_1135 = unuse_way == 2'h2 ? tag_0_0 : _GEN_923; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1136 = unuse_way == 2'h2 ? tag_0_1 : _GEN_924; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1137 = unuse_way == 2'h2 ? tag_0_2 : _GEN_925; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1138 = unuse_way == 2'h2 ? tag_0_3 : _GEN_926; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1139 = unuse_way == 2'h2 ? tag_0_4 : _GEN_927; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1140 = unuse_way == 2'h2 ? tag_0_5 : _GEN_928; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1141 = unuse_way == 2'h2 ? tag_0_6 : _GEN_929; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1142 = unuse_way == 2'h2 ? tag_0_7 : _GEN_930; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1143 = unuse_way == 2'h2 ? tag_0_8 : _GEN_931; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1144 = unuse_way == 2'h2 ? tag_0_9 : _GEN_932; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1145 = unuse_way == 2'h2 ? tag_0_10 : _GEN_933; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1146 = unuse_way == 2'h2 ? tag_0_11 : _GEN_934; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1147 = unuse_way == 2'h2 ? tag_0_12 : _GEN_935; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1148 = unuse_way == 2'h2 ? tag_0_13 : _GEN_936; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1149 = unuse_way == 2'h2 ? tag_0_14 : _GEN_937; // @[d_cache.scala 132:40 22:24]
  wire [31:0] _GEN_1150 = unuse_way == 2'h2 ? tag_0_15 : _GEN_938; // @[d_cache.scala 132:40 22:24]
  wire  _GEN_1151 = unuse_way == 2'h2 ? dirty_0_0 : _GEN_939; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1152 = unuse_way == 2'h2 ? dirty_0_1 : _GEN_940; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1153 = unuse_way == 2'h2 ? dirty_0_2 : _GEN_941; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1154 = unuse_way == 2'h2 ? dirty_0_3 : _GEN_942; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1155 = unuse_way == 2'h2 ? dirty_0_4 : _GEN_943; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1156 = unuse_way == 2'h2 ? dirty_0_5 : _GEN_944; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1157 = unuse_way == 2'h2 ? dirty_0_6 : _GEN_945; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1158 = unuse_way == 2'h2 ? dirty_0_7 : _GEN_946; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1159 = unuse_way == 2'h2 ? dirty_0_8 : _GEN_947; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1160 = unuse_way == 2'h2 ? dirty_0_9 : _GEN_948; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1161 = unuse_way == 2'h2 ? dirty_0_10 : _GEN_949; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1162 = unuse_way == 2'h2 ? dirty_0_11 : _GEN_950; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1163 = unuse_way == 2'h2 ? dirty_0_12 : _GEN_951; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1164 = unuse_way == 2'h2 ? dirty_0_13 : _GEN_952; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1165 = unuse_way == 2'h2 ? dirty_0_14 : _GEN_953; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1166 = unuse_way == 2'h2 ? dirty_0_15 : _GEN_954; // @[d_cache.scala 132:40 26:26]
  wire  _GEN_1167 = unuse_way == 2'h2 ? valid_0_0 : _GEN_955; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1168 = unuse_way == 2'h2 ? valid_0_1 : _GEN_956; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1169 = unuse_way == 2'h2 ? valid_0_2 : _GEN_957; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1170 = unuse_way == 2'h2 ? valid_0_3 : _GEN_958; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1171 = unuse_way == 2'h2 ? valid_0_4 : _GEN_959; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1172 = unuse_way == 2'h2 ? valid_0_5 : _GEN_960; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1173 = unuse_way == 2'h2 ? valid_0_6 : _GEN_961; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1174 = unuse_way == 2'h2 ? valid_0_7 : _GEN_962; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1175 = unuse_way == 2'h2 ? valid_0_8 : _GEN_963; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1176 = unuse_way == 2'h2 ? valid_0_9 : _GEN_964; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1177 = unuse_way == 2'h2 ? valid_0_10 : _GEN_965; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1178 = unuse_way == 2'h2 ? valid_0_11 : _GEN_966; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1179 = unuse_way == 2'h2 ? valid_0_12 : _GEN_967; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1180 = unuse_way == 2'h2 ? valid_0_13 : _GEN_968; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1181 = unuse_way == 2'h2 ? valid_0_14 : _GEN_969; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1182 = unuse_way == 2'h2 ? valid_0_15 : _GEN_970; // @[d_cache.scala 132:40 24:26]
  wire  _GEN_1183 = unuse_way == 2'h2 ? dirty_1_0 : _GEN_1020; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1184 = unuse_way == 2'h2 ? dirty_1_1 : _GEN_1021; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1185 = unuse_way == 2'h2 ? dirty_1_2 : _GEN_1022; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1186 = unuse_way == 2'h2 ? dirty_1_3 : _GEN_1023; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1187 = unuse_way == 2'h2 ? dirty_1_4 : _GEN_1024; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1188 = unuse_way == 2'h2 ? dirty_1_5 : _GEN_1025; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1189 = unuse_way == 2'h2 ? dirty_1_6 : _GEN_1026; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1190 = unuse_way == 2'h2 ? dirty_1_7 : _GEN_1027; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1191 = unuse_way == 2'h2 ? dirty_1_8 : _GEN_1028; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1192 = unuse_way == 2'h2 ? dirty_1_9 : _GEN_1029; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1193 = unuse_way == 2'h2 ? dirty_1_10 : _GEN_1030; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1194 = unuse_way == 2'h2 ? dirty_1_11 : _GEN_1031; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1195 = unuse_way == 2'h2 ? dirty_1_12 : _GEN_1032; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1196 = unuse_way == 2'h2 ? dirty_1_13 : _GEN_1033; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1197 = unuse_way == 2'h2 ? dirty_1_14 : _GEN_1034; // @[d_cache.scala 132:40 27:26]
  wire  _GEN_1198 = unuse_way == 2'h2 ? dirty_1_15 : _GEN_1035; // @[d_cache.scala 132:40 27:26]
  wire [3:0] _GEN_1199 = unuse_way == 2'h1 ? 4'h1 : _GEN_1052; // @[d_cache.scala 126:34 127:23]
  wire [127:0] _GEN_1200 = unuse_way == 2'h1 ? _GEN_275 : _GEN_1119; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1201 = unuse_way == 2'h1 ? _GEN_276 : _GEN_1120; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1202 = unuse_way == 2'h1 ? _GEN_277 : _GEN_1121; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1203 = unuse_way == 2'h1 ? _GEN_278 : _GEN_1122; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1204 = unuse_way == 2'h1 ? _GEN_279 : _GEN_1123; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1205 = unuse_way == 2'h1 ? _GEN_280 : _GEN_1124; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1206 = unuse_way == 2'h1 ? _GEN_281 : _GEN_1125; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1207 = unuse_way == 2'h1 ? _GEN_282 : _GEN_1126; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1208 = unuse_way == 2'h1 ? _GEN_283 : _GEN_1127; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1209 = unuse_way == 2'h1 ? _GEN_284 : _GEN_1128; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1210 = unuse_way == 2'h1 ? _GEN_285 : _GEN_1129; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1211 = unuse_way == 2'h1 ? _GEN_286 : _GEN_1130; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1212 = unuse_way == 2'h1 ? _GEN_287 : _GEN_1131; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1213 = unuse_way == 2'h1 ? _GEN_288 : _GEN_1132; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1214 = unuse_way == 2'h1 ? _GEN_289 : _GEN_1133; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1215 = unuse_way == 2'h1 ? _GEN_290 : _GEN_1134; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1216 = unuse_way == 2'h1 ? _GEN_291 : _GEN_1135; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1217 = unuse_way == 2'h1 ? _GEN_292 : _GEN_1136; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1218 = unuse_way == 2'h1 ? _GEN_293 : _GEN_1137; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1219 = unuse_way == 2'h1 ? _GEN_294 : _GEN_1138; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1220 = unuse_way == 2'h1 ? _GEN_295 : _GEN_1139; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1221 = unuse_way == 2'h1 ? _GEN_296 : _GEN_1140; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1222 = unuse_way == 2'h1 ? _GEN_297 : _GEN_1141; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1223 = unuse_way == 2'h1 ? _GEN_298 : _GEN_1142; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1224 = unuse_way == 2'h1 ? _GEN_299 : _GEN_1143; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1225 = unuse_way == 2'h1 ? _GEN_300 : _GEN_1144; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1226 = unuse_way == 2'h1 ? _GEN_301 : _GEN_1145; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1227 = unuse_way == 2'h1 ? _GEN_302 : _GEN_1146; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1228 = unuse_way == 2'h1 ? _GEN_303 : _GEN_1147; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1229 = unuse_way == 2'h1 ? _GEN_304 : _GEN_1148; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1230 = unuse_way == 2'h1 ? _GEN_305 : _GEN_1149; // @[d_cache.scala 126:34]
  wire [31:0] _GEN_1231 = unuse_way == 2'h1 ? _GEN_306 : _GEN_1150; // @[d_cache.scala 126:34]
  wire  _GEN_1232 = unuse_way == 2'h1 ? _GEN_307 : _GEN_1167; // @[d_cache.scala 126:34]
  wire  _GEN_1233 = unuse_way == 2'h1 ? _GEN_308 : _GEN_1168; // @[d_cache.scala 126:34]
  wire  _GEN_1234 = unuse_way == 2'h1 ? _GEN_309 : _GEN_1169; // @[d_cache.scala 126:34]
  wire  _GEN_1235 = unuse_way == 2'h1 ? _GEN_310 : _GEN_1170; // @[d_cache.scala 126:34]
  wire  _GEN_1236 = unuse_way == 2'h1 ? _GEN_311 : _GEN_1171; // @[d_cache.scala 126:34]
  wire  _GEN_1237 = unuse_way == 2'h1 ? _GEN_312 : _GEN_1172; // @[d_cache.scala 126:34]
  wire  _GEN_1238 = unuse_way == 2'h1 ? _GEN_313 : _GEN_1173; // @[d_cache.scala 126:34]
  wire  _GEN_1239 = unuse_way == 2'h1 ? _GEN_314 : _GEN_1174; // @[d_cache.scala 126:34]
  wire  _GEN_1240 = unuse_way == 2'h1 ? _GEN_315 : _GEN_1175; // @[d_cache.scala 126:34]
  wire  _GEN_1241 = unuse_way == 2'h1 ? _GEN_316 : _GEN_1176; // @[d_cache.scala 126:34]
  wire  _GEN_1242 = unuse_way == 2'h1 ? _GEN_317 : _GEN_1177; // @[d_cache.scala 126:34]
  wire  _GEN_1243 = unuse_way == 2'h1 ? _GEN_318 : _GEN_1178; // @[d_cache.scala 126:34]
  wire  _GEN_1244 = unuse_way == 2'h1 ? _GEN_319 : _GEN_1179; // @[d_cache.scala 126:34]
  wire  _GEN_1245 = unuse_way == 2'h1 ? _GEN_320 : _GEN_1180; // @[d_cache.scala 126:34]
  wire  _GEN_1246 = unuse_way == 2'h1 ? _GEN_321 : _GEN_1181; // @[d_cache.scala 126:34]
  wire  _GEN_1247 = unuse_way == 2'h1 ? _GEN_322 : _GEN_1182; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1248 = unuse_way == 2'h1 ? _GEN_339 : _GEN_1101; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1249 = unuse_way == 2'h1 ? _GEN_340 : _GEN_1102; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1250 = unuse_way == 2'h1 ? _GEN_341 : _GEN_1103; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1251 = unuse_way == 2'h1 ? _GEN_342 : _GEN_1104; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1252 = unuse_way == 2'h1 ? _GEN_343 : _GEN_1105; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1253 = unuse_way == 2'h1 ? _GEN_344 : _GEN_1106; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1254 = unuse_way == 2'h1 ? _GEN_345 : _GEN_1107; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1255 = unuse_way == 2'h1 ? _GEN_346 : _GEN_1108; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1256 = unuse_way == 2'h1 ? _GEN_347 : _GEN_1109; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1257 = unuse_way == 2'h1 ? _GEN_348 : _GEN_1110; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1258 = unuse_way == 2'h1 ? _GEN_349 : _GEN_1111; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1259 = unuse_way == 2'h1 ? _GEN_350 : _GEN_1112; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1260 = unuse_way == 2'h1 ? _GEN_351 : _GEN_1113; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1261 = unuse_way == 2'h1 ? _GEN_352 : _GEN_1114; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1262 = unuse_way == 2'h1 ? _GEN_353 : _GEN_1115; // @[d_cache.scala 126:34]
  wire [1:0] _GEN_1263 = unuse_way == 2'h1 ? _GEN_354 : _GEN_1116; // @[d_cache.scala 126:34]
  wire [127:0] _GEN_1264 = unuse_way == 2'h1 ? ram_1_0 : _GEN_1053; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1265 = unuse_way == 2'h1 ? ram_1_1 : _GEN_1054; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1266 = unuse_way == 2'h1 ? ram_1_2 : _GEN_1055; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1267 = unuse_way == 2'h1 ? ram_1_3 : _GEN_1056; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1268 = unuse_way == 2'h1 ? ram_1_4 : _GEN_1057; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1269 = unuse_way == 2'h1 ? ram_1_5 : _GEN_1058; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1270 = unuse_way == 2'h1 ? ram_1_6 : _GEN_1059; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1271 = unuse_way == 2'h1 ? ram_1_7 : _GEN_1060; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1272 = unuse_way == 2'h1 ? ram_1_8 : _GEN_1061; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1273 = unuse_way == 2'h1 ? ram_1_9 : _GEN_1062; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1274 = unuse_way == 2'h1 ? ram_1_10 : _GEN_1063; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1275 = unuse_way == 2'h1 ? ram_1_11 : _GEN_1064; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1276 = unuse_way == 2'h1 ? ram_1_12 : _GEN_1065; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1277 = unuse_way == 2'h1 ? ram_1_13 : _GEN_1066; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1278 = unuse_way == 2'h1 ? ram_1_14 : _GEN_1067; // @[d_cache.scala 126:34 20:24]
  wire [127:0] _GEN_1279 = unuse_way == 2'h1 ? ram_1_15 : _GEN_1068; // @[d_cache.scala 126:34 20:24]
  wire [31:0] _GEN_1280 = unuse_way == 2'h1 ? tag_1_0 : _GEN_1069; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1281 = unuse_way == 2'h1 ? tag_1_1 : _GEN_1070; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1282 = unuse_way == 2'h1 ? tag_1_2 : _GEN_1071; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1283 = unuse_way == 2'h1 ? tag_1_3 : _GEN_1072; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1284 = unuse_way == 2'h1 ? tag_1_4 : _GEN_1073; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1285 = unuse_way == 2'h1 ? tag_1_5 : _GEN_1074; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1286 = unuse_way == 2'h1 ? tag_1_6 : _GEN_1075; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1287 = unuse_way == 2'h1 ? tag_1_7 : _GEN_1076; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1288 = unuse_way == 2'h1 ? tag_1_8 : _GEN_1077; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1289 = unuse_way == 2'h1 ? tag_1_9 : _GEN_1078; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1290 = unuse_way == 2'h1 ? tag_1_10 : _GEN_1079; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1291 = unuse_way == 2'h1 ? tag_1_11 : _GEN_1080; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1292 = unuse_way == 2'h1 ? tag_1_12 : _GEN_1081; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1293 = unuse_way == 2'h1 ? tag_1_13 : _GEN_1082; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1294 = unuse_way == 2'h1 ? tag_1_14 : _GEN_1083; // @[d_cache.scala 126:34 23:24]
  wire [31:0] _GEN_1295 = unuse_way == 2'h1 ? tag_1_15 : _GEN_1084; // @[d_cache.scala 126:34 23:24]
  wire  _GEN_1296 = unuse_way == 2'h1 ? valid_1_0 : _GEN_1085; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1297 = unuse_way == 2'h1 ? valid_1_1 : _GEN_1086; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1298 = unuse_way == 2'h1 ? valid_1_2 : _GEN_1087; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1299 = unuse_way == 2'h1 ? valid_1_3 : _GEN_1088; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1300 = unuse_way == 2'h1 ? valid_1_4 : _GEN_1089; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1301 = unuse_way == 2'h1 ? valid_1_5 : _GEN_1090; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1302 = unuse_way == 2'h1 ? valid_1_6 : _GEN_1091; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1303 = unuse_way == 2'h1 ? valid_1_7 : _GEN_1092; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1304 = unuse_way == 2'h1 ? valid_1_8 : _GEN_1093; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1305 = unuse_way == 2'h1 ? valid_1_9 : _GEN_1094; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1306 = unuse_way == 2'h1 ? valid_1_10 : _GEN_1095; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1307 = unuse_way == 2'h1 ? valid_1_11 : _GEN_1096; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1308 = unuse_way == 2'h1 ? valid_1_12 : _GEN_1097; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1309 = unuse_way == 2'h1 ? valid_1_13 : _GEN_1098; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1310 = unuse_way == 2'h1 ? valid_1_14 : _GEN_1099; // @[d_cache.scala 126:34 25:26]
  wire  _GEN_1311 = unuse_way == 2'h1 ? valid_1_15 : _GEN_1100; // @[d_cache.scala 126:34 25:26]
  wire [127:0] _GEN_1312 = unuse_way == 2'h1 ? write_back_data : _GEN_1117; // @[d_cache.scala 126:34 31:34]
  wire [39:0] _GEN_1313 = unuse_way == 2'h1 ? {{8'd0}, write_back_addr} : _GEN_1118; // @[d_cache.scala 126:34 32:34]
  wire  _GEN_1314 = unuse_way == 2'h1 ? dirty_0_0 : _GEN_1151; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1315 = unuse_way == 2'h1 ? dirty_0_1 : _GEN_1152; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1316 = unuse_way == 2'h1 ? dirty_0_2 : _GEN_1153; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1317 = unuse_way == 2'h1 ? dirty_0_3 : _GEN_1154; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1318 = unuse_way == 2'h1 ? dirty_0_4 : _GEN_1155; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1319 = unuse_way == 2'h1 ? dirty_0_5 : _GEN_1156; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1320 = unuse_way == 2'h1 ? dirty_0_6 : _GEN_1157; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1321 = unuse_way == 2'h1 ? dirty_0_7 : _GEN_1158; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1322 = unuse_way == 2'h1 ? dirty_0_8 : _GEN_1159; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1323 = unuse_way == 2'h1 ? dirty_0_9 : _GEN_1160; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1324 = unuse_way == 2'h1 ? dirty_0_10 : _GEN_1161; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1325 = unuse_way == 2'h1 ? dirty_0_11 : _GEN_1162; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1326 = unuse_way == 2'h1 ? dirty_0_12 : _GEN_1163; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1327 = unuse_way == 2'h1 ? dirty_0_13 : _GEN_1164; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1328 = unuse_way == 2'h1 ? dirty_0_14 : _GEN_1165; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1329 = unuse_way == 2'h1 ? dirty_0_15 : _GEN_1166; // @[d_cache.scala 126:34 26:26]
  wire  _GEN_1330 = unuse_way == 2'h1 ? dirty_1_0 : _GEN_1183; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1331 = unuse_way == 2'h1 ? dirty_1_1 : _GEN_1184; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1332 = unuse_way == 2'h1 ? dirty_1_2 : _GEN_1185; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1333 = unuse_way == 2'h1 ? dirty_1_3 : _GEN_1186; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1334 = unuse_way == 2'h1 ? dirty_1_4 : _GEN_1187; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1335 = unuse_way == 2'h1 ? dirty_1_5 : _GEN_1188; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1336 = unuse_way == 2'h1 ? dirty_1_6 : _GEN_1189; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1337 = unuse_way == 2'h1 ? dirty_1_7 : _GEN_1190; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1338 = unuse_way == 2'h1 ? dirty_1_8 : _GEN_1191; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1339 = unuse_way == 2'h1 ? dirty_1_9 : _GEN_1192; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1340 = unuse_way == 2'h1 ? dirty_1_10 : _GEN_1193; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1341 = unuse_way == 2'h1 ? dirty_1_11 : _GEN_1194; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1342 = unuse_way == 2'h1 ? dirty_1_12 : _GEN_1195; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1343 = unuse_way == 2'h1 ? dirty_1_13 : _GEN_1196; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1344 = unuse_way == 2'h1 ? dirty_1_14 : _GEN_1197; // @[d_cache.scala 126:34 27:26]
  wire  _GEN_1345 = unuse_way == 2'h1 ? dirty_1_15 : _GEN_1198; // @[d_cache.scala 126:34 27:26]
  wire [127:0] _write_back_data_T = {{64'd0}, write_back_data[127:64]}; // @[d_cache.scala 179:52]
  wire [127:0] _GEN_1346 = io_from_axi_wready ? _write_back_data_T : write_back_data; // @[d_cache.scala 178:37 179:33 31:34]
  wire [3:0] _GEN_1347 = io_from_axi_bvalid ? 4'h1 : state; // @[d_cache.scala 181:37 182:23 60:24]
  wire [3:0] _GEN_1348 = io_from_axi_rvalid ? 4'h0 : state; // @[d_cache.scala 186:37 187:23 60:24]
  wire [3:0] _GEN_1350 = 4'h8 == state ? _GEN_274 : state; // @[d_cache.scala 65:18 60:24]
  wire [3:0] _GEN_1351 = 4'h7 == state ? _GEN_1348 : _GEN_1350; // @[d_cache.scala 65:18]
  wire [127:0] _GEN_1352 = 4'h6 == state ? _GEN_1346 : write_back_data; // @[d_cache.scala 65:18 31:34]
  wire [3:0] _GEN_1353 = 4'h6 == state ? _GEN_1347 : _GEN_1351; // @[d_cache.scala 65:18]
  wire [3:0] _GEN_1354 = 4'h5 == state ? _GEN_1199 : _GEN_1353; // @[d_cache.scala 65:18]
  wire [127:0] _GEN_1355 = 4'h5 == state ? _GEN_1200 : ram_0_0; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1356 = 4'h5 == state ? _GEN_1201 : ram_0_1; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1357 = 4'h5 == state ? _GEN_1202 : ram_0_2; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1358 = 4'h5 == state ? _GEN_1203 : ram_0_3; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1359 = 4'h5 == state ? _GEN_1204 : ram_0_4; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1360 = 4'h5 == state ? _GEN_1205 : ram_0_5; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1361 = 4'h5 == state ? _GEN_1206 : ram_0_6; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1362 = 4'h5 == state ? _GEN_1207 : ram_0_7; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1363 = 4'h5 == state ? _GEN_1208 : ram_0_8; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1364 = 4'h5 == state ? _GEN_1209 : ram_0_9; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1365 = 4'h5 == state ? _GEN_1210 : ram_0_10; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1366 = 4'h5 == state ? _GEN_1211 : ram_0_11; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1367 = 4'h5 == state ? _GEN_1212 : ram_0_12; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1368 = 4'h5 == state ? _GEN_1213 : ram_0_13; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1369 = 4'h5 == state ? _GEN_1214 : ram_0_14; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1370 = 4'h5 == state ? _GEN_1215 : ram_0_15; // @[d_cache.scala 65:18 19:24]
  wire [31:0] _GEN_1371 = 4'h5 == state ? _GEN_1216 : tag_0_0; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1372 = 4'h5 == state ? _GEN_1217 : tag_0_1; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1373 = 4'h5 == state ? _GEN_1218 : tag_0_2; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1374 = 4'h5 == state ? _GEN_1219 : tag_0_3; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1375 = 4'h5 == state ? _GEN_1220 : tag_0_4; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1376 = 4'h5 == state ? _GEN_1221 : tag_0_5; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1377 = 4'h5 == state ? _GEN_1222 : tag_0_6; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1378 = 4'h5 == state ? _GEN_1223 : tag_0_7; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1379 = 4'h5 == state ? _GEN_1224 : tag_0_8; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1380 = 4'h5 == state ? _GEN_1225 : tag_0_9; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1381 = 4'h5 == state ? _GEN_1226 : tag_0_10; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1382 = 4'h5 == state ? _GEN_1227 : tag_0_11; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1383 = 4'h5 == state ? _GEN_1228 : tag_0_12; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1384 = 4'h5 == state ? _GEN_1229 : tag_0_13; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1385 = 4'h5 == state ? _GEN_1230 : tag_0_14; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1386 = 4'h5 == state ? _GEN_1231 : tag_0_15; // @[d_cache.scala 65:18 22:24]
  wire  _GEN_1387 = 4'h5 == state ? _GEN_1232 : valid_0_0; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1388 = 4'h5 == state ? _GEN_1233 : valid_0_1; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1389 = 4'h5 == state ? _GEN_1234 : valid_0_2; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1390 = 4'h5 == state ? _GEN_1235 : valid_0_3; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1391 = 4'h5 == state ? _GEN_1236 : valid_0_4; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1392 = 4'h5 == state ? _GEN_1237 : valid_0_5; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1393 = 4'h5 == state ? _GEN_1238 : valid_0_6; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1394 = 4'h5 == state ? _GEN_1239 : valid_0_7; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1395 = 4'h5 == state ? _GEN_1240 : valid_0_8; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1396 = 4'h5 == state ? _GEN_1241 : valid_0_9; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1397 = 4'h5 == state ? _GEN_1242 : valid_0_10; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1398 = 4'h5 == state ? _GEN_1243 : valid_0_11; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1399 = 4'h5 == state ? _GEN_1244 : valid_0_12; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1400 = 4'h5 == state ? _GEN_1245 : valid_0_13; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1401 = 4'h5 == state ? _GEN_1246 : valid_0_14; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1402 = 4'h5 == state ? _GEN_1247 : valid_0_15; // @[d_cache.scala 65:18 24:26]
  wire [1:0] _GEN_1403 = 4'h5 == state ? _GEN_1248 : quene_0; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1404 = 4'h5 == state ? _GEN_1249 : quene_1; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1405 = 4'h5 == state ? _GEN_1250 : quene_2; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1406 = 4'h5 == state ? _GEN_1251 : quene_3; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1407 = 4'h5 == state ? _GEN_1252 : quene_4; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1408 = 4'h5 == state ? _GEN_1253 : quene_5; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1409 = 4'h5 == state ? _GEN_1254 : quene_6; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1410 = 4'h5 == state ? _GEN_1255 : quene_7; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1411 = 4'h5 == state ? _GEN_1256 : quene_8; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1412 = 4'h5 == state ? _GEN_1257 : quene_9; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1413 = 4'h5 == state ? _GEN_1258 : quene_10; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1414 = 4'h5 == state ? _GEN_1259 : quene_11; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1415 = 4'h5 == state ? _GEN_1260 : quene_12; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1416 = 4'h5 == state ? _GEN_1261 : quene_13; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1417 = 4'h5 == state ? _GEN_1262 : quene_14; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1418 = 4'h5 == state ? _GEN_1263 : quene_15; // @[d_cache.scala 65:18 39:24]
  wire [127:0] _GEN_1419 = 4'h5 == state ? _GEN_1264 : ram_1_0; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1420 = 4'h5 == state ? _GEN_1265 : ram_1_1; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1421 = 4'h5 == state ? _GEN_1266 : ram_1_2; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1422 = 4'h5 == state ? _GEN_1267 : ram_1_3; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1423 = 4'h5 == state ? _GEN_1268 : ram_1_4; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1424 = 4'h5 == state ? _GEN_1269 : ram_1_5; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1425 = 4'h5 == state ? _GEN_1270 : ram_1_6; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1426 = 4'h5 == state ? _GEN_1271 : ram_1_7; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1427 = 4'h5 == state ? _GEN_1272 : ram_1_8; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1428 = 4'h5 == state ? _GEN_1273 : ram_1_9; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1429 = 4'h5 == state ? _GEN_1274 : ram_1_10; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1430 = 4'h5 == state ? _GEN_1275 : ram_1_11; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1431 = 4'h5 == state ? _GEN_1276 : ram_1_12; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1432 = 4'h5 == state ? _GEN_1277 : ram_1_13; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1433 = 4'h5 == state ? _GEN_1278 : ram_1_14; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1434 = 4'h5 == state ? _GEN_1279 : ram_1_15; // @[d_cache.scala 65:18 20:24]
  wire [31:0] _GEN_1435 = 4'h5 == state ? _GEN_1280 : tag_1_0; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1436 = 4'h5 == state ? _GEN_1281 : tag_1_1; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1437 = 4'h5 == state ? _GEN_1282 : tag_1_2; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1438 = 4'h5 == state ? _GEN_1283 : tag_1_3; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1439 = 4'h5 == state ? _GEN_1284 : tag_1_4; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1440 = 4'h5 == state ? _GEN_1285 : tag_1_5; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1441 = 4'h5 == state ? _GEN_1286 : tag_1_6; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1442 = 4'h5 == state ? _GEN_1287 : tag_1_7; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1443 = 4'h5 == state ? _GEN_1288 : tag_1_8; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1444 = 4'h5 == state ? _GEN_1289 : tag_1_9; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1445 = 4'h5 == state ? _GEN_1290 : tag_1_10; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1446 = 4'h5 == state ? _GEN_1291 : tag_1_11; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1447 = 4'h5 == state ? _GEN_1292 : tag_1_12; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1448 = 4'h5 == state ? _GEN_1293 : tag_1_13; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1449 = 4'h5 == state ? _GEN_1294 : tag_1_14; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1450 = 4'h5 == state ? _GEN_1295 : tag_1_15; // @[d_cache.scala 65:18 23:24]
  wire  _GEN_1451 = 4'h5 == state ? _GEN_1296 : valid_1_0; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1452 = 4'h5 == state ? _GEN_1297 : valid_1_1; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1453 = 4'h5 == state ? _GEN_1298 : valid_1_2; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1454 = 4'h5 == state ? _GEN_1299 : valid_1_3; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1455 = 4'h5 == state ? _GEN_1300 : valid_1_4; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1456 = 4'h5 == state ? _GEN_1301 : valid_1_5; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1457 = 4'h5 == state ? _GEN_1302 : valid_1_6; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1458 = 4'h5 == state ? _GEN_1303 : valid_1_7; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1459 = 4'h5 == state ? _GEN_1304 : valid_1_8; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1460 = 4'h5 == state ? _GEN_1305 : valid_1_9; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1461 = 4'h5 == state ? _GEN_1306 : valid_1_10; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1462 = 4'h5 == state ? _GEN_1307 : valid_1_11; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1463 = 4'h5 == state ? _GEN_1308 : valid_1_12; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1464 = 4'h5 == state ? _GEN_1309 : valid_1_13; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1465 = 4'h5 == state ? _GEN_1310 : valid_1_14; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1466 = 4'h5 == state ? _GEN_1311 : valid_1_15; // @[d_cache.scala 65:18 25:26]
  wire [127:0] _GEN_1467 = 4'h5 == state ? _GEN_1312 : _GEN_1352; // @[d_cache.scala 65:18]
  wire [39:0] _GEN_1468 = 4'h5 == state ? _GEN_1313 : {{8'd0}, write_back_addr}; // @[d_cache.scala 65:18 32:34]
  wire  _GEN_1469 = 4'h5 == state ? _GEN_1314 : dirty_0_0; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1470 = 4'h5 == state ? _GEN_1315 : dirty_0_1; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1471 = 4'h5 == state ? _GEN_1316 : dirty_0_2; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1472 = 4'h5 == state ? _GEN_1317 : dirty_0_3; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1473 = 4'h5 == state ? _GEN_1318 : dirty_0_4; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1474 = 4'h5 == state ? _GEN_1319 : dirty_0_5; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1475 = 4'h5 == state ? _GEN_1320 : dirty_0_6; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1476 = 4'h5 == state ? _GEN_1321 : dirty_0_7; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1477 = 4'h5 == state ? _GEN_1322 : dirty_0_8; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1478 = 4'h5 == state ? _GEN_1323 : dirty_0_9; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1479 = 4'h5 == state ? _GEN_1324 : dirty_0_10; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1480 = 4'h5 == state ? _GEN_1325 : dirty_0_11; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1481 = 4'h5 == state ? _GEN_1326 : dirty_0_12; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1482 = 4'h5 == state ? _GEN_1327 : dirty_0_13; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1483 = 4'h5 == state ? _GEN_1328 : dirty_0_14; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1484 = 4'h5 == state ? _GEN_1329 : dirty_0_15; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1485 = 4'h5 == state ? _GEN_1330 : dirty_1_0; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1486 = 4'h5 == state ? _GEN_1331 : dirty_1_1; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1487 = 4'h5 == state ? _GEN_1332 : dirty_1_2; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1488 = 4'h5 == state ? _GEN_1333 : dirty_1_3; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1489 = 4'h5 == state ? _GEN_1334 : dirty_1_4; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1490 = 4'h5 == state ? _GEN_1335 : dirty_1_5; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1491 = 4'h5 == state ? _GEN_1336 : dirty_1_6; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1492 = 4'h5 == state ? _GEN_1337 : dirty_1_7; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1493 = 4'h5 == state ? _GEN_1338 : dirty_1_8; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1494 = 4'h5 == state ? _GEN_1339 : dirty_1_9; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1495 = 4'h5 == state ? _GEN_1340 : dirty_1_10; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1496 = 4'h5 == state ? _GEN_1341 : dirty_1_11; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1497 = 4'h5 == state ? _GEN_1342 : dirty_1_12; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1498 = 4'h5 == state ? _GEN_1343 : dirty_1_13; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1499 = 4'h5 == state ? _GEN_1344 : dirty_1_14; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1500 = 4'h5 == state ? _GEN_1345 : dirty_1_15; // @[d_cache.scala 65:18 27:26]
  wire [3:0] _GEN_1501 = 4'h4 == state ? _GEN_274 : _GEN_1354; // @[d_cache.scala 65:18]
  wire [127:0] _GEN_1502 = 4'h4 == state ? ram_0_0 : _GEN_1355; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1503 = 4'h4 == state ? ram_0_1 : _GEN_1356; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1504 = 4'h4 == state ? ram_0_2 : _GEN_1357; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1505 = 4'h4 == state ? ram_0_3 : _GEN_1358; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1506 = 4'h4 == state ? ram_0_4 : _GEN_1359; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1507 = 4'h4 == state ? ram_0_5 : _GEN_1360; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1508 = 4'h4 == state ? ram_0_6 : _GEN_1361; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1509 = 4'h4 == state ? ram_0_7 : _GEN_1362; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1510 = 4'h4 == state ? ram_0_8 : _GEN_1363; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1511 = 4'h4 == state ? ram_0_9 : _GEN_1364; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1512 = 4'h4 == state ? ram_0_10 : _GEN_1365; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1513 = 4'h4 == state ? ram_0_11 : _GEN_1366; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1514 = 4'h4 == state ? ram_0_12 : _GEN_1367; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1515 = 4'h4 == state ? ram_0_13 : _GEN_1368; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1516 = 4'h4 == state ? ram_0_14 : _GEN_1369; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1517 = 4'h4 == state ? ram_0_15 : _GEN_1370; // @[d_cache.scala 65:18 19:24]
  wire [31:0] _GEN_1518 = 4'h4 == state ? tag_0_0 : _GEN_1371; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1519 = 4'h4 == state ? tag_0_1 : _GEN_1372; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1520 = 4'h4 == state ? tag_0_2 : _GEN_1373; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1521 = 4'h4 == state ? tag_0_3 : _GEN_1374; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1522 = 4'h4 == state ? tag_0_4 : _GEN_1375; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1523 = 4'h4 == state ? tag_0_5 : _GEN_1376; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1524 = 4'h4 == state ? tag_0_6 : _GEN_1377; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1525 = 4'h4 == state ? tag_0_7 : _GEN_1378; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1526 = 4'h4 == state ? tag_0_8 : _GEN_1379; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1527 = 4'h4 == state ? tag_0_9 : _GEN_1380; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1528 = 4'h4 == state ? tag_0_10 : _GEN_1381; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1529 = 4'h4 == state ? tag_0_11 : _GEN_1382; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1530 = 4'h4 == state ? tag_0_12 : _GEN_1383; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1531 = 4'h4 == state ? tag_0_13 : _GEN_1384; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1532 = 4'h4 == state ? tag_0_14 : _GEN_1385; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1533 = 4'h4 == state ? tag_0_15 : _GEN_1386; // @[d_cache.scala 65:18 22:24]
  wire  _GEN_1534 = 4'h4 == state ? valid_0_0 : _GEN_1387; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1535 = 4'h4 == state ? valid_0_1 : _GEN_1388; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1536 = 4'h4 == state ? valid_0_2 : _GEN_1389; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1537 = 4'h4 == state ? valid_0_3 : _GEN_1390; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1538 = 4'h4 == state ? valid_0_4 : _GEN_1391; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1539 = 4'h4 == state ? valid_0_5 : _GEN_1392; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1540 = 4'h4 == state ? valid_0_6 : _GEN_1393; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1541 = 4'h4 == state ? valid_0_7 : _GEN_1394; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1542 = 4'h4 == state ? valid_0_8 : _GEN_1395; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1543 = 4'h4 == state ? valid_0_9 : _GEN_1396; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1544 = 4'h4 == state ? valid_0_10 : _GEN_1397; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1545 = 4'h4 == state ? valid_0_11 : _GEN_1398; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1546 = 4'h4 == state ? valid_0_12 : _GEN_1399; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1547 = 4'h4 == state ? valid_0_13 : _GEN_1400; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1548 = 4'h4 == state ? valid_0_14 : _GEN_1401; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1549 = 4'h4 == state ? valid_0_15 : _GEN_1402; // @[d_cache.scala 65:18 24:26]
  wire [1:0] _GEN_1550 = 4'h4 == state ? quene_0 : _GEN_1403; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1551 = 4'h4 == state ? quene_1 : _GEN_1404; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1552 = 4'h4 == state ? quene_2 : _GEN_1405; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1553 = 4'h4 == state ? quene_3 : _GEN_1406; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1554 = 4'h4 == state ? quene_4 : _GEN_1407; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1555 = 4'h4 == state ? quene_5 : _GEN_1408; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1556 = 4'h4 == state ? quene_6 : _GEN_1409; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1557 = 4'h4 == state ? quene_7 : _GEN_1410; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1558 = 4'h4 == state ? quene_8 : _GEN_1411; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1559 = 4'h4 == state ? quene_9 : _GEN_1412; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1560 = 4'h4 == state ? quene_10 : _GEN_1413; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1561 = 4'h4 == state ? quene_11 : _GEN_1414; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1562 = 4'h4 == state ? quene_12 : _GEN_1415; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1563 = 4'h4 == state ? quene_13 : _GEN_1416; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1564 = 4'h4 == state ? quene_14 : _GEN_1417; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1565 = 4'h4 == state ? quene_15 : _GEN_1418; // @[d_cache.scala 65:18 39:24]
  wire [127:0] _GEN_1566 = 4'h4 == state ? ram_1_0 : _GEN_1419; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1567 = 4'h4 == state ? ram_1_1 : _GEN_1420; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1568 = 4'h4 == state ? ram_1_2 : _GEN_1421; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1569 = 4'h4 == state ? ram_1_3 : _GEN_1422; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1570 = 4'h4 == state ? ram_1_4 : _GEN_1423; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1571 = 4'h4 == state ? ram_1_5 : _GEN_1424; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1572 = 4'h4 == state ? ram_1_6 : _GEN_1425; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1573 = 4'h4 == state ? ram_1_7 : _GEN_1426; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1574 = 4'h4 == state ? ram_1_8 : _GEN_1427; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1575 = 4'h4 == state ? ram_1_9 : _GEN_1428; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1576 = 4'h4 == state ? ram_1_10 : _GEN_1429; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1577 = 4'h4 == state ? ram_1_11 : _GEN_1430; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1578 = 4'h4 == state ? ram_1_12 : _GEN_1431; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1579 = 4'h4 == state ? ram_1_13 : _GEN_1432; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1580 = 4'h4 == state ? ram_1_14 : _GEN_1433; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1581 = 4'h4 == state ? ram_1_15 : _GEN_1434; // @[d_cache.scala 65:18 20:24]
  wire [31:0] _GEN_1582 = 4'h4 == state ? tag_1_0 : _GEN_1435; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1583 = 4'h4 == state ? tag_1_1 : _GEN_1436; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1584 = 4'h4 == state ? tag_1_2 : _GEN_1437; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1585 = 4'h4 == state ? tag_1_3 : _GEN_1438; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1586 = 4'h4 == state ? tag_1_4 : _GEN_1439; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1587 = 4'h4 == state ? tag_1_5 : _GEN_1440; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1588 = 4'h4 == state ? tag_1_6 : _GEN_1441; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1589 = 4'h4 == state ? tag_1_7 : _GEN_1442; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1590 = 4'h4 == state ? tag_1_8 : _GEN_1443; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1591 = 4'h4 == state ? tag_1_9 : _GEN_1444; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1592 = 4'h4 == state ? tag_1_10 : _GEN_1445; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1593 = 4'h4 == state ? tag_1_11 : _GEN_1446; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1594 = 4'h4 == state ? tag_1_12 : _GEN_1447; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1595 = 4'h4 == state ? tag_1_13 : _GEN_1448; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1596 = 4'h4 == state ? tag_1_14 : _GEN_1449; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1597 = 4'h4 == state ? tag_1_15 : _GEN_1450; // @[d_cache.scala 65:18 23:24]
  wire  _GEN_1598 = 4'h4 == state ? valid_1_0 : _GEN_1451; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1599 = 4'h4 == state ? valid_1_1 : _GEN_1452; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1600 = 4'h4 == state ? valid_1_2 : _GEN_1453; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1601 = 4'h4 == state ? valid_1_3 : _GEN_1454; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1602 = 4'h4 == state ? valid_1_4 : _GEN_1455; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1603 = 4'h4 == state ? valid_1_5 : _GEN_1456; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1604 = 4'h4 == state ? valid_1_6 : _GEN_1457; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1605 = 4'h4 == state ? valid_1_7 : _GEN_1458; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1606 = 4'h4 == state ? valid_1_8 : _GEN_1459; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1607 = 4'h4 == state ? valid_1_9 : _GEN_1460; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1608 = 4'h4 == state ? valid_1_10 : _GEN_1461; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1609 = 4'h4 == state ? valid_1_11 : _GEN_1462; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1610 = 4'h4 == state ? valid_1_12 : _GEN_1463; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1611 = 4'h4 == state ? valid_1_13 : _GEN_1464; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1612 = 4'h4 == state ? valid_1_14 : _GEN_1465; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1613 = 4'h4 == state ? valid_1_15 : _GEN_1466; // @[d_cache.scala 65:18 25:26]
  wire [127:0] _GEN_1614 = 4'h4 == state ? write_back_data : _GEN_1467; // @[d_cache.scala 65:18 31:34]
  wire [39:0] _GEN_1615 = 4'h4 == state ? {{8'd0}, write_back_addr} : _GEN_1468; // @[d_cache.scala 65:18 32:34]
  wire  _GEN_1616 = 4'h4 == state ? dirty_0_0 : _GEN_1469; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1617 = 4'h4 == state ? dirty_0_1 : _GEN_1470; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1618 = 4'h4 == state ? dirty_0_2 : _GEN_1471; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1619 = 4'h4 == state ? dirty_0_3 : _GEN_1472; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1620 = 4'h4 == state ? dirty_0_4 : _GEN_1473; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1621 = 4'h4 == state ? dirty_0_5 : _GEN_1474; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1622 = 4'h4 == state ? dirty_0_6 : _GEN_1475; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1623 = 4'h4 == state ? dirty_0_7 : _GEN_1476; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1624 = 4'h4 == state ? dirty_0_8 : _GEN_1477; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1625 = 4'h4 == state ? dirty_0_9 : _GEN_1478; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1626 = 4'h4 == state ? dirty_0_10 : _GEN_1479; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1627 = 4'h4 == state ? dirty_0_11 : _GEN_1480; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1628 = 4'h4 == state ? dirty_0_12 : _GEN_1481; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1629 = 4'h4 == state ? dirty_0_13 : _GEN_1482; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1630 = 4'h4 == state ? dirty_0_14 : _GEN_1483; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1631 = 4'h4 == state ? dirty_0_15 : _GEN_1484; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1632 = 4'h4 == state ? dirty_1_0 : _GEN_1485; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1633 = 4'h4 == state ? dirty_1_1 : _GEN_1486; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1634 = 4'h4 == state ? dirty_1_2 : _GEN_1487; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1635 = 4'h4 == state ? dirty_1_3 : _GEN_1488; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1636 = 4'h4 == state ? dirty_1_4 : _GEN_1489; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1637 = 4'h4 == state ? dirty_1_5 : _GEN_1490; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1638 = 4'h4 == state ? dirty_1_6 : _GEN_1491; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1639 = 4'h4 == state ? dirty_1_7 : _GEN_1492; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1640 = 4'h4 == state ? dirty_1_8 : _GEN_1493; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1641 = 4'h4 == state ? dirty_1_9 : _GEN_1494; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1642 = 4'h4 == state ? dirty_1_10 : _GEN_1495; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1643 = 4'h4 == state ? dirty_1_11 : _GEN_1496; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1644 = 4'h4 == state ? dirty_1_12 : _GEN_1497; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1645 = 4'h4 == state ? dirty_1_13 : _GEN_1498; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1646 = 4'h4 == state ? dirty_1_14 : _GEN_1499; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1647 = 4'h4 == state ? dirty_1_15 : _GEN_1500; // @[d_cache.scala 65:18 27:26]
  wire [63:0] _GEN_1648 = 4'h3 == state ? _GEN_270 : receive_data_0; // @[d_cache.scala 65:18 37:31]
  wire [63:0] _GEN_1649 = 4'h3 == state ? _GEN_271 : receive_data_1; // @[d_cache.scala 65:18 37:31]
  wire [2:0] _GEN_1650 = 4'h3 == state ? _GEN_272 : receive_num; // @[d_cache.scala 65:18 38:30]
  wire [3:0] _GEN_1651 = 4'h3 == state ? _GEN_273 : _GEN_1501; // @[d_cache.scala 65:18]
  wire [127:0] _GEN_1652 = 4'h3 == state ? ram_0_0 : _GEN_1502; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1653 = 4'h3 == state ? ram_0_1 : _GEN_1503; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1654 = 4'h3 == state ? ram_0_2 : _GEN_1504; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1655 = 4'h3 == state ? ram_0_3 : _GEN_1505; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1656 = 4'h3 == state ? ram_0_4 : _GEN_1506; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1657 = 4'h3 == state ? ram_0_5 : _GEN_1507; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1658 = 4'h3 == state ? ram_0_6 : _GEN_1508; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1659 = 4'h3 == state ? ram_0_7 : _GEN_1509; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1660 = 4'h3 == state ? ram_0_8 : _GEN_1510; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1661 = 4'h3 == state ? ram_0_9 : _GEN_1511; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1662 = 4'h3 == state ? ram_0_10 : _GEN_1512; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1663 = 4'h3 == state ? ram_0_11 : _GEN_1513; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1664 = 4'h3 == state ? ram_0_12 : _GEN_1514; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1665 = 4'h3 == state ? ram_0_13 : _GEN_1515; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1666 = 4'h3 == state ? ram_0_14 : _GEN_1516; // @[d_cache.scala 65:18 19:24]
  wire [127:0] _GEN_1667 = 4'h3 == state ? ram_0_15 : _GEN_1517; // @[d_cache.scala 65:18 19:24]
  wire [31:0] _GEN_1668 = 4'h3 == state ? tag_0_0 : _GEN_1518; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1669 = 4'h3 == state ? tag_0_1 : _GEN_1519; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1670 = 4'h3 == state ? tag_0_2 : _GEN_1520; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1671 = 4'h3 == state ? tag_0_3 : _GEN_1521; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1672 = 4'h3 == state ? tag_0_4 : _GEN_1522; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1673 = 4'h3 == state ? tag_0_5 : _GEN_1523; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1674 = 4'h3 == state ? tag_0_6 : _GEN_1524; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1675 = 4'h3 == state ? tag_0_7 : _GEN_1525; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1676 = 4'h3 == state ? tag_0_8 : _GEN_1526; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1677 = 4'h3 == state ? tag_0_9 : _GEN_1527; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1678 = 4'h3 == state ? tag_0_10 : _GEN_1528; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1679 = 4'h3 == state ? tag_0_11 : _GEN_1529; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1680 = 4'h3 == state ? tag_0_12 : _GEN_1530; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1681 = 4'h3 == state ? tag_0_13 : _GEN_1531; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1682 = 4'h3 == state ? tag_0_14 : _GEN_1532; // @[d_cache.scala 65:18 22:24]
  wire [31:0] _GEN_1683 = 4'h3 == state ? tag_0_15 : _GEN_1533; // @[d_cache.scala 65:18 22:24]
  wire  _GEN_1684 = 4'h3 == state ? valid_0_0 : _GEN_1534; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1685 = 4'h3 == state ? valid_0_1 : _GEN_1535; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1686 = 4'h3 == state ? valid_0_2 : _GEN_1536; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1687 = 4'h3 == state ? valid_0_3 : _GEN_1537; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1688 = 4'h3 == state ? valid_0_4 : _GEN_1538; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1689 = 4'h3 == state ? valid_0_5 : _GEN_1539; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1690 = 4'h3 == state ? valid_0_6 : _GEN_1540; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1691 = 4'h3 == state ? valid_0_7 : _GEN_1541; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1692 = 4'h3 == state ? valid_0_8 : _GEN_1542; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1693 = 4'h3 == state ? valid_0_9 : _GEN_1543; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1694 = 4'h3 == state ? valid_0_10 : _GEN_1544; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1695 = 4'h3 == state ? valid_0_11 : _GEN_1545; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1696 = 4'h3 == state ? valid_0_12 : _GEN_1546; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1697 = 4'h3 == state ? valid_0_13 : _GEN_1547; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1698 = 4'h3 == state ? valid_0_14 : _GEN_1548; // @[d_cache.scala 65:18 24:26]
  wire  _GEN_1699 = 4'h3 == state ? valid_0_15 : _GEN_1549; // @[d_cache.scala 65:18 24:26]
  wire [1:0] _GEN_1700 = 4'h3 == state ? quene_0 : _GEN_1550; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1701 = 4'h3 == state ? quene_1 : _GEN_1551; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1702 = 4'h3 == state ? quene_2 : _GEN_1552; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1703 = 4'h3 == state ? quene_3 : _GEN_1553; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1704 = 4'h3 == state ? quene_4 : _GEN_1554; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1705 = 4'h3 == state ? quene_5 : _GEN_1555; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1706 = 4'h3 == state ? quene_6 : _GEN_1556; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1707 = 4'h3 == state ? quene_7 : _GEN_1557; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1708 = 4'h3 == state ? quene_8 : _GEN_1558; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1709 = 4'h3 == state ? quene_9 : _GEN_1559; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1710 = 4'h3 == state ? quene_10 : _GEN_1560; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1711 = 4'h3 == state ? quene_11 : _GEN_1561; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1712 = 4'h3 == state ? quene_12 : _GEN_1562; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1713 = 4'h3 == state ? quene_13 : _GEN_1563; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1714 = 4'h3 == state ? quene_14 : _GEN_1564; // @[d_cache.scala 65:18 39:24]
  wire [1:0] _GEN_1715 = 4'h3 == state ? quene_15 : _GEN_1565; // @[d_cache.scala 65:18 39:24]
  wire [127:0] _GEN_1716 = 4'h3 == state ? ram_1_0 : _GEN_1566; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1717 = 4'h3 == state ? ram_1_1 : _GEN_1567; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1718 = 4'h3 == state ? ram_1_2 : _GEN_1568; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1719 = 4'h3 == state ? ram_1_3 : _GEN_1569; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1720 = 4'h3 == state ? ram_1_4 : _GEN_1570; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1721 = 4'h3 == state ? ram_1_5 : _GEN_1571; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1722 = 4'h3 == state ? ram_1_6 : _GEN_1572; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1723 = 4'h3 == state ? ram_1_7 : _GEN_1573; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1724 = 4'h3 == state ? ram_1_8 : _GEN_1574; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1725 = 4'h3 == state ? ram_1_9 : _GEN_1575; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1726 = 4'h3 == state ? ram_1_10 : _GEN_1576; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1727 = 4'h3 == state ? ram_1_11 : _GEN_1577; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1728 = 4'h3 == state ? ram_1_12 : _GEN_1578; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1729 = 4'h3 == state ? ram_1_13 : _GEN_1579; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1730 = 4'h3 == state ? ram_1_14 : _GEN_1580; // @[d_cache.scala 65:18 20:24]
  wire [127:0] _GEN_1731 = 4'h3 == state ? ram_1_15 : _GEN_1581; // @[d_cache.scala 65:18 20:24]
  wire [31:0] _GEN_1732 = 4'h3 == state ? tag_1_0 : _GEN_1582; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1733 = 4'h3 == state ? tag_1_1 : _GEN_1583; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1734 = 4'h3 == state ? tag_1_2 : _GEN_1584; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1735 = 4'h3 == state ? tag_1_3 : _GEN_1585; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1736 = 4'h3 == state ? tag_1_4 : _GEN_1586; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1737 = 4'h3 == state ? tag_1_5 : _GEN_1587; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1738 = 4'h3 == state ? tag_1_6 : _GEN_1588; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1739 = 4'h3 == state ? tag_1_7 : _GEN_1589; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1740 = 4'h3 == state ? tag_1_8 : _GEN_1590; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1741 = 4'h3 == state ? tag_1_9 : _GEN_1591; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1742 = 4'h3 == state ? tag_1_10 : _GEN_1592; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1743 = 4'h3 == state ? tag_1_11 : _GEN_1593; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1744 = 4'h3 == state ? tag_1_12 : _GEN_1594; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1745 = 4'h3 == state ? tag_1_13 : _GEN_1595; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1746 = 4'h3 == state ? tag_1_14 : _GEN_1596; // @[d_cache.scala 65:18 23:24]
  wire [31:0] _GEN_1747 = 4'h3 == state ? tag_1_15 : _GEN_1597; // @[d_cache.scala 65:18 23:24]
  wire  _GEN_1748 = 4'h3 == state ? valid_1_0 : _GEN_1598; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1749 = 4'h3 == state ? valid_1_1 : _GEN_1599; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1750 = 4'h3 == state ? valid_1_2 : _GEN_1600; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1751 = 4'h3 == state ? valid_1_3 : _GEN_1601; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1752 = 4'h3 == state ? valid_1_4 : _GEN_1602; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1753 = 4'h3 == state ? valid_1_5 : _GEN_1603; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1754 = 4'h3 == state ? valid_1_6 : _GEN_1604; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1755 = 4'h3 == state ? valid_1_7 : _GEN_1605; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1756 = 4'h3 == state ? valid_1_8 : _GEN_1606; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1757 = 4'h3 == state ? valid_1_9 : _GEN_1607; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1758 = 4'h3 == state ? valid_1_10 : _GEN_1608; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1759 = 4'h3 == state ? valid_1_11 : _GEN_1609; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1760 = 4'h3 == state ? valid_1_12 : _GEN_1610; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1761 = 4'h3 == state ? valid_1_13 : _GEN_1611; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1762 = 4'h3 == state ? valid_1_14 : _GEN_1612; // @[d_cache.scala 65:18 25:26]
  wire  _GEN_1763 = 4'h3 == state ? valid_1_15 : _GEN_1613; // @[d_cache.scala 65:18 25:26]
  wire [127:0] _GEN_1764 = 4'h3 == state ? write_back_data : _GEN_1614; // @[d_cache.scala 65:18 31:34]
  wire [39:0] _GEN_1765 = 4'h3 == state ? {{8'd0}, write_back_addr} : _GEN_1615; // @[d_cache.scala 65:18 32:34]
  wire  _GEN_1766 = 4'h3 == state ? dirty_0_0 : _GEN_1616; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1767 = 4'h3 == state ? dirty_0_1 : _GEN_1617; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1768 = 4'h3 == state ? dirty_0_2 : _GEN_1618; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1769 = 4'h3 == state ? dirty_0_3 : _GEN_1619; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1770 = 4'h3 == state ? dirty_0_4 : _GEN_1620; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1771 = 4'h3 == state ? dirty_0_5 : _GEN_1621; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1772 = 4'h3 == state ? dirty_0_6 : _GEN_1622; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1773 = 4'h3 == state ? dirty_0_7 : _GEN_1623; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1774 = 4'h3 == state ? dirty_0_8 : _GEN_1624; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1775 = 4'h3 == state ? dirty_0_9 : _GEN_1625; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1776 = 4'h3 == state ? dirty_0_10 : _GEN_1626; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1777 = 4'h3 == state ? dirty_0_11 : _GEN_1627; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1778 = 4'h3 == state ? dirty_0_12 : _GEN_1628; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1779 = 4'h3 == state ? dirty_0_13 : _GEN_1629; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1780 = 4'h3 == state ? dirty_0_14 : _GEN_1630; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1781 = 4'h3 == state ? dirty_0_15 : _GEN_1631; // @[d_cache.scala 65:18 26:26]
  wire  _GEN_1782 = 4'h3 == state ? dirty_1_0 : _GEN_1632; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1783 = 4'h3 == state ? dirty_1_1 : _GEN_1633; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1784 = 4'h3 == state ? dirty_1_2 : _GEN_1634; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1785 = 4'h3 == state ? dirty_1_3 : _GEN_1635; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1786 = 4'h3 == state ? dirty_1_4 : _GEN_1636; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1787 = 4'h3 == state ? dirty_1_5 : _GEN_1637; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1788 = 4'h3 == state ? dirty_1_6 : _GEN_1638; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1789 = 4'h3 == state ? dirty_1_7 : _GEN_1639; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1790 = 4'h3 == state ? dirty_1_8 : _GEN_1640; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1791 = 4'h3 == state ? dirty_1_9 : _GEN_1641; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1792 = 4'h3 == state ? dirty_1_10 : _GEN_1642; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1793 = 4'h3 == state ? dirty_1_11 : _GEN_1643; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1794 = 4'h3 == state ? dirty_1_12 : _GEN_1644; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1795 = 4'h3 == state ? dirty_1_13 : _GEN_1645; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1796 = 4'h3 == state ? dirty_1_14 : _GEN_1646; // @[d_cache.scala 65:18 27:26]
  wire  _GEN_1797 = 4'h3 == state ? dirty_1_15 : _GEN_1647; // @[d_cache.scala 65:18 27:26]
  wire [39:0] _GEN_1947 = 4'h2 == state ? {{8'd0}, write_back_addr} : _GEN_1765; // @[d_cache.scala 65:18 32:34]
  wire [39:0] _GEN_2097 = 4'h1 == state ? {{8'd0}, write_back_addr} : _GEN_1947; // @[d_cache.scala 65:18 32:34]
  wire [39:0] _GEN_2247 = 4'h0 == state ? {{8'd0}, write_back_addr} : _GEN_2097; // @[d_cache.scala 65:18 32:34]
  wire [127:0] _io_to_lsu_rdata_T = _GEN_88 >> shift_bit; // @[d_cache.scala 215:49]
  wire [127:0] _io_to_lsu_rdata_T_1 = _GEN_136 >> shift_bit; // @[d_cache.scala 223:49]
  wire [127:0] _GEN_2248 = way1_hit ? _io_to_lsu_rdata_T_1 : 128'h0; // @[d_cache.scala 222:33 223:33 231:33]
  wire [127:0] _GEN_2251 = way0_hit ? _io_to_lsu_rdata_T : _GEN_2248; // @[d_cache.scala 214:23 215:33]
  wire  _GEN_2253 = way0_hit | way1_hit; // @[d_cache.scala 214:23 217:34]
  wire [63:0] _GEN_2485 = {{32'd0}, io_from_lsu_araddr}; // @[d_cache.scala 290:49]
  wire [63:0] _io_to_axi_araddr_T = _GEN_2485 & 64'hfffffffffffffff0; // @[d_cache.scala 290:49]
  wire  _T_32 = state == 4'h0 & _T_3; // @[d_cache.scala 358:27]
  wire [63:0] _GEN_2255 = state == 4'h0 & _T_3 ? io_from_axi_rdata : 64'h0; // @[d_cache.scala 358:117 359:23 362:29]
  wire  _GEN_2257 = state == 4'h0 & _T_3 & io_from_axi_rvalid; // @[d_cache.scala 358:117 359:23 364:30]
  wire  _GEN_2260 = state == 4'h0 & _T_3 & io_from_axi_bvalid; // @[d_cache.scala 358:117 359:23 367:30]
  wire  _GEN_2265 = state == 4'h0 & _T_3 & io_from_lsu_arvalid; // @[d_cache.scala 358:117 360:23 369:31]
  wire [31:0] _GEN_2267 = state == 4'h0 & _T_3 ? io_from_lsu_awaddr : 32'h0; // @[d_cache.scala 358:117 360:23 375:30]
  wire  _GEN_2271 = state == 4'h0 & _T_3 & io_from_lsu_awvalid; // @[d_cache.scala 358:117 360:23 376:31]
  wire [63:0] _GEN_2272 = state == 4'h0 & _T_3 ? io_from_lsu_wdata : 64'h0; // @[d_cache.scala 358:117 360:23 380:29]
  wire [7:0] _GEN_2273 = state == 4'h0 & _T_3 ? io_from_lsu_wstrb : 8'h0; // @[d_cache.scala 358:117 360:23 381:29]
  wire  _GEN_2275 = state == 4'h0 & _T_3 & io_from_lsu_wvalid; // @[d_cache.scala 358:117 360:23 383:30]
  wire [63:0] _GEN_2278 = state == 4'h7 ? io_from_axi_rdata : _GEN_2255; // @[d_cache.scala 354:30 355:19]
  wire  _GEN_2280 = state == 4'h7 ? io_from_axi_rvalid : _GEN_2257; // @[d_cache.scala 354:30 355:19]
  wire  _GEN_2283 = state == 4'h7 ? io_from_axi_bvalid : _GEN_2260; // @[d_cache.scala 354:30 355:19]
  wire  _GEN_2288 = state == 4'h7 ? io_from_lsu_arvalid : _GEN_2265; // @[d_cache.scala 354:30 356:19]
  wire [31:0] _GEN_2290 = state == 4'h7 ? io_from_lsu_awaddr : _GEN_2267; // @[d_cache.scala 354:30 356:19]
  wire  _GEN_2294 = state == 4'h7 ? io_from_lsu_awvalid : _GEN_2271; // @[d_cache.scala 354:30 356:19]
  wire [63:0] _GEN_2295 = state == 4'h7 ? io_from_lsu_wdata : _GEN_2272; // @[d_cache.scala 354:30 356:19]
  wire [7:0] _GEN_2296 = state == 4'h7 ? io_from_lsu_wstrb : _GEN_2273; // @[d_cache.scala 354:30 356:19]
  wire  _GEN_2298 = state == 4'h7 ? io_from_lsu_wvalid : _GEN_2275; // @[d_cache.scala 354:30 356:19]
  wire  _GEN_2299 = state == 4'h7 | _T_32; // @[d_cache.scala 354:30 356:19]
  wire [63:0] _GEN_2300 = state == 4'h6 ? 64'h0 : _GEN_2278; // @[d_cache.scala 330:35 331:25]
  wire  _GEN_2302 = state == 4'h6 ? 1'h0 : _GEN_2280; // @[d_cache.scala 330:35 333:26]
  wire  _GEN_2305 = state == 4'h6 ? 1'h0 : _GEN_2283; // @[d_cache.scala 330:35 336:26]
  wire  _GEN_2307 = state == 4'h6 ? 1'h0 : _GEN_2288; // @[d_cache.scala 330:35 338:27]
  wire [31:0] _GEN_2308 = state == 4'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 330:35 339:26]
  wire [7:0] _GEN_2309 = state == 4'h6 ? 8'h1 : 8'h0; // @[d_cache.scala 330:35 340:25]
  wire  _GEN_2312 = state == 4'h6 ? 1'h0 : 1'h1; // @[d_cache.scala 330:35 343:26]
  wire [31:0] _GEN_2313 = state == 4'h6 ? write_back_addr : _GEN_2290; // @[d_cache.scala 330:35 344:26]
  wire  _GEN_2314 = state == 4'h6 | _GEN_2294; // @[d_cache.scala 330:35 345:27]
  wire [63:0] _GEN_2318 = state == 4'h6 ? write_back_data[63:0] : _GEN_2295; // @[d_cache.scala 330:35 349:25]
  wire [7:0] _GEN_2319 = state == 4'h6 ? 8'hff : _GEN_2296; // @[d_cache.scala 330:35 350:25]
  wire  _GEN_2321 = state == 4'h6 | _GEN_2298; // @[d_cache.scala 330:35 352:26]
  wire  _GEN_2322 = state == 4'h6 | _GEN_2299; // @[d_cache.scala 330:35 353:26]
  wire [63:0] _GEN_2323 = state == 4'h4 | state == 4'h8 ? 64'h0 : _GEN_2300; // @[d_cache.scala 305:50 306:25]
  wire  _GEN_2325 = state == 4'h4 | state == 4'h8 ? 1'h0 : _GEN_2302; // @[d_cache.scala 305:50 308:26]
  wire  _GEN_2328 = state == 4'h4 | state == 4'h8 ? io_from_axi_bvalid : _GEN_2305; // @[d_cache.scala 305:50 311:26]
  wire  _GEN_2330 = state == 4'h4 | state == 4'h8 ? 1'h0 : _GEN_2307; // @[d_cache.scala 305:50 313:27]
  wire [31:0] _GEN_2331 = state == 4'h4 | state == 4'h8 ? 32'h0 : _GEN_2308; // @[d_cache.scala 305:50 314:26]
  wire [7:0] _GEN_2332 = state == 4'h4 | state == 4'h8 ? 8'h0 : _GEN_2309; // @[d_cache.scala 305:50 315:25]
  wire  _GEN_2335 = state == 4'h4 | state == 4'h8 | _GEN_2312; // @[d_cache.scala 305:50 318:26]
  wire [31:0] _GEN_2336 = state == 4'h4 | state == 4'h8 ? io_from_lsu_awaddr : _GEN_2313; // @[d_cache.scala 305:50 319:26]
  wire  _GEN_2337 = state == 4'h4 | state == 4'h8 ? io_from_lsu_awvalid : _GEN_2314; // @[d_cache.scala 305:50 320:27]
  wire [63:0] _GEN_2341 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wdata : _GEN_2318; // @[d_cache.scala 305:50 324:25]
  wire [7:0] _GEN_2342 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wstrb : _GEN_2319; // @[d_cache.scala 305:50 325:25]
  wire  _GEN_2344 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wvalid : _GEN_2321; // @[d_cache.scala 305:50 327:26]
  wire  _GEN_2345 = state == 4'h4 | state == 4'h8 | _GEN_2322; // @[d_cache.scala 305:50 328:26]
  wire [63:0] _GEN_2346 = state == 4'h3 ? 64'h0 : _GEN_2323; // @[d_cache.scala 281:31 282:25]
  wire  _GEN_2348 = state == 4'h3 ? 1'h0 : _GEN_2325; // @[d_cache.scala 281:31 284:26]
  wire  _GEN_2351 = state == 4'h3 ? 1'h0 : _GEN_2328; // @[d_cache.scala 281:31 287:26]
  wire  _GEN_2353 = state == 4'h3 | _GEN_2330; // @[d_cache.scala 281:31 289:27]
  wire [63:0] _GEN_2354 = state == 4'h3 ? _io_to_axi_araddr_T : {{32'd0}, _GEN_2331}; // @[d_cache.scala 281:31 290:26]
  wire [7:0] _GEN_2355 = state == 4'h3 ? 8'h1 : _GEN_2332; // @[d_cache.scala 281:31 291:25]
  wire  _GEN_2358 = state == 4'h3 | _GEN_2335; // @[d_cache.scala 281:31 294:26]
  wire [31:0] _GEN_2359 = state == 4'h3 ? 32'h0 : _GEN_2336; // @[d_cache.scala 281:31 295:26]
  wire  _GEN_2360 = state == 4'h3 ? 1'h0 : _GEN_2337; // @[d_cache.scala 281:31 296:27]
  wire [7:0] _GEN_2361 = state == 4'h3 ? 8'h0 : _GEN_2332; // @[d_cache.scala 281:31 297:25]
  wire [63:0] _GEN_2364 = state == 4'h3 ? 64'h0 : _GEN_2341; // @[d_cache.scala 281:31 300:25]
  wire [7:0] _GEN_2365 = state == 4'h3 ? 8'h0 : _GEN_2342; // @[d_cache.scala 281:31 301:25]
  wire  _GEN_2367 = state == 4'h3 ? 1'h0 : _GEN_2344; // @[d_cache.scala 281:31 303:26]
  wire  _GEN_2368 = state == 4'h3 ? 1'h0 : _GEN_2345; // @[d_cache.scala 281:31 304:26]
  wire  _GEN_2369 = state == 4'h2 ? 1'h0 : _GEN_2353; // @[d_cache.scala 239:33 240:27]
  wire [63:0] _GEN_2370 = state == 4'h2 ? {{32'd0}, io_from_lsu_araddr} : _GEN_2354; // @[d_cache.scala 239:33 241:26]
  wire [7:0] _GEN_2371 = state == 4'h2 ? 8'h0 : _GEN_2355; // @[d_cache.scala 239:33 242:25]
  wire  _GEN_2374 = state == 4'h2 ? 1'h0 : _GEN_2358; // @[d_cache.scala 239:33 245:26]
  wire [31:0] _GEN_2375 = state == 4'h2 ? 32'h0 : _GEN_2359; // @[d_cache.scala 239:33 246:26]
  wire  _GEN_2376 = state == 4'h2 ? 1'h0 : _GEN_2360; // @[d_cache.scala 239:33 247:27]
  wire [7:0] _GEN_2377 = state == 4'h2 ? 8'h0 : _GEN_2361; // @[d_cache.scala 239:33 248:25]
  wire [63:0] _GEN_2380 = state == 4'h2 ? 64'h0 : _GEN_2364; // @[d_cache.scala 239:33 251:25]
  wire [7:0] _GEN_2381 = state == 4'h2 ? 8'h0 : _GEN_2365; // @[d_cache.scala 239:33 252:25]
  wire  _GEN_2383 = state == 4'h2 ? 1'h0 : _GEN_2367; // @[d_cache.scala 239:33 254:26]
  wire  _GEN_2384 = state == 4'h2 ? 1'h0 : _GEN_2368; // @[d_cache.scala 239:33 255:26]
  wire [63:0] _GEN_2385 = state == 4'h2 ? 64'h0 : _GEN_2346; // @[d_cache.scala 239:33]
  wire  _GEN_2387 = state == 4'h2 ? 1'h0 : _GEN_2348; // @[d_cache.scala 239:33]
  wire  _GEN_2391 = state == 4'h2 ? _GEN_2253 : _GEN_2351; // @[d_cache.scala 239:33]
  wire [63:0] _GEN_2393 = state == 4'h1 ? {{32'd0}, io_from_lsu_araddr} : _GEN_2370; // @[d_cache.scala 197:27 199:26]
  wire [127:0] _GEN_2408 = state == 4'h1 ? _GEN_2251 : {{64'd0}, _GEN_2385}; // @[d_cache.scala 197:27]
  wire [39:0] _GEN_2486 = reset ? 40'h0 : _GEN_2247; // @[d_cache.scala 32:{34,34}]
  assign io_to_lsu_rdata = _GEN_2408[63:0];
  assign io_to_lsu_rvalid = state == 4'h1 ? _GEN_2253 : _GEN_2387; // @[d_cache.scala 197:27]
  assign io_to_lsu_bvalid = state == 4'h1 ? 1'h0 : _GEN_2391; // @[d_cache.scala 197:27]
  assign io_to_axi_araddr = _GEN_2393[31:0];
  assign io_to_axi_arlen = state == 4'h1 ? 8'h0 : _GEN_2371; // @[d_cache.scala 197:27 200:25]
  assign io_to_axi_arvalid = state == 4'h1 ? 1'h0 : _GEN_2369; // @[d_cache.scala 197:27 198:27]
  assign io_to_axi_rready = state == 4'h1 ? 1'h0 : _GEN_2374; // @[d_cache.scala 197:27 203:26]
  assign io_to_axi_awaddr = state == 4'h1 ? 32'h0 : _GEN_2375; // @[d_cache.scala 197:27 204:26]
  assign io_to_axi_awlen = state == 4'h1 ? 8'h0 : _GEN_2377; // @[d_cache.scala 197:27 206:25]
  assign io_to_axi_awvalid = state == 4'h1 ? 1'h0 : _GEN_2376; // @[d_cache.scala 197:27 205:27]
  assign io_to_axi_wdata = state == 4'h1 ? 64'h0 : _GEN_2380; // @[d_cache.scala 197:27 209:25]
  assign io_to_axi_wstrb = state == 4'h1 ? 8'h0 : _GEN_2381; // @[d_cache.scala 197:27 210:25]
  assign io_to_axi_wvalid = state == 4'h1 ? 1'h0 : _GEN_2383; // @[d_cache.scala 197:27 212:26]
  assign io_to_axi_bready = state == 4'h1 ? 1'h0 : _GEN_2384; // @[d_cache.scala 197:27 213:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_0 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_0 <= _GEN_203;
        end else begin
          ram_0_0 <= _GEN_1652;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_1 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_1 <= _GEN_204;
        end else begin
          ram_0_1 <= _GEN_1653;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_2 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_2 <= _GEN_205;
        end else begin
          ram_0_2 <= _GEN_1654;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_3 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_3 <= _GEN_206;
        end else begin
          ram_0_3 <= _GEN_1655;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_4 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_4 <= _GEN_207;
        end else begin
          ram_0_4 <= _GEN_1656;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_5 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_5 <= _GEN_208;
        end else begin
          ram_0_5 <= _GEN_1657;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_6 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_6 <= _GEN_209;
        end else begin
          ram_0_6 <= _GEN_1658;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_7 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_7 <= _GEN_210;
        end else begin
          ram_0_7 <= _GEN_1659;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_8 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_8 <= _GEN_211;
        end else begin
          ram_0_8 <= _GEN_1660;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_9 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_9 <= _GEN_212;
        end else begin
          ram_0_9 <= _GEN_1661;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_10 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_10 <= _GEN_213;
        end else begin
          ram_0_10 <= _GEN_1662;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_11 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_11 <= _GEN_214;
        end else begin
          ram_0_11 <= _GEN_1663;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_12 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_12 <= _GEN_215;
        end else begin
          ram_0_12 <= _GEN_1664;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_13 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_13 <= _GEN_216;
        end else begin
          ram_0_13 <= _GEN_1665;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_14 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_14 <= _GEN_217;
        end else begin
          ram_0_14 <= _GEN_1666;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_15 <= 128'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_0_15 <= _GEN_218;
        end else begin
          ram_0_15 <= _GEN_1667;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_0 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_0 <= _GEN_235;
        end else begin
          ram_1_0 <= _GEN_1716;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_1 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_1 <= _GEN_236;
        end else begin
          ram_1_1 <= _GEN_1717;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_2 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_2 <= _GEN_237;
        end else begin
          ram_1_2 <= _GEN_1718;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_3 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_3 <= _GEN_238;
        end else begin
          ram_1_3 <= _GEN_1719;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_4 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_4 <= _GEN_239;
        end else begin
          ram_1_4 <= _GEN_1720;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_5 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_5 <= _GEN_240;
        end else begin
          ram_1_5 <= _GEN_1721;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_6 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_6 <= _GEN_241;
        end else begin
          ram_1_6 <= _GEN_1722;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_7 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_7 <= _GEN_242;
        end else begin
          ram_1_7 <= _GEN_1723;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_8 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_8 <= _GEN_243;
        end else begin
          ram_1_8 <= _GEN_1724;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_9 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_9 <= _GEN_244;
        end else begin
          ram_1_9 <= _GEN_1725;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_10 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_10 <= _GEN_245;
        end else begin
          ram_1_10 <= _GEN_1726;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_11 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_11 <= _GEN_246;
        end else begin
          ram_1_11 <= _GEN_1727;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_12 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_12 <= _GEN_247;
        end else begin
          ram_1_12 <= _GEN_1728;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_13 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_13 <= _GEN_248;
        end else begin
          ram_1_13 <= _GEN_1729;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_14 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_14 <= _GEN_249;
        end else begin
          ram_1_14 <= _GEN_1730;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_15 <= 128'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          ram_1_15 <= _GEN_250;
        end else begin
          ram_1_15 <= _GEN_1731;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_0 <= _GEN_1668;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_1 <= _GEN_1669;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_2 <= _GEN_1670;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_3 <= _GEN_1671;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_4 <= _GEN_1672;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_5 <= _GEN_1673;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_6 <= _GEN_1674;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_7 <= _GEN_1675;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_8 <= _GEN_1676;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_9 <= _GEN_1677;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_10 <= _GEN_1678;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_11 <= _GEN_1679;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_12 <= _GEN_1680;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_13 <= _GEN_1681;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_14 <= _GEN_1682;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_0_15 <= _GEN_1683;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_0 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_0 <= _GEN_1732;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_1 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_1 <= _GEN_1733;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_2 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_2 <= _GEN_1734;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_3 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_3 <= _GEN_1735;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_4 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_4 <= _GEN_1736;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_5 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_5 <= _GEN_1737;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_6 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_6 <= _GEN_1738;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_7 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_7 <= _GEN_1739;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_8 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_8 <= _GEN_1740;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_9 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_9 <= _GEN_1741;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_10 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_10 <= _GEN_1742;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_11 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_11 <= _GEN_1743;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_12 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_12 <= _GEN_1744;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_13 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_13 <= _GEN_1745;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_14 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_14 <= _GEN_1746;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 23:24]
      tag_1_15 <= 32'h0; // @[d_cache.scala 23:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          tag_1_15 <= _GEN_1747;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_0 <= _GEN_1684;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_1 <= _GEN_1685;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_2 <= _GEN_1686;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_3 <= _GEN_1687;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_4 <= _GEN_1688;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_5 <= _GEN_1689;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_6 <= _GEN_1690;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_7 <= _GEN_1691;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_8 <= _GEN_1692;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_9 <= _GEN_1693;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_10 <= _GEN_1694;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_11 <= _GEN_1695;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_12 <= _GEN_1696;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_13 <= _GEN_1697;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_14 <= _GEN_1698;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 24:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_0_15 <= _GEN_1699;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_0 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_0 <= _GEN_1748;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_1 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_1 <= _GEN_1749;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_2 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_2 <= _GEN_1750;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_3 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_3 <= _GEN_1751;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_4 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_4 <= _GEN_1752;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_5 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_5 <= _GEN_1753;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_6 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_6 <= _GEN_1754;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_7 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_7 <= _GEN_1755;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_8 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_8 <= _GEN_1756;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_9 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_9 <= _GEN_1757;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_10 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_10 <= _GEN_1758;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_11 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_11 <= _GEN_1759;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_12 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_12 <= _GEN_1760;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_13 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_13 <= _GEN_1761;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_14 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_14 <= _GEN_1762;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:26]
      valid_1_15 <= 1'h0; // @[d_cache.scala 25:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          valid_1_15 <= _GEN_1763;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_0 <= _GEN_219;
        end else begin
          dirty_0_0 <= _GEN_1766;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_1 <= _GEN_220;
        end else begin
          dirty_0_1 <= _GEN_1767;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_2 <= _GEN_221;
        end else begin
          dirty_0_2 <= _GEN_1768;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_3 <= _GEN_222;
        end else begin
          dirty_0_3 <= _GEN_1769;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_4 <= _GEN_223;
        end else begin
          dirty_0_4 <= _GEN_1770;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_5 <= _GEN_224;
        end else begin
          dirty_0_5 <= _GEN_1771;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_6 <= _GEN_225;
        end else begin
          dirty_0_6 <= _GEN_1772;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_7 <= _GEN_226;
        end else begin
          dirty_0_7 <= _GEN_1773;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_8 <= _GEN_227;
        end else begin
          dirty_0_8 <= _GEN_1774;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_9 <= _GEN_228;
        end else begin
          dirty_0_9 <= _GEN_1775;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_10 <= _GEN_229;
        end else begin
          dirty_0_10 <= _GEN_1776;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_11 <= _GEN_230;
        end else begin
          dirty_0_11 <= _GEN_1777;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_12 <= _GEN_231;
        end else begin
          dirty_0_12 <= _GEN_1778;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_13 <= _GEN_232;
        end else begin
          dirty_0_13 <= _GEN_1779;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_14 <= _GEN_233;
        end else begin
          dirty_0_14 <= _GEN_1780;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 26:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_0_15 <= _GEN_234;
        end else begin
          dirty_0_15 <= _GEN_1781;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_0 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_0 <= _GEN_251;
        end else begin
          dirty_1_0 <= _GEN_1782;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_1 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_1 <= _GEN_252;
        end else begin
          dirty_1_1 <= _GEN_1783;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_2 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_2 <= _GEN_253;
        end else begin
          dirty_1_2 <= _GEN_1784;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_3 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_3 <= _GEN_254;
        end else begin
          dirty_1_3 <= _GEN_1785;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_4 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_4 <= _GEN_255;
        end else begin
          dirty_1_4 <= _GEN_1786;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_5 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_5 <= _GEN_256;
        end else begin
          dirty_1_5 <= _GEN_1787;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_6 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_6 <= _GEN_257;
        end else begin
          dirty_1_6 <= _GEN_1788;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_7 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_7 <= _GEN_258;
        end else begin
          dirty_1_7 <= _GEN_1789;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_8 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_8 <= _GEN_259;
        end else begin
          dirty_1_8 <= _GEN_1790;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_9 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_9 <= _GEN_260;
        end else begin
          dirty_1_9 <= _GEN_1791;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_10 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_10 <= _GEN_261;
        end else begin
          dirty_1_10 <= _GEN_1792;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_11 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_11 <= _GEN_262;
        end else begin
          dirty_1_11 <= _GEN_1793;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_12 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_12 <= _GEN_263;
        end else begin
          dirty_1_12 <= _GEN_1794;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_13 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_13 <= _GEN_264;
        end else begin
          dirty_1_13 <= _GEN_1795;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_14 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_14 <= _GEN_265;
        end else begin
          dirty_1_14 <= _GEN_1796;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:26]
      dirty_1_15 <= 1'h0; // @[d_cache.scala 27:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (4'h2 == state) begin // @[d_cache.scala 65:18]
          dirty_1_15 <= _GEN_266;
        end else begin
          dirty_1_15 <= _GEN_1797;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:34]
      write_back_data <= 128'h0; // @[d_cache.scala 31:34]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          write_back_data <= _GEN_1764;
        end
      end
    end
    write_back_addr <= _GEN_2486[31:0]; // @[d_cache.scala 32:{34,34}]
    if (reset) begin // @[d_cache.scala 37:31]
      receive_data_0 <= 64'h0; // @[d_cache.scala 37:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          receive_data_0 <= _GEN_1648;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:31]
      receive_data_1 <= 64'h0; // @[d_cache.scala 37:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          receive_data_1 <= _GEN_1649;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 38:30]
      receive_num <= 3'h0; // @[d_cache.scala 38:30]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (4'h1 == state) begin // @[d_cache.scala 65:18]
        if (!(way0_hit)) begin // @[d_cache.scala 76:27]
          receive_num <= _GEN_69;
        end
      end else if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
        receive_num <= _GEN_1650;
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_0 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_0 <= _GEN_1700;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_1 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_1 <= _GEN_1701;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_2 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_2 <= _GEN_1702;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_3 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_3 <= _GEN_1703;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_4 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_4 <= _GEN_1704;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_5 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_5 <= _GEN_1705;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_6 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_6 <= _GEN_1706;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_7 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_7 <= _GEN_1707;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_8 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_8 <= _GEN_1708;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_9 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_9 <= _GEN_1709;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_10 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_10 <= _GEN_1710;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_11 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_11 <= _GEN_1711;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_12 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_12 <= _GEN_1712;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_13 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_13 <= _GEN_1713;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_14 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_14 <= _GEN_1714;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 39:24]
      quene_15 <= 2'h0; // @[d_cache.scala 39:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 65:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 65:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 65:18]
          quene_15 <= _GEN_1715;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 60:24]
      state <= 4'h0; // @[d_cache.scala 60:24]
    end else if (4'h0 == state) begin // @[d_cache.scala 65:18]
      if ((io_from_lsu_arvalid | io_from_lsu_awvalid) & io_from_lsu_araddr >= 32'ha0000000) begin // @[d_cache.scala 67:99]
        state <= 4'h0; // @[d_cache.scala 68:23]
      end else if (io_from_lsu_arvalid) begin // @[d_cache.scala 69:44]
        state <= 4'h1; // @[d_cache.scala 70:23]
      end else begin
        state <= _GEN_64;
      end
    end else if (4'h1 == state) begin // @[d_cache.scala 65:18]
      if (way0_hit) begin // @[d_cache.scala 76:27]
        state <= 4'h0;
      end else begin
        state <= _GEN_68;
      end
    end else if (4'h2 == state) begin // @[d_cache.scala 65:18]
      state <= _GEN_202;
    end else begin
      state <= _GEN_1651;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  ram_0_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  ram_0_1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  ram_0_2 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  ram_0_3 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  ram_0_4 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  ram_0_5 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  ram_0_6 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  ram_0_7 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  ram_0_8 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  ram_0_9 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  ram_0_10 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  ram_0_11 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  ram_0_12 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  ram_0_13 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  ram_0_14 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  ram_0_15 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  ram_1_0 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  ram_1_1 = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  ram_1_2 = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  ram_1_3 = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  ram_1_4 = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  ram_1_5 = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  ram_1_6 = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  ram_1_7 = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  ram_1_8 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  ram_1_9 = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  ram_1_10 = _RAND_26[127:0];
  _RAND_27 = {4{`RANDOM}};
  ram_1_11 = _RAND_27[127:0];
  _RAND_28 = {4{`RANDOM}};
  ram_1_12 = _RAND_28[127:0];
  _RAND_29 = {4{`RANDOM}};
  ram_1_13 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  ram_1_14 = _RAND_30[127:0];
  _RAND_31 = {4{`RANDOM}};
  ram_1_15 = _RAND_31[127:0];
  _RAND_32 = {1{`RANDOM}};
  tag_0_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  tag_0_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  tag_0_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  tag_0_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  tag_0_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  tag_0_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  tag_0_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  tag_0_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  tag_0_8 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  tag_0_9 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  tag_0_10 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  tag_0_11 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  tag_0_12 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  tag_0_13 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  tag_0_14 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  tag_0_15 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  tag_1_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  tag_1_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  tag_1_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  tag_1_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  tag_1_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  tag_1_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  tag_1_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  tag_1_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  tag_1_8 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  tag_1_9 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  tag_1_10 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  tag_1_11 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  tag_1_12 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  tag_1_13 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  tag_1_14 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  tag_1_15 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  valid_0_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_0_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_0_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_0_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_0_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_0_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_0_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_0_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_0_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_0_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_0_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_0_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_0_12 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_0_13 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_0_14 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_0_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_1_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_1_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_1_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_1_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_1_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_1_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_1_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_1_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_1_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_1_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_1_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_1_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_1_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_1_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_1_15 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  dirty_0_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  dirty_0_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dirty_0_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  dirty_0_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  dirty_0_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dirty_0_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  dirty_0_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  dirty_0_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dirty_0_8 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  dirty_0_9 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  dirty_0_10 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  dirty_0_11 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  dirty_0_12 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  dirty_0_13 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dirty_0_14 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  dirty_0_15 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  dirty_1_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  dirty_1_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  dirty_1_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  dirty_1_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dirty_1_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  dirty_1_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  dirty_1_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  dirty_1_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  dirty_1_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  dirty_1_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  dirty_1_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  dirty_1_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  dirty_1_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  dirty_1_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  dirty_1_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  dirty_1_15 = _RAND_127[0:0];
  _RAND_128 = {4{`RANDOM}};
  write_back_data = _RAND_128[127:0];
  _RAND_129 = {1{`RANDOM}};
  write_back_addr = _RAND_129[31:0];
  _RAND_130 = {2{`RANDOM}};
  receive_data_0 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  receive_data_1 = _RAND_131[63:0];
  _RAND_132 = {1{`RANDOM}};
  receive_num = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  quene_0 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  quene_1 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  quene_2 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  quene_3 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  quene_4 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  quene_5 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  quene_6 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  quene_7 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  quene_8 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  quene_9 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  quene_10 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  quene_11 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  quene_12 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  quene_13 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  quene_14 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  quene_15 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  state = _RAND_149[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI(
  input         clock,
  input         reset,
  input  [31:0] io_axi_in_araddr,
  input  [7:0]  io_axi_in_arlen,
  input         io_axi_in_arvalid,
  input         io_axi_in_rready,
  input  [31:0] io_axi_in_awaddr,
  input  [7:0]  io_axi_in_awlen,
  input         io_axi_in_awvalid,
  input  [63:0] io_axi_in_wdata,
  input  [7:0]  io_axi_in_wstrb,
  input         io_axi_in_wvalid,
  input         io_axi_in_bready,
  output [63:0] io_axi_out_rdata,
  output        io_axi_out_rlast,
  output        io_axi_out_rvalid,
  output        io_axi_out_wready,
  output        io_axi_out_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] Mem_modle_Raddr; // @[AXI.scala 30:27]
  wire [63:0] Mem_modle_Rdata; // @[AXI.scala 30:27]
  wire [63:0] Mem_modle_Waddr; // @[AXI.scala 30:27]
  wire [63:0] Mem_modle_Wdata; // @[AXI.scala 30:27]
  wire [7:0] Mem_modle_Wmask; // @[AXI.scala 30:27]
  wire  Mem_modle_Write_en; // @[AXI.scala 30:27]
  wire  Mem_modle_Read_en; // @[AXI.scala 30:27]
  reg  axi_wready; // @[AXI.scala 14:29]
  reg  axi_bvalid; // @[AXI.scala 17:29]
  reg  axi_rvalid; // @[AXI.scala 21:29]
  reg [7:0] arlen; // @[AXI.scala 22:24]
  reg [7:0] awlen; // @[AXI.scala 23:24]
  reg [63:0] araddr; // @[AXI.scala 24:25]
  reg [63:0] awaddr; // @[AXI.scala 25:25]
  reg [2:0] state; // @[AXI.scala 28:24]
  wire  _GEN_4 = io_axi_in_arvalid | axi_rvalid; // @[AXI.scala 55:42 60:28 21:29]
  wire  _GEN_7 = io_axi_in_awvalid & io_axi_in_wvalid | axi_wready; // @[AXI.scala 43:56 46:28 14:29]
  wire [63:0] _awaddr_T_1 = awaddr + 64'h8; // @[AXI.scala 72:38]
  wire [7:0] _awlen_T_1 = awlen - 8'h1; // @[AXI.scala 73:36]
  wire [63:0] _GEN_14 = io_axi_in_wvalid & axi_wready ? _awaddr_T_1 : awaddr; // @[AXI.scala 25:25 71:60 72:28]
  wire [7:0] _GEN_15 = io_axi_in_wvalid & axi_wready ? _awlen_T_1 : awlen; // @[AXI.scala 23:24 71:60 73:27]
  wire  _GEN_18 = awlen == 8'h0 | axi_bvalid; // @[AXI.scala 64:30 68:28 17:29]
  wire  _T_7 = arlen == 8'h0; // @[AXI.scala 78:23]
  wire [2:0] _GEN_22 = io_axi_in_rready ? 3'h0 : state; // @[AXI.scala 28:24 79:39 80:27]
  wire  _GEN_24 = io_axi_in_rready ? 1'h0 : axi_rvalid; // @[AXI.scala 21:29 79:39 82:32]
  wire [63:0] _araddr_T_1 = araddr + 64'h8; // @[AXI.scala 86:38]
  wire [7:0] _arlen_T_1 = arlen - 8'h1; // @[AXI.scala 87:36]
  wire [63:0] _GEN_25 = io_axi_in_rready ? _araddr_T_1 : araddr; // @[AXI.scala 24:25 85:39 86:28]
  wire [7:0] _GEN_26 = io_axi_in_rready ? _arlen_T_1 : arlen; // @[AXI.scala 22:24 85:39 87:27]
  wire [2:0] _GEN_27 = arlen == 8'h0 ? _GEN_22 : state; // @[AXI.scala 28:24 78:30]
  wire  _GEN_29 = arlen == 8'h0 ? _GEN_24 : axi_rvalid; // @[AXI.scala 21:29 78:30]
  wire [63:0] _GEN_30 = arlen == 8'h0 ? araddr : _GEN_25; // @[AXI.scala 24:25 78:30]
  wire [7:0] _GEN_31 = arlen == 8'h0 ? arlen : _GEN_26; // @[AXI.scala 22:24 78:30]
  wire [2:0] _GEN_32 = io_axi_in_bready ? 3'h0 : state; // @[AXI.scala 92:35 93:23 28:24]
  wire  _GEN_33 = io_axi_in_bready ? 1'h0 : axi_bvalid; // @[AXI.scala 92:35 94:28 17:29]
  wire [2:0] _GEN_35 = 3'h3 == state ? _GEN_32 : state; // @[AXI.scala 41:18 28:24]
  wire  _GEN_36 = 3'h3 == state ? _GEN_33 : axi_bvalid; // @[AXI.scala 41:18 17:29]
  MEM Mem_modle ( // @[AXI.scala 30:27]
    .Raddr(Mem_modle_Raddr),
    .Rdata(Mem_modle_Rdata),
    .Waddr(Mem_modle_Waddr),
    .Wdata(Mem_modle_Wdata),
    .Wmask(Mem_modle_Wmask),
    .Write_en(Mem_modle_Write_en),
    .Read_en(Mem_modle_Read_en)
  );
  assign io_axi_out_rdata = Mem_modle_Rdata; // @[AXI.scala 108:22]
  assign io_axi_out_rlast = state == 3'h1 & _T_7; // @[AXI.scala 110:41]
  assign io_axi_out_rvalid = axi_rvalid; // @[AXI.scala 109:23]
  assign io_axi_out_wready = axi_wready; // @[AXI.scala 112:23]
  assign io_axi_out_bvalid = axi_bvalid; // @[AXI.scala 113:23]
  assign Mem_modle_Raddr = araddr; // @[AXI.scala 31:24]
  assign Mem_modle_Waddr = awaddr; // @[AXI.scala 32:24]
  assign Mem_modle_Wdata = io_axi_in_wdata; // @[AXI.scala 33:24]
  assign Mem_modle_Wmask = io_axi_in_wstrb; // @[AXI.scala 34:24]
  assign Mem_modle_Write_en = axi_wready; // @[AXI.scala 35:27]
  assign Mem_modle_Read_en = axi_rvalid; // @[AXI.scala 36:26]
  always @(posedge clock) begin
    if (reset) begin // @[AXI.scala 14:29]
      axi_wready <= 1'h0; // @[AXI.scala 14:29]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      axi_wready <= _GEN_7;
    end else if (3'h2 == state) begin // @[AXI.scala 41:18]
      if (awlen == 8'h0) begin // @[AXI.scala 64:30]
        axi_wready <= 1'h0; // @[AXI.scala 65:28]
      end
    end
    if (reset) begin // @[AXI.scala 17:29]
      axi_bvalid <= 1'h0; // @[AXI.scala 17:29]
    end else if (!(3'h0 == state)) begin // @[AXI.scala 41:18]
      if (3'h2 == state) begin // @[AXI.scala 41:18]
        axi_bvalid <= _GEN_18;
      end else if (!(3'h1 == state)) begin // @[AXI.scala 41:18]
        axi_bvalid <= _GEN_36;
      end
    end
    if (reset) begin // @[AXI.scala 21:29]
      axi_rvalid <= 1'h0; // @[AXI.scala 21:29]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 43:56]
        axi_rvalid <= _GEN_4;
      end
    end else if (!(3'h2 == state)) begin // @[AXI.scala 41:18]
      if (3'h1 == state) begin // @[AXI.scala 41:18]
        axi_rvalid <= _GEN_29;
      end
    end
    if (reset) begin // @[AXI.scala 22:24]
      arlen <= 8'h0; // @[AXI.scala 22:24]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 43:56]
        if (io_axi_in_arvalid) begin // @[AXI.scala 55:42]
          arlen <= io_axi_in_arlen; // @[AXI.scala 57:23]
        end
      end
    end else if (!(3'h2 == state)) begin // @[AXI.scala 41:18]
      if (3'h1 == state) begin // @[AXI.scala 41:18]
        arlen <= _GEN_31;
      end
    end
    if (reset) begin // @[AXI.scala 23:24]
      awlen <= 8'h0; // @[AXI.scala 23:24]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 43:56]
        awlen <= io_axi_in_awlen; // @[AXI.scala 48:23]
      end
    end else if (3'h2 == state) begin // @[AXI.scala 41:18]
      if (!(awlen == 8'h0)) begin // @[AXI.scala 64:30]
        awlen <= _GEN_15;
      end
    end
    if (reset) begin // @[AXI.scala 24:25]
      araddr <= 64'h0; // @[AXI.scala 24:25]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 43:56]
        if (io_axi_in_arvalid) begin // @[AXI.scala 55:42]
          araddr <= {{32'd0}, io_axi_in_araddr}; // @[AXI.scala 58:24]
        end
      end
    end else if (!(3'h2 == state)) begin // @[AXI.scala 41:18]
      if (3'h1 == state) begin // @[AXI.scala 41:18]
        araddr <= _GEN_30;
      end
    end
    if (reset) begin // @[AXI.scala 25:25]
      awaddr <= 64'h0; // @[AXI.scala 25:25]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 43:56]
        awaddr <= {{32'd0}, io_axi_in_awaddr}; // @[AXI.scala 49:24]
      end
    end else if (3'h2 == state) begin // @[AXI.scala 41:18]
      if (!(awlen == 8'h0)) begin // @[AXI.scala 64:30]
        awaddr <= _GEN_14;
      end
    end
    if (reset) begin // @[AXI.scala 28:24]
      state <= 3'h0; // @[AXI.scala 28:24]
    end else if (3'h0 == state) begin // @[AXI.scala 41:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 43:56]
        state <= 3'h2; // @[AXI.scala 44:23]
      end else if (io_axi_in_arvalid) begin // @[AXI.scala 55:42]
        state <= 3'h1; // @[AXI.scala 56:23]
      end
    end else if (3'h2 == state) begin // @[AXI.scala 41:18]
      if (awlen == 8'h0) begin // @[AXI.scala 64:30]
        state <= 3'h3; // @[AXI.scala 69:23]
      end
    end else if (3'h1 == state) begin // @[AXI.scala 41:18]
      state <= _GEN_27;
    end else begin
      state <= _GEN_35;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_wready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_bvalid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_rvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  arlen = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  awlen = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  araddr = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  awaddr = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input         clock,
  input         reset,
  output [31:0] io_inst,
  output [63:0] io_pc,
  output        io_step
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  Register_clock; // @[top.scala 15:25]
  wire [4:0] Register_io_raddr1; // @[top.scala 15:25]
  wire [4:0] Register_io_raddr2; // @[top.scala 15:25]
  wire [63:0] Register_io_rdata1; // @[top.scala 15:25]
  wire [63:0] Register_io_rdata2; // @[top.scala 15:25]
  wire  Register_io_we; // @[top.scala 15:25]
  wire [4:0] Register_io_waddr; // @[top.scala 15:25]
  wire [63:0] Register_io_wdata; // @[top.scala 15:25]
  wire  IFU_clock; // @[top.scala 16:21]
  wire  IFU_reset; // @[top.scala 16:21]
  wire  IFU_io_ds_allowin; // @[top.scala 16:21]
  wire  IFU_io_ds_ready_go; // @[top.scala 16:21]
  wire  IFU_io_ds_valid; // @[top.scala 16:21]
  wire  IFU_io_br_taken; // @[top.scala 16:21]
  wire [63:0] IFU_io_br_target; // @[top.scala 16:21]
  wire [63:0] IFU_io_to_ds_pc; // @[top.scala 16:21]
  wire  IFU_io_fs_to_ds_valid; // @[top.scala 16:21]
  wire [31:0] IFU_io_inst; // @[top.scala 16:21]
  wire  IFU_io_axi_in_arready; // @[top.scala 16:21]
  wire [63:0] IFU_io_axi_in_rdata; // @[top.scala 16:21]
  wire  IFU_io_axi_in_rvalid; // @[top.scala 16:21]
  wire [31:0] IFU_io_axi_out_araddr; // @[top.scala 16:21]
  wire  IFU_io_axi_out_arvalid; // @[top.scala 16:21]
  wire  IFU_io_axi_out_rready; // @[top.scala 16:21]
  wire  IFU_io_fence; // @[top.scala 16:21]
  wire  IFU_io_clear_cache; // @[top.scala 16:21]
  wire  IFU_io_cache_init; // @[top.scala 16:21]
  wire  IDU_clock; // @[top.scala 17:21]
  wire  IDU_reset; // @[top.scala 17:21]
  wire [63:0] IDU_io_pc; // @[top.scala 17:21]
  wire  IDU_io_fs_to_ds_valid; // @[top.scala 17:21]
  wire  IDU_io_ds_to_es_valid; // @[top.scala 17:21]
  wire  IDU_io_es_allowin; // @[top.scala 17:21]
  wire [31:0] IDU_io_from_fs_inst; // @[top.scala 17:21]
  wire  IDU_io_br_taken; // @[top.scala 17:21]
  wire [63:0] IDU_io_br_target; // @[top.scala 17:21]
  wire  IDU_io_ds_allowin; // @[top.scala 17:21]
  wire  IDU_io_ds_ready_go; // @[top.scala 17:21]
  wire  IDU_io_fence; // @[top.scala 17:21]
  wire [4:0] IDU_io_raddr1; // @[top.scala 17:21]
  wire [4:0] IDU_io_raddr2; // @[top.scala 17:21]
  wire [63:0] IDU_io_rdata1; // @[top.scala 17:21]
  wire [63:0] IDU_io_rdata2; // @[top.scala 17:21]
  wire [63:0] IDU_io_to_es_pc; // @[top.scala 17:21]
  wire [31:0] IDU_io_ALUop; // @[top.scala 17:21]
  wire [63:0] IDU_io_src1; // @[top.scala 17:21]
  wire [63:0] IDU_io_src2; // @[top.scala 17:21]
  wire [4:0] IDU_io_rf_dst; // @[top.scala 17:21]
  wire [63:0] IDU_io_store_data; // @[top.scala 17:21]
  wire  IDU_io_ctrl_sign_reg_write; // @[top.scala 17:21]
  wire  IDU_io_ctrl_sign_Writemem_en; // @[top.scala 17:21]
  wire  IDU_io_ctrl_sign_Readmem_en; // @[top.scala 17:21]
  wire [7:0] IDU_io_ctrl_sign_Wmask; // @[top.scala 17:21]
  wire [2:0] IDU_io_load_type; // @[top.scala 17:21]
  wire  IDU_io_es_ld; // @[top.scala 17:21]
  wire [63:0] IDU_io_es_fwd_res; // @[top.scala 17:21]
  wire [63:0] IDU_io_ms_fwd_res; // @[top.scala 17:21]
  wire [63:0] IDU_io_ws_fwd_res; // @[top.scala 17:21]
  wire  IDU_io_es_fwd_ready; // @[top.scala 17:21]
  wire  IDU_io_ms_fwd_ready; // @[top.scala 17:21]
  wire  IDU_io_es_rf_we; // @[top.scala 17:21]
  wire  IDU_io_ms_rf_we; // @[top.scala 17:21]
  wire  IDU_io_ws_rf_we; // @[top.scala 17:21]
  wire  IDU_io_es_valid; // @[top.scala 17:21]
  wire  IDU_io_ms_valid; // @[top.scala 17:21]
  wire  IDU_io_ws_valid; // @[top.scala 17:21]
  wire [4:0] IDU_io_es_rf_dst; // @[top.scala 17:21]
  wire [4:0] IDU_io_ms_rf_dst; // @[top.scala 17:21]
  wire [4:0] IDU_io_ws_rf_dst; // @[top.scala 17:21]
  wire  IDU_io_ds_valid; // @[top.scala 17:21]
  wire  EXU_clock; // @[top.scala 18:21]
  wire  EXU_reset; // @[top.scala 18:21]
  wire [63:0] EXU_io_pc; // @[top.scala 18:21]
  wire  EXU_io_ds_to_es_valid; // @[top.scala 18:21]
  wire  EXU_io_ms_allowin; // @[top.scala 18:21]
  wire  EXU_io_es_allowin; // @[top.scala 18:21]
  wire [31:0] EXU_io_ALUop; // @[top.scala 18:21]
  wire [63:0] EXU_io_src1_value; // @[top.scala 18:21]
  wire [63:0] EXU_io_src2_value; // @[top.scala 18:21]
  wire [4:0] EXU_io_rf_dst; // @[top.scala 18:21]
  wire [63:0] EXU_io_store_data; // @[top.scala 18:21]
  wire  EXU_io_es_to_ms_valid; // @[top.scala 18:21]
  wire [2:0] EXU_io_load_type; // @[top.scala 18:21]
  wire [63:0] EXU_io_to_ms_pc; // @[top.scala 18:21]
  wire [63:0] EXU_io_to_ms_alures; // @[top.scala 18:21]
  wire [63:0] EXU_io_to_ms_store_data; // @[top.scala 18:21]
  wire  EXU_io_to_ms_wen; // @[top.scala 18:21]
  wire [7:0] EXU_io_to_ms_wstrb; // @[top.scala 18:21]
  wire  EXU_io_to_ms_ren; // @[top.scala 18:21]
  wire [63:0] EXU_io_to_ms_maddr; // @[top.scala 18:21]
  wire [4:0] EXU_io_to_ms_rf_dst; // @[top.scala 18:21]
  wire  EXU_io_to_ms_rf_we; // @[top.scala 18:21]
  wire [2:0] EXU_io_to_ms_load_type; // @[top.scala 18:21]
  wire  EXU_io_ctrl_sign_reg_write; // @[top.scala 18:21]
  wire  EXU_io_ctrl_sign_Writemem_en; // @[top.scala 18:21]
  wire  EXU_io_ctrl_sign_Readmem_en; // @[top.scala 18:21]
  wire [7:0] EXU_io_ctrl_sign_Wmask; // @[top.scala 18:21]
  wire  EXU_io_es_valid; // @[top.scala 18:21]
  wire  EXU_io_es_rf_we; // @[top.scala 18:21]
  wire [4:0] EXU_io_es_rf_dst; // @[top.scala 18:21]
  wire  EXU_io_es_fwd_ready; // @[top.scala 18:21]
  wire [63:0] EXU_io_es_fwd_res; // @[top.scala 18:21]
  wire  EXU_io_es_ld; // @[top.scala 18:21]
  wire  LSU_clock; // @[top.scala 19:21]
  wire  LSU_reset; // @[top.scala 19:21]
  wire [63:0] LSU_io_pc; // @[top.scala 19:21]
  wire  LSU_io_es_to_ms_valid; // @[top.scala 19:21]
  wire  LSU_io_ms_allowin; // @[top.scala 19:21]
  wire  LSU_io_rf_we; // @[top.scala 19:21]
  wire [4:0] LSU_io_rf_dst; // @[top.scala 19:21]
  wire [63:0] LSU_io_alu_res; // @[top.scala 19:21]
  wire [63:0] LSU_io_store_data; // @[top.scala 19:21]
  wire [2:0] LSU_io_load_type; // @[top.scala 19:21]
  wire  LSU_io_wen; // @[top.scala 19:21]
  wire [7:0] LSU_io_wstrb; // @[top.scala 19:21]
  wire  LSU_io_ren; // @[top.scala 19:21]
  wire [63:0] LSU_io_maddr; // @[top.scala 19:21]
  wire [63:0] LSU_io_to_ws_pc; // @[top.scala 19:21]
  wire [63:0] LSU_io_ms_final_res; // @[top.scala 19:21]
  wire  LSU_io_ms_to_ws_valid; // @[top.scala 19:21]
  wire  LSU_io_to_ws_rf_we; // @[top.scala 19:21]
  wire [4:0] LSU_io_to_ws_rf_dst; // @[top.scala 19:21]
  wire  LSU_io_ms_valid; // @[top.scala 19:21]
  wire  LSU_io_ms_rf_we; // @[top.scala 19:21]
  wire [4:0] LSU_io_ms_rf_dst; // @[top.scala 19:21]
  wire  LSU_io_ms_fwd_ready; // @[top.scala 19:21]
  wire [63:0] LSU_io_ms_fwd_res; // @[top.scala 19:21]
  wire [63:0] LSU_io_axi_in_rdata; // @[top.scala 19:21]
  wire  LSU_io_axi_in_rvalid; // @[top.scala 19:21]
  wire  LSU_io_axi_in_bvalid; // @[top.scala 19:21]
  wire [31:0] LSU_io_axi_out_araddr; // @[top.scala 19:21]
  wire  LSU_io_axi_out_arvalid; // @[top.scala 19:21]
  wire [31:0] LSU_io_axi_out_awaddr; // @[top.scala 19:21]
  wire  LSU_io_axi_out_awvalid; // @[top.scala 19:21]
  wire [63:0] LSU_io_axi_out_wdata; // @[top.scala 19:21]
  wire [7:0] LSU_io_axi_out_wstrb; // @[top.scala 19:21]
  wire  LSU_io_axi_out_wvalid; // @[top.scala 19:21]
  wire  WBU_clock; // @[top.scala 20:21]
  wire  WBU_reset; // @[top.scala 20:21]
  wire [63:0] WBU_io_pc; // @[top.scala 20:21]
  wire  WBU_io_ms_to_ws_valid; // @[top.scala 20:21]
  wire [63:0] WBU_io_ms_final_res; // @[top.scala 20:21]
  wire  WBU_io_rf_we; // @[top.scala 20:21]
  wire [4:0] WBU_io_rf_dst; // @[top.scala 20:21]
  wire  WBU_io_we; // @[top.scala 20:21]
  wire [4:0] WBU_io_waddr; // @[top.scala 20:21]
  wire [63:0] WBU_io_wdata; // @[top.scala 20:21]
  wire  WBU_io_ws_valid; // @[top.scala 20:21]
  wire  WBU_io_ws_rf_we; // @[top.scala 20:21]
  wire [4:0] WBU_io_ws_rf_dst; // @[top.scala 20:21]
  wire [63:0] WBU_io_ws_fwd_res; // @[top.scala 20:21]
  wire [63:0] WBU_io_ws_pc; // @[top.scala 20:21]
  wire  arbiter_clock; // @[top.scala 21:25]
  wire  arbiter_reset; // @[top.scala 21:25]
  wire [31:0] arbiter_io_ifu_axi_in_araddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_ifu_axi_in_arlen; // @[top.scala 21:25]
  wire  arbiter_io_ifu_axi_in_arvalid; // @[top.scala 21:25]
  wire  arbiter_io_ifu_axi_in_rready; // @[top.scala 21:25]
  wire [63:0] arbiter_io_ifu_axi_out_rdata; // @[top.scala 21:25]
  wire  arbiter_io_ifu_axi_out_rlast; // @[top.scala 21:25]
  wire  arbiter_io_ifu_axi_out_rvalid; // @[top.scala 21:25]
  wire [31:0] arbiter_io_lsu_axi_in_araddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_lsu_axi_in_arlen; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_arvalid; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_rready; // @[top.scala 21:25]
  wire [31:0] arbiter_io_lsu_axi_in_awaddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_lsu_axi_in_awlen; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_awvalid; // @[top.scala 21:25]
  wire [63:0] arbiter_io_lsu_axi_in_wdata; // @[top.scala 21:25]
  wire [7:0] arbiter_io_lsu_axi_in_wstrb; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_wvalid; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_in_bready; // @[top.scala 21:25]
  wire [63:0] arbiter_io_lsu_axi_out_rdata; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_out_rlast; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_out_rvalid; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_out_wready; // @[top.scala 21:25]
  wire  arbiter_io_lsu_axi_out_bvalid; // @[top.scala 21:25]
  wire [63:0] arbiter_io_axi_in_rdata; // @[top.scala 21:25]
  wire  arbiter_io_axi_in_rlast; // @[top.scala 21:25]
  wire  arbiter_io_axi_in_rvalid; // @[top.scala 21:25]
  wire  arbiter_io_axi_in_wready; // @[top.scala 21:25]
  wire  arbiter_io_axi_in_bvalid; // @[top.scala 21:25]
  wire [31:0] arbiter_io_axi_out_araddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_axi_out_arlen; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_arvalid; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_rready; // @[top.scala 21:25]
  wire [31:0] arbiter_io_axi_out_awaddr; // @[top.scala 21:25]
  wire [7:0] arbiter_io_axi_out_awlen; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_awvalid; // @[top.scala 21:25]
  wire [63:0] arbiter_io_axi_out_wdata; // @[top.scala 21:25]
  wire [7:0] arbiter_io_axi_out_wstrb; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_wvalid; // @[top.scala 21:25]
  wire  arbiter_io_axi_out_bready; // @[top.scala 21:25]
  wire  i_cache_clock; // @[top.scala 22:25]
  wire  i_cache_reset; // @[top.scala 22:25]
  wire [31:0] i_cache_io_from_ifu_araddr; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_from_ifu_rready; // @[top.scala 22:25]
  wire  i_cache_io_to_ifu_arready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_to_ifu_rdata; // @[top.scala 22:25]
  wire  i_cache_io_to_ifu_rvalid; // @[top.scala 22:25]
  wire [31:0] i_cache_io_to_axi_araddr; // @[top.scala 22:25]
  wire [7:0] i_cache_io_to_axi_arlen; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_arvalid; // @[top.scala 22:25]
  wire  i_cache_io_to_axi_rready; // @[top.scala 22:25]
  wire [63:0] i_cache_io_from_axi_rdata; // @[top.scala 22:25]
  wire  i_cache_io_from_axi_rlast; // @[top.scala 22:25]
  wire  i_cache_io_from_axi_rvalid; // @[top.scala 22:25]
  wire  i_cache_io_cache_init; // @[top.scala 22:25]
  wire  i_cache_io_clear_cache; // @[top.scala 22:25]
  wire  d_cache_clock; // @[top.scala 23:25]
  wire  d_cache_reset; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_araddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_arvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_from_lsu_awaddr; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_awvalid; // @[top.scala 23:25]
  wire [63:0] d_cache_io_from_lsu_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_from_lsu_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_from_lsu_wvalid; // @[top.scala 23:25]
  wire [63:0] d_cache_io_to_lsu_rdata; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_lsu_bvalid; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_araddr; // @[top.scala 23:25]
  wire [7:0] d_cache_io_to_axi_arlen; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_arvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_rready; // @[top.scala 23:25]
  wire [31:0] d_cache_io_to_axi_awaddr; // @[top.scala 23:25]
  wire [7:0] d_cache_io_to_axi_awlen; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_awvalid; // @[top.scala 23:25]
  wire [63:0] d_cache_io_to_axi_wdata; // @[top.scala 23:25]
  wire [7:0] d_cache_io_to_axi_wstrb; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_wvalid; // @[top.scala 23:25]
  wire  d_cache_io_to_axi_bready; // @[top.scala 23:25]
  wire [63:0] d_cache_io_from_axi_rdata; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_rlast; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_rvalid; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_wready; // @[top.scala 23:25]
  wire  d_cache_io_from_axi_bvalid; // @[top.scala 23:25]
  wire  axi_clock; // @[top.scala 24:21]
  wire  axi_reset; // @[top.scala 24:21]
  wire [31:0] axi_io_axi_in_araddr; // @[top.scala 24:21]
  wire [7:0] axi_io_axi_in_arlen; // @[top.scala 24:21]
  wire  axi_io_axi_in_arvalid; // @[top.scala 24:21]
  wire  axi_io_axi_in_rready; // @[top.scala 24:21]
  wire [31:0] axi_io_axi_in_awaddr; // @[top.scala 24:21]
  wire [7:0] axi_io_axi_in_awlen; // @[top.scala 24:21]
  wire  axi_io_axi_in_awvalid; // @[top.scala 24:21]
  wire [63:0] axi_io_axi_in_wdata; // @[top.scala 24:21]
  wire [7:0] axi_io_axi_in_wstrb; // @[top.scala 24:21]
  wire  axi_io_axi_in_wvalid; // @[top.scala 24:21]
  wire  axi_io_axi_in_bready; // @[top.scala 24:21]
  wire [63:0] axi_io_axi_out_rdata; // @[top.scala 24:21]
  wire  axi_io_axi_out_rlast; // @[top.scala 24:21]
  wire  axi_io_axi_out_rvalid; // @[top.scala 24:21]
  wire  axi_io_axi_out_wready; // @[top.scala 24:21]
  wire  axi_io_axi_out_bvalid; // @[top.scala 24:21]
  wire [31:0] dpi_flag; // @[top.scala 116:21]
  wire [31:0] dpi_ecall_flag; // @[top.scala 116:21]
  wire [63:0] dpi_pc; // @[top.scala 116:21]
  reg  diff_step; // @[top.scala 113:28]
  wire [63:0] _dpi_io_pc_T = IDU_io_ds_valid ? EXU_io_pc : IDU_io_pc; // @[top.scala 119:96]
  wire [63:0] _dpi_io_pc_T_1 = EXU_io_es_valid ? LSU_io_pc : _dpi_io_pc_T; // @[top.scala 119:72]
  wire [63:0] _dpi_io_pc_T_2 = LSU_io_ms_valid ? WBU_io_pc : _dpi_io_pc_T_1; // @[top.scala 119:48]
  Register Register ( // @[top.scala 15:25]
    .clock(Register_clock),
    .io_raddr1(Register_io_raddr1),
    .io_raddr2(Register_io_raddr2),
    .io_rdata1(Register_io_rdata1),
    .io_rdata2(Register_io_rdata2),
    .io_we(Register_io_we),
    .io_waddr(Register_io_waddr),
    .io_wdata(Register_io_wdata)
  );
  IFU IFU ( // @[top.scala 16:21]
    .clock(IFU_clock),
    .reset(IFU_reset),
    .io_ds_allowin(IFU_io_ds_allowin),
    .io_ds_ready_go(IFU_io_ds_ready_go),
    .io_ds_valid(IFU_io_ds_valid),
    .io_br_taken(IFU_io_br_taken),
    .io_br_target(IFU_io_br_target),
    .io_to_ds_pc(IFU_io_to_ds_pc),
    .io_fs_to_ds_valid(IFU_io_fs_to_ds_valid),
    .io_inst(IFU_io_inst),
    .io_axi_in_arready(IFU_io_axi_in_arready),
    .io_axi_in_rdata(IFU_io_axi_in_rdata),
    .io_axi_in_rvalid(IFU_io_axi_in_rvalid),
    .io_axi_out_araddr(IFU_io_axi_out_araddr),
    .io_axi_out_arvalid(IFU_io_axi_out_arvalid),
    .io_axi_out_rready(IFU_io_axi_out_rready),
    .io_fence(IFU_io_fence),
    .io_clear_cache(IFU_io_clear_cache),
    .io_cache_init(IFU_io_cache_init)
  );
  IDU IDU ( // @[top.scala 17:21]
    .clock(IDU_clock),
    .reset(IDU_reset),
    .io_pc(IDU_io_pc),
    .io_fs_to_ds_valid(IDU_io_fs_to_ds_valid),
    .io_ds_to_es_valid(IDU_io_ds_to_es_valid),
    .io_es_allowin(IDU_io_es_allowin),
    .io_from_fs_inst(IDU_io_from_fs_inst),
    .io_br_taken(IDU_io_br_taken),
    .io_br_target(IDU_io_br_target),
    .io_ds_allowin(IDU_io_ds_allowin),
    .io_ds_ready_go(IDU_io_ds_ready_go),
    .io_fence(IDU_io_fence),
    .io_raddr1(IDU_io_raddr1),
    .io_raddr2(IDU_io_raddr2),
    .io_rdata1(IDU_io_rdata1),
    .io_rdata2(IDU_io_rdata2),
    .io_to_es_pc(IDU_io_to_es_pc),
    .io_ALUop(IDU_io_ALUop),
    .io_src1(IDU_io_src1),
    .io_src2(IDU_io_src2),
    .io_rf_dst(IDU_io_rf_dst),
    .io_store_data(IDU_io_store_data),
    .io_ctrl_sign_reg_write(IDU_io_ctrl_sign_reg_write),
    .io_ctrl_sign_Writemem_en(IDU_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(IDU_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(IDU_io_ctrl_sign_Wmask),
    .io_load_type(IDU_io_load_type),
    .io_es_ld(IDU_io_es_ld),
    .io_es_fwd_res(IDU_io_es_fwd_res),
    .io_ms_fwd_res(IDU_io_ms_fwd_res),
    .io_ws_fwd_res(IDU_io_ws_fwd_res),
    .io_es_fwd_ready(IDU_io_es_fwd_ready),
    .io_ms_fwd_ready(IDU_io_ms_fwd_ready),
    .io_es_rf_we(IDU_io_es_rf_we),
    .io_ms_rf_we(IDU_io_ms_rf_we),
    .io_ws_rf_we(IDU_io_ws_rf_we),
    .io_es_valid(IDU_io_es_valid),
    .io_ms_valid(IDU_io_ms_valid),
    .io_ws_valid(IDU_io_ws_valid),
    .io_es_rf_dst(IDU_io_es_rf_dst),
    .io_ms_rf_dst(IDU_io_ms_rf_dst),
    .io_ws_rf_dst(IDU_io_ws_rf_dst),
    .io_ds_valid(IDU_io_ds_valid)
  );
  EXU EXU ( // @[top.scala 18:21]
    .clock(EXU_clock),
    .reset(EXU_reset),
    .io_pc(EXU_io_pc),
    .io_ds_to_es_valid(EXU_io_ds_to_es_valid),
    .io_ms_allowin(EXU_io_ms_allowin),
    .io_es_allowin(EXU_io_es_allowin),
    .io_ALUop(EXU_io_ALUop),
    .io_src1_value(EXU_io_src1_value),
    .io_src2_value(EXU_io_src2_value),
    .io_rf_dst(EXU_io_rf_dst),
    .io_store_data(EXU_io_store_data),
    .io_es_to_ms_valid(EXU_io_es_to_ms_valid),
    .io_load_type(EXU_io_load_type),
    .io_to_ms_pc(EXU_io_to_ms_pc),
    .io_to_ms_alures(EXU_io_to_ms_alures),
    .io_to_ms_store_data(EXU_io_to_ms_store_data),
    .io_to_ms_wen(EXU_io_to_ms_wen),
    .io_to_ms_wstrb(EXU_io_to_ms_wstrb),
    .io_to_ms_ren(EXU_io_to_ms_ren),
    .io_to_ms_maddr(EXU_io_to_ms_maddr),
    .io_to_ms_rf_dst(EXU_io_to_ms_rf_dst),
    .io_to_ms_rf_we(EXU_io_to_ms_rf_we),
    .io_to_ms_load_type(EXU_io_to_ms_load_type),
    .io_ctrl_sign_reg_write(EXU_io_ctrl_sign_reg_write),
    .io_ctrl_sign_Writemem_en(EXU_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(EXU_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(EXU_io_ctrl_sign_Wmask),
    .io_es_valid(EXU_io_es_valid),
    .io_es_rf_we(EXU_io_es_rf_we),
    .io_es_rf_dst(EXU_io_es_rf_dst),
    .io_es_fwd_ready(EXU_io_es_fwd_ready),
    .io_es_fwd_res(EXU_io_es_fwd_res),
    .io_es_ld(EXU_io_es_ld)
  );
  LSU LSU ( // @[top.scala 19:21]
    .clock(LSU_clock),
    .reset(LSU_reset),
    .io_pc(LSU_io_pc),
    .io_es_to_ms_valid(LSU_io_es_to_ms_valid),
    .io_ms_allowin(LSU_io_ms_allowin),
    .io_rf_we(LSU_io_rf_we),
    .io_rf_dst(LSU_io_rf_dst),
    .io_alu_res(LSU_io_alu_res),
    .io_store_data(LSU_io_store_data),
    .io_load_type(LSU_io_load_type),
    .io_wen(LSU_io_wen),
    .io_wstrb(LSU_io_wstrb),
    .io_ren(LSU_io_ren),
    .io_maddr(LSU_io_maddr),
    .io_to_ws_pc(LSU_io_to_ws_pc),
    .io_ms_final_res(LSU_io_ms_final_res),
    .io_ms_to_ws_valid(LSU_io_ms_to_ws_valid),
    .io_to_ws_rf_we(LSU_io_to_ws_rf_we),
    .io_to_ws_rf_dst(LSU_io_to_ws_rf_dst),
    .io_ms_valid(LSU_io_ms_valid),
    .io_ms_rf_we(LSU_io_ms_rf_we),
    .io_ms_rf_dst(LSU_io_ms_rf_dst),
    .io_ms_fwd_ready(LSU_io_ms_fwd_ready),
    .io_ms_fwd_res(LSU_io_ms_fwd_res),
    .io_axi_in_rdata(LSU_io_axi_in_rdata),
    .io_axi_in_rvalid(LSU_io_axi_in_rvalid),
    .io_axi_in_bvalid(LSU_io_axi_in_bvalid),
    .io_axi_out_araddr(LSU_io_axi_out_araddr),
    .io_axi_out_arvalid(LSU_io_axi_out_arvalid),
    .io_axi_out_awaddr(LSU_io_axi_out_awaddr),
    .io_axi_out_awvalid(LSU_io_axi_out_awvalid),
    .io_axi_out_wdata(LSU_io_axi_out_wdata),
    .io_axi_out_wstrb(LSU_io_axi_out_wstrb),
    .io_axi_out_wvalid(LSU_io_axi_out_wvalid)
  );
  WBU WBU ( // @[top.scala 20:21]
    .clock(WBU_clock),
    .reset(WBU_reset),
    .io_pc(WBU_io_pc),
    .io_ms_to_ws_valid(WBU_io_ms_to_ws_valid),
    .io_ms_final_res(WBU_io_ms_final_res),
    .io_rf_we(WBU_io_rf_we),
    .io_rf_dst(WBU_io_rf_dst),
    .io_we(WBU_io_we),
    .io_waddr(WBU_io_waddr),
    .io_wdata(WBU_io_wdata),
    .io_ws_valid(WBU_io_ws_valid),
    .io_ws_rf_we(WBU_io_ws_rf_we),
    .io_ws_rf_dst(WBU_io_ws_rf_dst),
    .io_ws_fwd_res(WBU_io_ws_fwd_res),
    .io_ws_pc(WBU_io_ws_pc)
  );
  AXI_ARBITER arbiter ( // @[top.scala 21:25]
    .clock(arbiter_clock),
    .reset(arbiter_reset),
    .io_ifu_axi_in_araddr(arbiter_io_ifu_axi_in_araddr),
    .io_ifu_axi_in_arlen(arbiter_io_ifu_axi_in_arlen),
    .io_ifu_axi_in_arvalid(arbiter_io_ifu_axi_in_arvalid),
    .io_ifu_axi_in_rready(arbiter_io_ifu_axi_in_rready),
    .io_ifu_axi_out_rdata(arbiter_io_ifu_axi_out_rdata),
    .io_ifu_axi_out_rlast(arbiter_io_ifu_axi_out_rlast),
    .io_ifu_axi_out_rvalid(arbiter_io_ifu_axi_out_rvalid),
    .io_lsu_axi_in_araddr(arbiter_io_lsu_axi_in_araddr),
    .io_lsu_axi_in_arlen(arbiter_io_lsu_axi_in_arlen),
    .io_lsu_axi_in_arvalid(arbiter_io_lsu_axi_in_arvalid),
    .io_lsu_axi_in_rready(arbiter_io_lsu_axi_in_rready),
    .io_lsu_axi_in_awaddr(arbiter_io_lsu_axi_in_awaddr),
    .io_lsu_axi_in_awlen(arbiter_io_lsu_axi_in_awlen),
    .io_lsu_axi_in_awvalid(arbiter_io_lsu_axi_in_awvalid),
    .io_lsu_axi_in_wdata(arbiter_io_lsu_axi_in_wdata),
    .io_lsu_axi_in_wstrb(arbiter_io_lsu_axi_in_wstrb),
    .io_lsu_axi_in_wvalid(arbiter_io_lsu_axi_in_wvalid),
    .io_lsu_axi_in_bready(arbiter_io_lsu_axi_in_bready),
    .io_lsu_axi_out_rdata(arbiter_io_lsu_axi_out_rdata),
    .io_lsu_axi_out_rlast(arbiter_io_lsu_axi_out_rlast),
    .io_lsu_axi_out_rvalid(arbiter_io_lsu_axi_out_rvalid),
    .io_lsu_axi_out_wready(arbiter_io_lsu_axi_out_wready),
    .io_lsu_axi_out_bvalid(arbiter_io_lsu_axi_out_bvalid),
    .io_axi_in_rdata(arbiter_io_axi_in_rdata),
    .io_axi_in_rlast(arbiter_io_axi_in_rlast),
    .io_axi_in_rvalid(arbiter_io_axi_in_rvalid),
    .io_axi_in_wready(arbiter_io_axi_in_wready),
    .io_axi_in_bvalid(arbiter_io_axi_in_bvalid),
    .io_axi_out_araddr(arbiter_io_axi_out_araddr),
    .io_axi_out_arlen(arbiter_io_axi_out_arlen),
    .io_axi_out_arvalid(arbiter_io_axi_out_arvalid),
    .io_axi_out_rready(arbiter_io_axi_out_rready),
    .io_axi_out_awaddr(arbiter_io_axi_out_awaddr),
    .io_axi_out_awlen(arbiter_io_axi_out_awlen),
    .io_axi_out_awvalid(arbiter_io_axi_out_awvalid),
    .io_axi_out_wdata(arbiter_io_axi_out_wdata),
    .io_axi_out_wstrb(arbiter_io_axi_out_wstrb),
    .io_axi_out_wvalid(arbiter_io_axi_out_wvalid),
    .io_axi_out_bready(arbiter_io_axi_out_bready)
  );
  I_CACHE i_cache ( // @[top.scala 22:25]
    .clock(i_cache_clock),
    .reset(i_cache_reset),
    .io_from_ifu_araddr(i_cache_io_from_ifu_araddr),
    .io_from_ifu_arvalid(i_cache_io_from_ifu_arvalid),
    .io_from_ifu_rready(i_cache_io_from_ifu_rready),
    .io_to_ifu_arready(i_cache_io_to_ifu_arready),
    .io_to_ifu_rdata(i_cache_io_to_ifu_rdata),
    .io_to_ifu_rvalid(i_cache_io_to_ifu_rvalid),
    .io_to_axi_araddr(i_cache_io_to_axi_araddr),
    .io_to_axi_arlen(i_cache_io_to_axi_arlen),
    .io_to_axi_arvalid(i_cache_io_to_axi_arvalid),
    .io_to_axi_rready(i_cache_io_to_axi_rready),
    .io_from_axi_rdata(i_cache_io_from_axi_rdata),
    .io_from_axi_rlast(i_cache_io_from_axi_rlast),
    .io_from_axi_rvalid(i_cache_io_from_axi_rvalid),
    .io_cache_init(i_cache_io_cache_init),
    .io_clear_cache(i_cache_io_clear_cache)
  );
  D_CACHE d_cache ( // @[top.scala 23:25]
    .clock(d_cache_clock),
    .reset(d_cache_reset),
    .io_from_lsu_araddr(d_cache_io_from_lsu_araddr),
    .io_from_lsu_arvalid(d_cache_io_from_lsu_arvalid),
    .io_from_lsu_awaddr(d_cache_io_from_lsu_awaddr),
    .io_from_lsu_awvalid(d_cache_io_from_lsu_awvalid),
    .io_from_lsu_wdata(d_cache_io_from_lsu_wdata),
    .io_from_lsu_wstrb(d_cache_io_from_lsu_wstrb),
    .io_from_lsu_wvalid(d_cache_io_from_lsu_wvalid),
    .io_to_lsu_rdata(d_cache_io_to_lsu_rdata),
    .io_to_lsu_rvalid(d_cache_io_to_lsu_rvalid),
    .io_to_lsu_bvalid(d_cache_io_to_lsu_bvalid),
    .io_to_axi_araddr(d_cache_io_to_axi_araddr),
    .io_to_axi_arlen(d_cache_io_to_axi_arlen),
    .io_to_axi_arvalid(d_cache_io_to_axi_arvalid),
    .io_to_axi_rready(d_cache_io_to_axi_rready),
    .io_to_axi_awaddr(d_cache_io_to_axi_awaddr),
    .io_to_axi_awlen(d_cache_io_to_axi_awlen),
    .io_to_axi_awvalid(d_cache_io_to_axi_awvalid),
    .io_to_axi_wdata(d_cache_io_to_axi_wdata),
    .io_to_axi_wstrb(d_cache_io_to_axi_wstrb),
    .io_to_axi_wvalid(d_cache_io_to_axi_wvalid),
    .io_to_axi_bready(d_cache_io_to_axi_bready),
    .io_from_axi_rdata(d_cache_io_from_axi_rdata),
    .io_from_axi_rlast(d_cache_io_from_axi_rlast),
    .io_from_axi_rvalid(d_cache_io_from_axi_rvalid),
    .io_from_axi_wready(d_cache_io_from_axi_wready),
    .io_from_axi_bvalid(d_cache_io_from_axi_bvalid)
  );
  AXI axi ( // @[top.scala 24:21]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_axi_in_araddr(axi_io_axi_in_araddr),
    .io_axi_in_arlen(axi_io_axi_in_arlen),
    .io_axi_in_arvalid(axi_io_axi_in_arvalid),
    .io_axi_in_rready(axi_io_axi_in_rready),
    .io_axi_in_awaddr(axi_io_axi_in_awaddr),
    .io_axi_in_awlen(axi_io_axi_in_awlen),
    .io_axi_in_awvalid(axi_io_axi_in_awvalid),
    .io_axi_in_wdata(axi_io_axi_in_wdata),
    .io_axi_in_wstrb(axi_io_axi_in_wstrb),
    .io_axi_in_wvalid(axi_io_axi_in_wvalid),
    .io_axi_in_bready(axi_io_axi_in_bready),
    .io_axi_out_rdata(axi_io_axi_out_rdata),
    .io_axi_out_rlast(axi_io_axi_out_rlast),
    .io_axi_out_rvalid(axi_io_axi_out_rvalid),
    .io_axi_out_wready(axi_io_axi_out_wready),
    .io_axi_out_bvalid(axi_io_axi_out_bvalid)
  );
  DPI dpi ( // @[top.scala 116:21]
    .flag(dpi_flag),
    .ecall_flag(dpi_ecall_flag),
    .pc(dpi_pc)
  );
  assign io_inst = IFU_io_inst; // @[top.scala 112:13]
  assign io_pc = IFU_io_to_ds_pc; // @[top.scala 110:11]
  assign io_step = diff_step; // @[top.scala 115:13]
  assign Register_clock = clock;
  assign Register_io_raddr1 = IDU_io_raddr1; // @[top.scala 56:20]
  assign Register_io_raddr2 = IDU_io_raddr2; // @[top.scala 57:20]
  assign Register_io_we = WBU_io_we; // @[top.scala 106:16]
  assign Register_io_waddr = WBU_io_waddr; // @[top.scala 107:19]
  assign Register_io_wdata = WBU_io_wdata; // @[top.scala 108:19]
  assign IFU_clock = clock;
  assign IFU_reset = reset;
  assign IFU_io_ds_allowin = IDU_io_ds_allowin; // @[top.scala 44:20]
  assign IFU_io_ds_ready_go = IDU_io_ds_ready_go; // @[top.scala 43:21]
  assign IFU_io_ds_valid = IDU_io_ds_valid; // @[top.scala 42:18]
  assign IFU_io_br_taken = IDU_io_br_taken; // @[top.scala 45:18]
  assign IFU_io_br_target = IDU_io_br_target; // @[top.scala 46:19]
  assign IFU_io_axi_in_arready = i_cache_io_to_ifu_arready; // @[top.scala 29:16]
  assign IFU_io_axi_in_rdata = i_cache_io_to_ifu_rdata; // @[top.scala 29:16]
  assign IFU_io_axi_in_rvalid = i_cache_io_to_ifu_rvalid; // @[top.scala 29:16]
  assign IFU_io_fence = IDU_io_fence; // @[top.scala 48:15]
  assign IFU_io_cache_init = i_cache_io_cache_init; // @[top.scala 49:20]
  assign IDU_clock = clock;
  assign IDU_reset = reset;
  assign IDU_io_pc = IFU_io_to_ds_pc; // @[top.scala 52:12]
  assign IDU_io_fs_to_ds_valid = IFU_io_fs_to_ds_valid; // @[top.scala 53:24]
  assign IDU_io_es_allowin = EXU_io_es_allowin; // @[top.scala 54:20]
  assign IDU_io_from_fs_inst = IFU_io_inst; // @[top.scala 55:22]
  assign IDU_io_rdata1 = Register_io_rdata1; // @[top.scala 58:16]
  assign IDU_io_rdata2 = Register_io_rdata2; // @[top.scala 59:16]
  assign IDU_io_es_ld = EXU_io_es_ld; // @[top.scala 75:15]
  assign IDU_io_es_fwd_res = EXU_io_es_fwd_res; // @[top.scala 70:20]
  assign IDU_io_ms_fwd_res = LSU_io_ms_fwd_res; // @[top.scala 72:20]
  assign IDU_io_ws_fwd_res = WBU_io_ws_fwd_res; // @[top.scala 74:20]
  assign IDU_io_es_fwd_ready = EXU_io_es_fwd_ready; // @[top.scala 69:22]
  assign IDU_io_ms_fwd_ready = LSU_io_ms_fwd_ready; // @[top.scala 71:22]
  assign IDU_io_es_rf_we = EXU_io_es_rf_we; // @[top.scala 62:18]
  assign IDU_io_ms_rf_we = LSU_io_ms_rf_we; // @[top.scala 65:18]
  assign IDU_io_ws_rf_we = WBU_io_ws_rf_we; // @[top.scala 68:18]
  assign IDU_io_es_valid = EXU_io_es_valid; // @[top.scala 60:18]
  assign IDU_io_ms_valid = LSU_io_ms_valid; // @[top.scala 63:18]
  assign IDU_io_ws_valid = WBU_io_ws_valid; // @[top.scala 66:18]
  assign IDU_io_es_rf_dst = EXU_io_es_rf_dst; // @[top.scala 61:19]
  assign IDU_io_ms_rf_dst = LSU_io_ms_rf_dst; // @[top.scala 64:19]
  assign IDU_io_ws_rf_dst = WBU_io_ws_rf_dst; // @[top.scala 67:19]
  assign EXU_clock = clock;
  assign EXU_reset = reset;
  assign EXU_io_pc = IDU_io_to_es_pc; // @[top.scala 77:12]
  assign EXU_io_ds_to_es_valid = IDU_io_ds_to_es_valid; // @[top.scala 78:24]
  assign EXU_io_ms_allowin = LSU_io_ms_allowin; // @[top.scala 79:20]
  assign EXU_io_ALUop = IDU_io_ALUop; // @[top.scala 80:15]
  assign EXU_io_src1_value = IDU_io_src1; // @[top.scala 81:20]
  assign EXU_io_src2_value = IDU_io_src2; // @[top.scala 82:20]
  assign EXU_io_rf_dst = IDU_io_rf_dst; // @[top.scala 83:16]
  assign EXU_io_store_data = IDU_io_store_data; // @[top.scala 84:20]
  assign EXU_io_load_type = IDU_io_load_type; // @[top.scala 86:19]
  assign EXU_io_ctrl_sign_reg_write = IDU_io_ctrl_sign_reg_write; // @[top.scala 85:19]
  assign EXU_io_ctrl_sign_Writemem_en = IDU_io_ctrl_sign_Writemem_en; // @[top.scala 85:19]
  assign EXU_io_ctrl_sign_Readmem_en = IDU_io_ctrl_sign_Readmem_en; // @[top.scala 85:19]
  assign EXU_io_ctrl_sign_Wmask = IDU_io_ctrl_sign_Wmask; // @[top.scala 85:19]
  assign LSU_clock = clock;
  assign LSU_reset = reset;
  assign LSU_io_pc = EXU_io_to_ms_pc; // @[top.scala 88:12]
  assign LSU_io_es_to_ms_valid = EXU_io_es_to_ms_valid; // @[top.scala 89:24]
  assign LSU_io_rf_we = EXU_io_to_ms_rf_we; // @[top.scala 91:15]
  assign LSU_io_rf_dst = EXU_io_to_ms_rf_dst; // @[top.scala 92:16]
  assign LSU_io_alu_res = EXU_io_to_ms_alures; // @[top.scala 93:17]
  assign LSU_io_store_data = EXU_io_to_ms_store_data; // @[top.scala 94:20]
  assign LSU_io_load_type = EXU_io_to_ms_load_type; // @[top.scala 99:19]
  assign LSU_io_wen = EXU_io_to_ms_wen; // @[top.scala 95:13]
  assign LSU_io_wstrb = EXU_io_to_ms_wstrb; // @[top.scala 96:15]
  assign LSU_io_ren = EXU_io_to_ms_ren; // @[top.scala 97:13]
  assign LSU_io_maddr = EXU_io_to_ms_maddr; // @[top.scala 98:15]
  assign LSU_io_axi_in_rdata = d_cache_io_to_lsu_rdata; // @[top.scala 34:16]
  assign LSU_io_axi_in_rvalid = d_cache_io_to_lsu_rvalid; // @[top.scala 34:16]
  assign LSU_io_axi_in_bvalid = d_cache_io_to_lsu_bvalid; // @[top.scala 34:16]
  assign WBU_clock = clock;
  assign WBU_reset = reset;
  assign WBU_io_pc = LSU_io_to_ws_pc; // @[top.scala 101:12]
  assign WBU_io_ms_to_ws_valid = LSU_io_ms_to_ws_valid; // @[top.scala 102:24]
  assign WBU_io_ms_final_res = LSU_io_ms_final_res; // @[top.scala 103:22]
  assign WBU_io_rf_we = LSU_io_to_ws_rf_we; // @[top.scala 104:15]
  assign WBU_io_rf_dst = LSU_io_to_ws_rf_dst; // @[top.scala 105:16]
  assign arbiter_clock = clock;
  assign arbiter_reset = reset;
  assign arbiter_io_ifu_axi_in_araddr = i_cache_io_to_axi_araddr; // @[top.scala 27:27]
  assign arbiter_io_ifu_axi_in_arlen = i_cache_io_to_axi_arlen; // @[top.scala 27:27]
  assign arbiter_io_ifu_axi_in_arvalid = i_cache_io_to_axi_arvalid; // @[top.scala 27:27]
  assign arbiter_io_ifu_axi_in_rready = i_cache_io_to_axi_rready; // @[top.scala 27:27]
  assign arbiter_io_lsu_axi_in_araddr = d_cache_io_to_axi_araddr; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_arlen = d_cache_io_to_axi_arlen; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_arvalid = d_cache_io_to_axi_arvalid; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_rready = d_cache_io_to_axi_rready; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_awaddr = d_cache_io_to_axi_awaddr; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_awlen = d_cache_io_to_axi_awlen; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_awvalid = d_cache_io_to_axi_awvalid; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_wdata = d_cache_io_to_axi_wdata; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_wstrb = d_cache_io_to_axi_wstrb; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_wvalid = d_cache_io_to_axi_wvalid; // @[top.scala 32:27]
  assign arbiter_io_lsu_axi_in_bready = d_cache_io_to_axi_bready; // @[top.scala 32:27]
  assign arbiter_io_axi_in_rdata = axi_io_axi_out_rdata; // @[top.scala 37:23]
  assign arbiter_io_axi_in_rlast = axi_io_axi_out_rlast; // @[top.scala 37:23]
  assign arbiter_io_axi_in_rvalid = axi_io_axi_out_rvalid; // @[top.scala 37:23]
  assign arbiter_io_axi_in_wready = axi_io_axi_out_wready; // @[top.scala 37:23]
  assign arbiter_io_axi_in_bvalid = axi_io_axi_out_bvalid; // @[top.scala 37:23]
  assign i_cache_clock = clock;
  assign i_cache_reset = reset;
  assign i_cache_io_from_ifu_araddr = IFU_io_axi_out_araddr; // @[top.scala 30:25]
  assign i_cache_io_from_ifu_arvalid = IFU_io_axi_out_arvalid; // @[top.scala 30:25]
  assign i_cache_io_from_ifu_rready = IFU_io_axi_out_rready; // @[top.scala 30:25]
  assign i_cache_io_from_axi_rdata = arbiter_io_ifu_axi_out_rdata; // @[top.scala 28:25]
  assign i_cache_io_from_axi_rlast = arbiter_io_ifu_axi_out_rlast; // @[top.scala 28:25]
  assign i_cache_io_from_axi_rvalid = arbiter_io_ifu_axi_out_rvalid; // @[top.scala 28:25]
  assign i_cache_io_clear_cache = IFU_io_clear_cache; // @[top.scala 50:28]
  assign d_cache_clock = clock;
  assign d_cache_reset = reset;
  assign d_cache_io_from_lsu_araddr = LSU_io_axi_out_araddr; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_arvalid = LSU_io_axi_out_arvalid; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_awaddr = LSU_io_axi_out_awaddr; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_awvalid = LSU_io_axi_out_awvalid; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_wdata = LSU_io_axi_out_wdata; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_wstrb = LSU_io_axi_out_wstrb; // @[top.scala 35:25]
  assign d_cache_io_from_lsu_wvalid = LSU_io_axi_out_wvalid; // @[top.scala 35:25]
  assign d_cache_io_from_axi_rdata = arbiter_io_lsu_axi_out_rdata; // @[top.scala 33:25]
  assign d_cache_io_from_axi_rlast = arbiter_io_lsu_axi_out_rlast; // @[top.scala 33:25]
  assign d_cache_io_from_axi_rvalid = arbiter_io_lsu_axi_out_rvalid; // @[top.scala 33:25]
  assign d_cache_io_from_axi_wready = arbiter_io_lsu_axi_out_wready; // @[top.scala 33:25]
  assign d_cache_io_from_axi_bvalid = arbiter_io_lsu_axi_out_bvalid; // @[top.scala 33:25]
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_axi_in_araddr = arbiter_io_axi_out_araddr; // @[top.scala 38:19]
  assign axi_io_axi_in_arlen = arbiter_io_axi_out_arlen; // @[top.scala 38:19]
  assign axi_io_axi_in_arvalid = arbiter_io_axi_out_arvalid; // @[top.scala 38:19]
  assign axi_io_axi_in_rready = arbiter_io_axi_out_rready; // @[top.scala 38:19]
  assign axi_io_axi_in_awaddr = arbiter_io_axi_out_awaddr; // @[top.scala 38:19]
  assign axi_io_axi_in_awlen = arbiter_io_axi_out_awlen; // @[top.scala 38:19]
  assign axi_io_axi_in_awvalid = arbiter_io_axi_out_awvalid; // @[top.scala 38:19]
  assign axi_io_axi_in_wdata = arbiter_io_axi_out_wdata; // @[top.scala 38:19]
  assign axi_io_axi_in_wstrb = arbiter_io_axi_out_wstrb; // @[top.scala 38:19]
  assign axi_io_axi_in_wvalid = arbiter_io_axi_out_wvalid; // @[top.scala 38:19]
  assign axi_io_axi_in_bready = arbiter_io_axi_out_bready; // @[top.scala 38:19]
  assign dpi_flag = {{31'd0}, IDU_io_ALUop == 32'h2}; // @[top.scala 117:17]
  assign dpi_ecall_flag = {{31'd0}, IDU_io_ALUop == 32'h3d}; // @[top.scala 118:23]
  assign dpi_pc = WBU_io_ws_valid ? WBU_io_ws_pc : _dpi_io_pc_T_2; // @[top.scala 119:21]
  always @(posedge clock) begin
    if (reset) begin // @[top.scala 113:28]
      diff_step <= 1'h0; // @[top.scala 113:28]
    end else begin
      diff_step <= WBU_io_ws_valid; // @[top.scala 114:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  diff_step = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
