module AXI(
  input         clock,
  input         reset,
  input  [31:0] io_axi_in_araddr,
  input         io_axi_in_arvalid,
  input         io_axi_in_rready,
  input  [31:0] io_axi_in_awaddr,
  input         io_axi_in_awvalid,
  input  [31:0] io_axi_in_wdata,
  input  [7:0]  io_axi_in_wstrb,
  input         io_axi_in_wvalid,
  input         io_axi_in_bready,
  output        io_axi_out_arready,
  output [63:0] io_axi_out_rdata,
  output        io_axi_out_rvalid,
  output        io_axi_out_awready,
  output        io_axi_out_wready,
  output        io_axi_out_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] Mem_modle_Raddr; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Rdata; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Waddr; // @[AXI.scala 26:27]
  wire [63:0] Mem_modle_Wdata; // @[AXI.scala 26:27]
  wire [7:0] Mem_modle_Wmask; // @[AXI.scala 26:27]
  wire  Mem_modle_Write_en; // @[AXI.scala 26:27]
  wire  Mem_modle_Read_en; // @[AXI.scala 26:27]
  reg  axi_awready; // @[AXI.scala 13:30]
  reg  axi_wready; // @[AXI.scala 14:29]
  reg  axi_bvalid; // @[AXI.scala 17:29]
  reg  axi_arready; // @[AXI.scala 19:30]
  reg  axi_rvalid; // @[AXI.scala 21:29]
  reg [2:0] state; // @[AXI.scala 24:24]
  wire  _GEN_1 = io_axi_in_arvalid ? 1'h0 : axi_arready; // @[AXI.scala 49:42 51:29 19:30]
  wire  _GEN_2 = io_axi_in_arvalid | axi_rvalid; // @[AXI.scala 49:42 52:28 21:29]
  wire  _GEN_4 = io_axi_in_awvalid & io_axi_in_wvalid ? 1'h0 : axi_awready; // @[AXI.scala 39:56 41:29 13:30]
  wire  _GEN_5 = io_axi_in_awvalid & io_axi_in_wvalid ? 1'h0 : axi_wready; // @[AXI.scala 39:56 42:28 14:29]
  wire  _GEN_6 = io_axi_in_awvalid & io_axi_in_wvalid | axi_bvalid; // @[AXI.scala 39:56 43:28 17:29]
  wire  _GEN_7 = io_axi_in_awvalid & io_axi_in_wvalid ? axi_arready : _GEN_1; // @[AXI.scala 19:30 39:56]
  wire  _GEN_11 = io_axi_in_bready | axi_awready; // @[AXI.scala 56:35 59:29 13:30]
  wire  _GEN_12 = io_axi_in_bready | axi_wready; // @[AXI.scala 56:35 60:28 14:29]
  wire [2:0] _GEN_13 = io_axi_in_rready ? 3'h0 : state; // @[AXI.scala 64:35 65:23 24:24]
  wire  _GEN_14 = io_axi_in_rready | axi_arready; // @[AXI.scala 64:35 66:29 19:30]
  wire  _GEN_15 = io_axi_in_rready ? 1'h0 : axi_rvalid; // @[AXI.scala 64:35 67:28 21:29]
  wire  _GEN_17 = 3'h4 == state ? _GEN_14 : axi_arready; // @[AXI.scala 37:18 19:30]
  wire  _GEN_21 = 3'h3 == state ? _GEN_11 : axi_awready; // @[AXI.scala 37:18 13:30]
  wire  _GEN_22 = 3'h3 == state ? _GEN_12 : axi_wready; // @[AXI.scala 37:18 14:29]
  wire  _GEN_23 = 3'h3 == state ? axi_arready : _GEN_17; // @[AXI.scala 37:18 19:30]
  wire  _GEN_26 = 3'h0 == state ? _GEN_4 : _GEN_21; // @[AXI.scala 37:18]
  wire  _GEN_27 = 3'h0 == state ? _GEN_5 : _GEN_22; // @[AXI.scala 37:18]
  wire  _GEN_29 = 3'h0 == state ? _GEN_7 : _GEN_23; // @[AXI.scala 37:18]
  MEM Mem_modle ( // @[AXI.scala 26:27]
    .Raddr(Mem_modle_Raddr),
    .Rdata(Mem_modle_Rdata),
    .Waddr(Mem_modle_Waddr),
    .Wdata(Mem_modle_Wdata),
    .Wmask(Mem_modle_Wmask),
    .Write_en(Mem_modle_Write_en),
    .Read_en(Mem_modle_Read_en)
  );
  assign io_axi_out_arready = axi_arready; // @[AXI.scala 71:24]
  assign io_axi_out_rdata = Mem_modle_Rdata; // @[AXI.scala 72:22]
  assign io_axi_out_rvalid = axi_rvalid; // @[AXI.scala 73:23]
  assign io_axi_out_awready = axi_awready; // @[AXI.scala 74:24]
  assign io_axi_out_wready = axi_wready; // @[AXI.scala 75:23]
  assign io_axi_out_bvalid = axi_bvalid; // @[AXI.scala 76:23]
  assign Mem_modle_Raddr = {32'h0,io_axi_in_araddr}; // @[Cat.scala 31:58]
  assign Mem_modle_Waddr = {{32'd0}, io_axi_in_awaddr}; // @[AXI.scala 28:24]
  assign Mem_modle_Wdata = {{32'd0}, io_axi_in_wdata}; // @[AXI.scala 29:24]
  assign Mem_modle_Wmask = io_axi_in_wstrb; // @[AXI.scala 30:24]
  assign Mem_modle_Write_en = axi_wready & io_axi_in_wvalid; // @[AXI.scala 31:48]
  assign Mem_modle_Read_en = axi_arready & io_axi_in_arvalid; // @[AXI.scala 32:48]
  always @(posedge clock) begin
    axi_awready <= reset | _GEN_26; // @[AXI.scala 13:{30,30}]
    axi_wready <= reset | _GEN_27; // @[AXI.scala 14:{29,29}]
    if (reset) begin // @[AXI.scala 17:29]
      axi_bvalid <= 1'h0; // @[AXI.scala 17:29]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      axi_bvalid <= _GEN_6;
    end else if (3'h3 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_bready) begin // @[AXI.scala 56:35]
        axi_bvalid <= 1'h0; // @[AXI.scala 58:28]
      end
    end
    axi_arready <= reset | _GEN_29; // @[AXI.scala 19:{30,30}]
    if (reset) begin // @[AXI.scala 21:29]
      axi_rvalid <= 1'h0; // @[AXI.scala 21:29]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      if (!(io_axi_in_awvalid & io_axi_in_wvalid)) begin // @[AXI.scala 39:56]
        axi_rvalid <= _GEN_2;
      end
    end else if (!(3'h3 == state)) begin // @[AXI.scala 37:18]
      if (3'h4 == state) begin // @[AXI.scala 37:18]
        axi_rvalid <= _GEN_15;
      end
    end
    if (reset) begin // @[AXI.scala 24:24]
      state <= 3'h0; // @[AXI.scala 24:24]
    end else if (3'h0 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_awvalid & io_axi_in_wvalid) begin // @[AXI.scala 39:56]
        state <= 3'h3; // @[AXI.scala 40:23]
      end else if (io_axi_in_arvalid) begin // @[AXI.scala 49:42]
        state <= 3'h4; // @[AXI.scala 50:23]
      end
    end else if (3'h3 == state) begin // @[AXI.scala 37:18]
      if (io_axi_in_bready) begin // @[AXI.scala 56:35]
        state <= 3'h0; // @[AXI.scala 57:23]
      end
    end else if (3'h4 == state) begin // @[AXI.scala 37:18]
      state <= _GEN_13;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_awready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_wready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_bvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  axi_arready = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  axi_rvalid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSU(
  input         clock,
  input         reset,
  input         io_inst_store,
  input         io_inst_load,
  input  [31:0] io_mem_addr,
  input  [63:0] io_mem_wdata,
  input  [7:0]  io_mem_wstrb,
  output [63:0] io_mem_rdata,
  input         io_axi_in_arready,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_awready,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [31:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  axi_arvalid; // @[LSU.scala 19:30]
  reg  axi_rready; // @[LSU.scala 22:29]
  reg  axi_awvalid; // @[LSU.scala 23:30]
  reg  axi_wvalid; // @[LSU.scala 24:29]
  reg  axi_bready; // @[LSU.scala 25:29]
  reg [1:0] state; // @[LSU.scala 28:24]
  wire  _GEN_1 = io_inst_store | axi_awvalid; // @[LSU.scala 36:38 38:29 23:30]
  wire  _GEN_2 = io_inst_store | axi_wvalid; // @[LSU.scala 36:38 39:28 24:29]
  wire  _GEN_3 = io_inst_store | axi_bready; // @[LSU.scala 36:38 40:28 25:29]
  wire  _GEN_5 = io_inst_load | axi_arvalid; // @[LSU.scala 32:31 34:29 19:30]
  wire  _GEN_6 = io_inst_load | axi_rready; // @[LSU.scala 32:31 35:28 22:29]
  wire  _GEN_9 = io_inst_load ? axi_bready : _GEN_3; // @[LSU.scala 25:29 32:31]
  wire  _GEN_11 = io_axi_in_bvalid ? 1'h0 : axi_bready; // @[LSU.scala 44:35 46:28 25:29]
  wire  _GEN_14 = io_axi_in_arready ? 1'h0 : axi_arvalid; // @[LSU.scala 56:36 57:29 19:30]
  wire [1:0] _GEN_15 = io_axi_in_rvalid ? 2'h0 : state; // @[LSU.scala 59:35 60:23 28:24]
  wire  _GEN_16 = io_axi_in_rvalid ? 1'h0 : axi_rready; // @[LSU.scala 59:35 61:28 22:29]
  wire  _GEN_19 = 2'h2 == state ? _GEN_16 : axi_rready; // @[LSU.scala 30:18 22:29]
  wire  _GEN_21 = 2'h1 == state ? _GEN_11 : axi_bready; // @[LSU.scala 30:18 25:29]
  wire  _GEN_25 = 2'h1 == state ? axi_rready : _GEN_19; // @[LSU.scala 30:18 22:29]
  wire  _GEN_28 = 2'h0 == state ? _GEN_6 : _GEN_25; // @[LSU.scala 30:18]
  wire  _GEN_31 = 2'h0 == state ? _GEN_9 : _GEN_21; // @[LSU.scala 30:18]
  assign io_mem_rdata = io_axi_in_rdata; // @[LSU.scala 72:18]
  assign io_axi_out_araddr = io_mem_addr; // @[LSU.scala 73:23]
  assign io_axi_out_arvalid = axi_arvalid; // @[LSU.scala 74:24]
  assign io_axi_out_rready = axi_rready; // @[LSU.scala 75:23]
  assign io_axi_out_awaddr = io_mem_addr; // @[LSU.scala 76:23]
  assign io_axi_out_awvalid = axi_awvalid; // @[LSU.scala 77:24]
  assign io_axi_out_wdata = io_mem_wdata[31:0]; // @[LSU.scala 78:22]
  assign io_axi_out_wstrb = io_mem_wstrb; // @[LSU.scala 79:22]
  assign io_axi_out_wvalid = axi_wvalid; // @[LSU.scala 80:23]
  assign io_axi_out_bready = axi_bready; // @[LSU.scala 81:23]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 19:30]
      axi_arvalid <= 1'h0; // @[LSU.scala 19:30]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      axi_arvalid <= _GEN_5;
    end else if (!(2'h1 == state)) begin // @[LSU.scala 30:18]
      if (2'h2 == state) begin // @[LSU.scala 30:18]
        axi_arvalid <= _GEN_14;
      end
    end
    axi_rready <= reset | _GEN_28; // @[LSU.scala 22:{29,29}]
    if (reset) begin // @[LSU.scala 23:30]
      axi_awvalid <= 1'h0; // @[LSU.scala 23:30]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (!(io_inst_load)) begin // @[LSU.scala 32:31]
        axi_awvalid <= _GEN_1;
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_awready) begin // @[LSU.scala 51:36]
        axi_awvalid <= 1'h0; // @[LSU.scala 52:29]
      end
    end
    if (reset) begin // @[LSU.scala 24:29]
      axi_wvalid <= 1'h0; // @[LSU.scala 24:29]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (!(io_inst_load)) begin // @[LSU.scala 32:31]
        axi_wvalid <= _GEN_2;
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_wready) begin // @[LSU.scala 48:35]
        axi_wvalid <= 1'h0; // @[LSU.scala 49:28]
      end
    end
    axi_bready <= reset | _GEN_31; // @[LSU.scala 25:{29,29}]
    if (reset) begin // @[LSU.scala 28:24]
      state <= 2'h0; // @[LSU.scala 28:24]
    end else if (2'h0 == state) begin // @[LSU.scala 30:18]
      if (io_inst_load) begin // @[LSU.scala 32:31]
        state <= 2'h2; // @[LSU.scala 33:23]
      end else if (io_inst_store) begin // @[LSU.scala 36:38]
        state <= 2'h1; // @[LSU.scala 37:23]
      end
    end else if (2'h1 == state) begin // @[LSU.scala 30:18]
      if (io_axi_in_bvalid) begin // @[LSU.scala 44:35]
        state <= 2'h0; // @[LSU.scala 45:23]
      end
    end else if (2'h2 == state) begin // @[LSU.scala 30:18]
      state <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_arvalid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  axi_rready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  axi_awvalid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  axi_wvalid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  axi_bready = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI_ARBITER(
  input         clock,
  input         reset,
  input  [31:0] io_ifu_axi_in_araddr,
  input         io_ifu_axi_in_arvalid,
  input         io_ifu_axi_in_rready,
  output [63:0] io_ifu_axi_out_rdata,
  output        io_ifu_axi_out_rvalid,
  input  [31:0] io_lsu_axi_in_araddr,
  input         io_lsu_axi_in_arvalid,
  input         io_lsu_axi_in_rready,
  input  [31:0] io_lsu_axi_in_awaddr,
  input         io_lsu_axi_in_awvalid,
  input  [31:0] io_lsu_axi_in_wdata,
  input  [7:0]  io_lsu_axi_in_wstrb,
  input         io_lsu_axi_in_wvalid,
  input         io_lsu_axi_in_bready,
  output        io_lsu_axi_out_arready,
  output [63:0] io_lsu_axi_out_rdata,
  output        io_lsu_axi_out_rvalid,
  output        io_lsu_axi_out_awready,
  output        io_lsu_axi_out_wready,
  output        io_lsu_axi_out_bvalid,
  input         io_axi_in_arready,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  input         io_axi_in_awready,
  input         io_axi_in_wready,
  input         io_axi_in_bvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready,
  output [31:0] io_axi_out_awaddr,
  output        io_axi_out_awvalid,
  output [31:0] io_axi_out_wdata,
  output [7:0]  io_axi_out_wstrb,
  output        io_axi_out_wvalid,
  output        io_axi_out_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[axi_arbiter.scala 18:24]
  wire  _T_1 = ~reset; // @[axi_arbiter.scala 38:11]
  wire [1:0] _GEN_0 = io_ifu_axi_in_arvalid ? 2'h1 : state; // @[axi_arbiter.scala 51:46 52:23 18:24]
  wire [31:0] _GEN_1 = io_ifu_axi_in_arvalid ? io_ifu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 51:46 53:28 57:28]
  wire  _GEN_3 = io_ifu_axi_in_arvalid & io_ifu_axi_in_rready; // @[axi_arbiter.scala 51:46 53:28 57:28]
  wire [63:0] _GEN_11 = io_ifu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 51:46 54:32 59:32]
  wire  _GEN_12 = io_ifu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 51:46 54:32 59:32]
  wire [31:0] _GEN_23 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_araddr : _GEN_1; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_24 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_arvalid : io_ifu_axi_in_arvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_25 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_rready : _GEN_3; // @[axi_arbiter.scala 46:46 48:28]
  wire [31:0] _GEN_26 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_27 = io_lsu_axi_in_arvalid & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire [31:0] _GEN_28 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wdata : 32'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire [7:0] _GEN_29 = io_lsu_axi_in_arvalid ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_30 = io_lsu_axi_in_arvalid & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_31 = io_lsu_axi_in_arvalid & io_lsu_axi_in_bready; // @[axi_arbiter.scala 46:46 48:28]
  wire  _GEN_32 = io_lsu_axi_in_arvalid & io_axi_in_arready; // @[axi_arbiter.scala 46:46 49:32]
  wire [63:0] _GEN_33 = io_lsu_axi_in_arvalid ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_34 = io_lsu_axi_in_arvalid & io_axi_in_rvalid; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_35 = io_lsu_axi_in_arvalid & io_axi_in_awready; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_36 = io_lsu_axi_in_arvalid & io_axi_in_wready; // @[axi_arbiter.scala 46:46 49:32]
  wire  _GEN_37 = io_lsu_axi_in_arvalid & io_axi_in_bvalid; // @[axi_arbiter.scala 46:46 49:32]
  wire [63:0] _GEN_39 = io_lsu_axi_in_arvalid ? 64'h0 : _GEN_11; // @[axi_arbiter.scala 46:46 50:32]
  wire  _GEN_40 = io_lsu_axi_in_arvalid ? 1'h0 : _GEN_12; // @[axi_arbiter.scala 46:46 50:32]
  wire [31:0] _GEN_45 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_araddr : _GEN_23; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_46 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_arvalid : _GEN_24; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_47 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_rready : _GEN_25; // @[axi_arbiter.scala 41:40 43:28]
  wire [31:0] _GEN_48 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awaddr : _GEN_26; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_49 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_awvalid : _GEN_27; // @[axi_arbiter.scala 41:40 43:28]
  wire [31:0] _GEN_50 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wdata : _GEN_28; // @[axi_arbiter.scala 41:40 43:28]
  wire [7:0] _GEN_51 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wstrb : _GEN_29; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_52 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_wvalid : _GEN_30; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_53 = io_lsu_axi_in_awvalid ? io_lsu_axi_in_bready : _GEN_31; // @[axi_arbiter.scala 41:40 43:28]
  wire  _GEN_54 = io_lsu_axi_in_awvalid ? io_axi_in_arready : _GEN_32; // @[axi_arbiter.scala 41:40 44:32]
  wire [63:0] _GEN_55 = io_lsu_axi_in_awvalid ? io_axi_in_rdata : _GEN_33; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_56 = io_lsu_axi_in_awvalid ? io_axi_in_rvalid : _GEN_34; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_57 = io_lsu_axi_in_awvalid ? io_axi_in_awready : _GEN_35; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_58 = io_lsu_axi_in_awvalid ? io_axi_in_wready : _GEN_36; // @[axi_arbiter.scala 41:40 44:32]
  wire  _GEN_59 = io_lsu_axi_in_awvalid ? io_axi_in_bvalid : _GEN_37; // @[axi_arbiter.scala 41:40 44:32]
  wire [63:0] _GEN_61 = io_lsu_axi_in_awvalid ? 64'h0 : _GEN_39; // @[axi_arbiter.scala 41:40 45:32]
  wire  _GEN_62 = io_lsu_axi_in_awvalid ? 1'h0 : _GEN_40; // @[axi_arbiter.scala 41:40 45:32]
  wire [1:0] _GEN_67 = io_lsu_axi_out_rvalid & io_lsu_axi_in_rready ? 2'h0 : state; // @[axi_arbiter.scala 74:64 75:23 18:24]
  wire [1:0] _GEN_68 = io_lsu_axi_out_bvalid & io_lsu_axi_in_bready ? 2'h0 : state; // @[axi_arbiter.scala 82:64 83:23 18:24]
  wire [31:0] _GEN_69 = state == 2'h3 ? io_lsu_axi_in_araddr : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_70 = state == 2'h3 & io_lsu_axi_in_arvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_71 = state == 2'h3 & io_lsu_axi_in_rready; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [31:0] _GEN_72 = state == 2'h3 ? io_lsu_axi_in_awaddr : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_73 = state == 2'h3 & io_lsu_axi_in_awvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [31:0] _GEN_74 = state == 2'h3 ? io_lsu_axi_in_wdata : 32'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire [7:0] _GEN_75 = state == 2'h3 ? io_lsu_axi_in_wstrb : 8'h0; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_76 = state == 2'h3 & io_lsu_axi_in_wvalid; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_77 = state == 2'h3 & io_lsu_axi_in_bready; // @[axi_arbiter.scala 78:39 79:24 87:24]
  wire  _GEN_78 = state == 2'h3 & io_axi_in_arready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire [63:0] _GEN_79 = state == 2'h3 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_80 = state == 2'h3 & io_axi_in_rvalid; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_81 = state == 2'h3 & io_axi_in_awready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_82 = state == 2'h3 & io_axi_in_wready; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire  _GEN_83 = state == 2'h3 & io_axi_in_bvalid; // @[axi_arbiter.scala 78:39 80:28 88:28]
  wire [1:0] _GEN_90 = state == 2'h3 ? _GEN_68 : state; // @[axi_arbiter.scala 18:24 78:39]
  wire [31:0] _GEN_91 = state == 2'h2 ? io_lsu_axi_in_araddr : _GEN_69; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_92 = state == 2'h2 ? io_lsu_axi_in_arvalid : _GEN_70; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_93 = state == 2'h2 ? io_lsu_axi_in_rready : _GEN_71; // @[axi_arbiter.scala 70:39 71:24]
  wire [31:0] _GEN_94 = state == 2'h2 ? io_lsu_axi_in_awaddr : _GEN_72; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_95 = state == 2'h2 ? io_lsu_axi_in_awvalid : _GEN_73; // @[axi_arbiter.scala 70:39 71:24]
  wire [31:0] _GEN_96 = state == 2'h2 ? io_lsu_axi_in_wdata : _GEN_74; // @[axi_arbiter.scala 70:39 71:24]
  wire [7:0] _GEN_97 = state == 2'h2 ? io_lsu_axi_in_wstrb : _GEN_75; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_98 = state == 2'h2 ? io_lsu_axi_in_wvalid : _GEN_76; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_99 = state == 2'h2 ? io_lsu_axi_in_bready : _GEN_77; // @[axi_arbiter.scala 70:39 71:24]
  wire  _GEN_100 = state == 2'h2 ? io_axi_in_arready : _GEN_78; // @[axi_arbiter.scala 70:39 72:28]
  wire [63:0] _GEN_101 = state == 2'h2 ? io_axi_in_rdata : _GEN_79; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_102 = state == 2'h2 ? io_axi_in_rvalid : _GEN_80; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_103 = state == 2'h2 ? io_axi_in_awready : _GEN_81; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_104 = state == 2'h2 ? io_axi_in_wready : _GEN_82; // @[axi_arbiter.scala 70:39 72:28]
  wire  _GEN_105 = state == 2'h2 ? io_axi_in_bvalid : _GEN_83; // @[axi_arbiter.scala 70:39 72:28]
  wire [31:0] _GEN_113 = state == 2'h1 ? io_ifu_axi_in_araddr : _GEN_91; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_114 = state == 2'h1 ? io_ifu_axi_in_arvalid : _GEN_92; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_115 = state == 2'h1 ? io_ifu_axi_in_rready : _GEN_93; // @[axi_arbiter.scala 62:39 63:24]
  wire [31:0] _GEN_116 = state == 2'h1 ? 32'h0 : _GEN_94; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_117 = state == 2'h1 ? 1'h0 : _GEN_95; // @[axi_arbiter.scala 62:39 63:24]
  wire [31:0] _GEN_118 = state == 2'h1 ? 32'h0 : _GEN_96; // @[axi_arbiter.scala 62:39 63:24]
  wire [7:0] _GEN_119 = state == 2'h1 ? 8'h0 : _GEN_97; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_120 = state == 2'h1 ? 1'h0 : _GEN_98; // @[axi_arbiter.scala 62:39 63:24]
  wire  _GEN_121 = state == 2'h1 ? 1'h0 : _GEN_99; // @[axi_arbiter.scala 62:39 63:24]
  wire [63:0] _GEN_123 = state == 2'h1 ? io_axi_in_rdata : 64'h0; // @[axi_arbiter.scala 62:39 64:28]
  wire  _GEN_124 = state == 2'h1 & io_axi_in_rvalid; // @[axi_arbiter.scala 62:39 64:28]
  wire  _GEN_128 = state == 2'h1 ? 1'h0 : _GEN_100; // @[axi_arbiter.scala 62:39 65:28]
  wire [63:0] _GEN_129 = state == 2'h1 ? 64'h0 : _GEN_101; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_130 = state == 2'h1 ? 1'h0 : _GEN_102; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_131 = state == 2'h1 ? 1'h0 : _GEN_103; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_132 = state == 2'h1 ? 1'h0 : _GEN_104; // @[axi_arbiter.scala 62:39 65:28]
  wire  _GEN_133 = state == 2'h1 ? 1'h0 : _GEN_105; // @[axi_arbiter.scala 62:39 65:28]
  assign io_ifu_axi_out_rdata = state == 2'h0 ? _GEN_61 : _GEN_123; // @[axi_arbiter.scala 40:27]
  assign io_ifu_axi_out_rvalid = state == 2'h0 ? _GEN_62 : _GEN_124; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_arready = state == 2'h0 ? _GEN_54 : _GEN_128; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_rdata = state == 2'h0 ? _GEN_55 : _GEN_129; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_rvalid = state == 2'h0 ? _GEN_56 : _GEN_130; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_awready = state == 2'h0 ? _GEN_57 : _GEN_131; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_wready = state == 2'h0 ? _GEN_58 : _GEN_132; // @[axi_arbiter.scala 40:27]
  assign io_lsu_axi_out_bvalid = state == 2'h0 ? _GEN_59 : _GEN_133; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_araddr = state == 2'h0 ? _GEN_45 : _GEN_113; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_arvalid = state == 2'h0 ? _GEN_46 : _GEN_114; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_rready = state == 2'h0 ? _GEN_47 : _GEN_115; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_awaddr = state == 2'h0 ? _GEN_48 : _GEN_116; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_awvalid = state == 2'h0 ? _GEN_49 : _GEN_117; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wdata = state == 2'h0 ? _GEN_50 : _GEN_118; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wstrb = state == 2'h0 ? _GEN_51 : _GEN_119; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_wvalid = state == 2'h0 ? _GEN_52 : _GEN_120; // @[axi_arbiter.scala 40:27]
  assign io_axi_out_bready = state == 2'h0 ? _GEN_53 : _GEN_121; // @[axi_arbiter.scala 40:27]
  always @(posedge clock) begin
    if (reset) begin // @[axi_arbiter.scala 18:24]
      state <= 2'h0; // @[axi_arbiter.scala 18:24]
    end else if (state == 2'h0) begin // @[axi_arbiter.scala 40:27]
      if (io_lsu_axi_in_awvalid) begin // @[axi_arbiter.scala 41:40]
        state <= 2'h3; // @[axi_arbiter.scala 42:23]
      end else if (io_lsu_axi_in_arvalid) begin // @[axi_arbiter.scala 46:46]
        state <= 2'h2; // @[axi_arbiter.scala 47:23]
      end else begin
        state <= _GEN_0;
      end
    end else if (state == 2'h1) begin // @[axi_arbiter.scala 62:39]
      if (io_ifu_axi_out_rvalid & io_ifu_axi_in_rready) begin // @[axi_arbiter.scala 66:64]
        state <= 2'h0; // @[axi_arbiter.scala 67:23]
      end
    end else if (state == 2'h2) begin // @[axi_arbiter.scala 70:39]
      state <= _GEN_67;
    end else begin
      state <= _GEN_90;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"arbiter state:%d\n",state); // @[axi_arbiter.scala 38:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"ifu_arvalid:%d lsu_awvalid:%d lsu_arvalid:%d\n",io_ifu_axi_in_arvalid,
            io_lsu_axi_in_awvalid,io_lsu_axi_in_arvalid); // @[axi_arbiter.scala 39:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU_AXI(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input         io_pc_valid,
  output        io_inst_valid,
  output [31:0] io_inst,
  output [31:0] io_inst_reg,
  input  [63:0] io_axi_in_rdata,
  input         io_axi_in_rvalid,
  output [31:0] io_axi_out_araddr,
  output        io_axi_out_arvalid,
  output        io_axi_out_rready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  inst_ready; // @[IFU_AXI.scala 19:29]
  wire  _GEN_0 = io_axi_in_rvalid & inst_ready ? 1'h0 : 1'h1; // @[IFU_AXI.scala 20:41 21:20 23:20]
  reg [31:0] inst_reg; // @[IFU_AXI.scala 25:27]
  assign io_inst_valid = io_axi_in_rvalid; // @[IFU_AXI.scala 41:19]
  assign io_inst = io_axi_in_rdata[31:0]; // @[IFU_AXI.scala 39:31]
  assign io_inst_reg = inst_reg; // @[IFU_AXI.scala 40:17]
  assign io_axi_out_araddr = io_pc[31:0]; // @[IFU_AXI.scala 29:31]
  assign io_axi_out_arvalid = io_pc_valid; // @[IFU_AXI.scala 30:24]
  assign io_axi_out_rready = inst_ready; // @[IFU_AXI.scala 31:23]
  always @(posedge clock) begin
    inst_ready <= reset | _GEN_0; // @[IFU_AXI.scala 19:{29,29}]
    if (reset) begin // @[IFU_AXI.scala 25:27]
      inst_reg <= 32'h0; // @[IFU_AXI.scala 25:27]
    end else if (io_axi_in_rvalid) begin // @[IFU_AXI.scala 26:27]
      inst_reg <= io_axi_in_rdata[31:0]; // @[IFU_AXI.scala 27:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst_ready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  inst_reg = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module I_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_ifu_araddr,
  input         io_from_ifu_arvalid,
  input         io_from_ifu_rready,
  output [63:0] io_to_ifu_rdata,
  output        io_to_ifu_rvalid,
  output [31:0] io_to_axi_araddr,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [63:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = ~reset; // @[cache.scala 14:11]
  reg [63:0] ram_0_0; // @[cache.scala 17:24]
  reg [63:0] ram_0_1; // @[cache.scala 17:24]
  reg [63:0] ram_0_2; // @[cache.scala 17:24]
  reg [63:0] ram_0_3; // @[cache.scala 17:24]
  reg [63:0] ram_0_4; // @[cache.scala 17:24]
  reg [63:0] ram_0_5; // @[cache.scala 17:24]
  reg [63:0] ram_0_6; // @[cache.scala 17:24]
  reg [63:0] ram_0_7; // @[cache.scala 17:24]
  reg [63:0] ram_0_8; // @[cache.scala 17:24]
  reg [63:0] ram_0_9; // @[cache.scala 17:24]
  reg [63:0] ram_0_10; // @[cache.scala 17:24]
  reg [63:0] ram_0_11; // @[cache.scala 17:24]
  reg [63:0] ram_0_12; // @[cache.scala 17:24]
  reg [63:0] ram_0_13; // @[cache.scala 17:24]
  reg [63:0] ram_0_14; // @[cache.scala 17:24]
  reg [63:0] ram_0_15; // @[cache.scala 17:24]
  reg [63:0] ram_0_16; // @[cache.scala 17:24]
  reg [63:0] ram_0_17; // @[cache.scala 17:24]
  reg [63:0] ram_0_18; // @[cache.scala 17:24]
  reg [63:0] ram_0_19; // @[cache.scala 17:24]
  reg [63:0] ram_0_20; // @[cache.scala 17:24]
  reg [63:0] ram_0_21; // @[cache.scala 17:24]
  reg [63:0] ram_0_22; // @[cache.scala 17:24]
  reg [63:0] ram_0_23; // @[cache.scala 17:24]
  reg [63:0] ram_0_24; // @[cache.scala 17:24]
  reg [63:0] ram_0_25; // @[cache.scala 17:24]
  reg [63:0] ram_0_26; // @[cache.scala 17:24]
  reg [63:0] ram_0_27; // @[cache.scala 17:24]
  reg [63:0] ram_0_28; // @[cache.scala 17:24]
  reg [63:0] ram_0_29; // @[cache.scala 17:24]
  reg [63:0] ram_0_30; // @[cache.scala 17:24]
  reg [63:0] ram_0_31; // @[cache.scala 17:24]
  reg [63:0] ram_0_32; // @[cache.scala 17:24]
  reg [63:0] ram_0_33; // @[cache.scala 17:24]
  reg [63:0] ram_0_34; // @[cache.scala 17:24]
  reg [63:0] ram_0_35; // @[cache.scala 17:24]
  reg [63:0] ram_0_36; // @[cache.scala 17:24]
  reg [63:0] ram_0_37; // @[cache.scala 17:24]
  reg [63:0] ram_0_38; // @[cache.scala 17:24]
  reg [63:0] ram_0_39; // @[cache.scala 17:24]
  reg [63:0] ram_0_40; // @[cache.scala 17:24]
  reg [63:0] ram_0_41; // @[cache.scala 17:24]
  reg [63:0] ram_0_42; // @[cache.scala 17:24]
  reg [63:0] ram_0_43; // @[cache.scala 17:24]
  reg [63:0] ram_0_44; // @[cache.scala 17:24]
  reg [63:0] ram_0_45; // @[cache.scala 17:24]
  reg [63:0] ram_0_46; // @[cache.scala 17:24]
  reg [63:0] ram_0_47; // @[cache.scala 17:24]
  reg [63:0] ram_0_48; // @[cache.scala 17:24]
  reg [63:0] ram_0_49; // @[cache.scala 17:24]
  reg [63:0] ram_0_50; // @[cache.scala 17:24]
  reg [63:0] ram_0_51; // @[cache.scala 17:24]
  reg [63:0] ram_0_52; // @[cache.scala 17:24]
  reg [63:0] ram_0_53; // @[cache.scala 17:24]
  reg [63:0] ram_0_54; // @[cache.scala 17:24]
  reg [63:0] ram_0_55; // @[cache.scala 17:24]
  reg [63:0] ram_0_56; // @[cache.scala 17:24]
  reg [63:0] ram_0_57; // @[cache.scala 17:24]
  reg [63:0] ram_0_58; // @[cache.scala 17:24]
  reg [63:0] ram_0_59; // @[cache.scala 17:24]
  reg [63:0] ram_0_60; // @[cache.scala 17:24]
  reg [63:0] ram_0_61; // @[cache.scala 17:24]
  reg [63:0] ram_0_62; // @[cache.scala 17:24]
  reg [63:0] ram_0_63; // @[cache.scala 17:24]
  reg [63:0] ram_0_64; // @[cache.scala 17:24]
  reg [63:0] ram_0_65; // @[cache.scala 17:24]
  reg [63:0] ram_0_66; // @[cache.scala 17:24]
  reg [63:0] ram_0_67; // @[cache.scala 17:24]
  reg [63:0] ram_0_68; // @[cache.scala 17:24]
  reg [63:0] ram_0_69; // @[cache.scala 17:24]
  reg [63:0] ram_0_70; // @[cache.scala 17:24]
  reg [63:0] ram_0_71; // @[cache.scala 17:24]
  reg [63:0] ram_0_72; // @[cache.scala 17:24]
  reg [63:0] ram_0_73; // @[cache.scala 17:24]
  reg [63:0] ram_0_74; // @[cache.scala 17:24]
  reg [63:0] ram_0_75; // @[cache.scala 17:24]
  reg [63:0] ram_0_76; // @[cache.scala 17:24]
  reg [63:0] ram_0_77; // @[cache.scala 17:24]
  reg [63:0] ram_0_78; // @[cache.scala 17:24]
  reg [63:0] ram_0_79; // @[cache.scala 17:24]
  reg [63:0] ram_0_80; // @[cache.scala 17:24]
  reg [63:0] ram_0_81; // @[cache.scala 17:24]
  reg [63:0] ram_0_82; // @[cache.scala 17:24]
  reg [63:0] ram_0_83; // @[cache.scala 17:24]
  reg [63:0] ram_0_84; // @[cache.scala 17:24]
  reg [63:0] ram_0_85; // @[cache.scala 17:24]
  reg [63:0] ram_0_86; // @[cache.scala 17:24]
  reg [63:0] ram_0_87; // @[cache.scala 17:24]
  reg [63:0] ram_0_88; // @[cache.scala 17:24]
  reg [63:0] ram_0_89; // @[cache.scala 17:24]
  reg [63:0] ram_0_90; // @[cache.scala 17:24]
  reg [63:0] ram_0_91; // @[cache.scala 17:24]
  reg [63:0] ram_0_92; // @[cache.scala 17:24]
  reg [63:0] ram_0_93; // @[cache.scala 17:24]
  reg [63:0] ram_0_94; // @[cache.scala 17:24]
  reg [63:0] ram_0_95; // @[cache.scala 17:24]
  reg [63:0] ram_0_96; // @[cache.scala 17:24]
  reg [63:0] ram_0_97; // @[cache.scala 17:24]
  reg [63:0] ram_0_98; // @[cache.scala 17:24]
  reg [63:0] ram_0_99; // @[cache.scala 17:24]
  reg [63:0] ram_0_100; // @[cache.scala 17:24]
  reg [63:0] ram_0_101; // @[cache.scala 17:24]
  reg [63:0] ram_0_102; // @[cache.scala 17:24]
  reg [63:0] ram_0_103; // @[cache.scala 17:24]
  reg [63:0] ram_0_104; // @[cache.scala 17:24]
  reg [63:0] ram_0_105; // @[cache.scala 17:24]
  reg [63:0] ram_0_106; // @[cache.scala 17:24]
  reg [63:0] ram_0_107; // @[cache.scala 17:24]
  reg [63:0] ram_0_108; // @[cache.scala 17:24]
  reg [63:0] ram_0_109; // @[cache.scala 17:24]
  reg [63:0] ram_0_110; // @[cache.scala 17:24]
  reg [63:0] ram_0_111; // @[cache.scala 17:24]
  reg [63:0] ram_0_112; // @[cache.scala 17:24]
  reg [63:0] ram_0_113; // @[cache.scala 17:24]
  reg [63:0] ram_0_114; // @[cache.scala 17:24]
  reg [63:0] ram_0_115; // @[cache.scala 17:24]
  reg [63:0] ram_0_116; // @[cache.scala 17:24]
  reg [63:0] ram_0_117; // @[cache.scala 17:24]
  reg [63:0] ram_0_118; // @[cache.scala 17:24]
  reg [63:0] ram_0_119; // @[cache.scala 17:24]
  reg [63:0] ram_0_120; // @[cache.scala 17:24]
  reg [63:0] ram_0_121; // @[cache.scala 17:24]
  reg [63:0] ram_0_122; // @[cache.scala 17:24]
  reg [63:0] ram_0_123; // @[cache.scala 17:24]
  reg [63:0] ram_0_124; // @[cache.scala 17:24]
  reg [63:0] ram_0_125; // @[cache.scala 17:24]
  reg [63:0] ram_0_126; // @[cache.scala 17:24]
  reg [63:0] ram_0_127; // @[cache.scala 17:24]
  reg [63:0] ram_1_0; // @[cache.scala 18:24]
  reg [63:0] ram_1_1; // @[cache.scala 18:24]
  reg [63:0] ram_1_2; // @[cache.scala 18:24]
  reg [63:0] ram_1_3; // @[cache.scala 18:24]
  reg [63:0] ram_1_4; // @[cache.scala 18:24]
  reg [63:0] ram_1_5; // @[cache.scala 18:24]
  reg [63:0] ram_1_6; // @[cache.scala 18:24]
  reg [63:0] ram_1_7; // @[cache.scala 18:24]
  reg [63:0] ram_1_8; // @[cache.scala 18:24]
  reg [63:0] ram_1_9; // @[cache.scala 18:24]
  reg [63:0] ram_1_10; // @[cache.scala 18:24]
  reg [63:0] ram_1_11; // @[cache.scala 18:24]
  reg [63:0] ram_1_12; // @[cache.scala 18:24]
  reg [63:0] ram_1_13; // @[cache.scala 18:24]
  reg [63:0] ram_1_14; // @[cache.scala 18:24]
  reg [63:0] ram_1_15; // @[cache.scala 18:24]
  reg [63:0] ram_1_16; // @[cache.scala 18:24]
  reg [63:0] ram_1_17; // @[cache.scala 18:24]
  reg [63:0] ram_1_18; // @[cache.scala 18:24]
  reg [63:0] ram_1_19; // @[cache.scala 18:24]
  reg [63:0] ram_1_20; // @[cache.scala 18:24]
  reg [63:0] ram_1_21; // @[cache.scala 18:24]
  reg [63:0] ram_1_22; // @[cache.scala 18:24]
  reg [63:0] ram_1_23; // @[cache.scala 18:24]
  reg [63:0] ram_1_24; // @[cache.scala 18:24]
  reg [63:0] ram_1_25; // @[cache.scala 18:24]
  reg [63:0] ram_1_26; // @[cache.scala 18:24]
  reg [63:0] ram_1_27; // @[cache.scala 18:24]
  reg [63:0] ram_1_28; // @[cache.scala 18:24]
  reg [63:0] ram_1_29; // @[cache.scala 18:24]
  reg [63:0] ram_1_30; // @[cache.scala 18:24]
  reg [63:0] ram_1_31; // @[cache.scala 18:24]
  reg [63:0] ram_1_32; // @[cache.scala 18:24]
  reg [63:0] ram_1_33; // @[cache.scala 18:24]
  reg [63:0] ram_1_34; // @[cache.scala 18:24]
  reg [63:0] ram_1_35; // @[cache.scala 18:24]
  reg [63:0] ram_1_36; // @[cache.scala 18:24]
  reg [63:0] ram_1_37; // @[cache.scala 18:24]
  reg [63:0] ram_1_38; // @[cache.scala 18:24]
  reg [63:0] ram_1_39; // @[cache.scala 18:24]
  reg [63:0] ram_1_40; // @[cache.scala 18:24]
  reg [63:0] ram_1_41; // @[cache.scala 18:24]
  reg [63:0] ram_1_42; // @[cache.scala 18:24]
  reg [63:0] ram_1_43; // @[cache.scala 18:24]
  reg [63:0] ram_1_44; // @[cache.scala 18:24]
  reg [63:0] ram_1_45; // @[cache.scala 18:24]
  reg [63:0] ram_1_46; // @[cache.scala 18:24]
  reg [63:0] ram_1_47; // @[cache.scala 18:24]
  reg [63:0] ram_1_48; // @[cache.scala 18:24]
  reg [63:0] ram_1_49; // @[cache.scala 18:24]
  reg [63:0] ram_1_50; // @[cache.scala 18:24]
  reg [63:0] ram_1_51; // @[cache.scala 18:24]
  reg [63:0] ram_1_52; // @[cache.scala 18:24]
  reg [63:0] ram_1_53; // @[cache.scala 18:24]
  reg [63:0] ram_1_54; // @[cache.scala 18:24]
  reg [63:0] ram_1_55; // @[cache.scala 18:24]
  reg [63:0] ram_1_56; // @[cache.scala 18:24]
  reg [63:0] ram_1_57; // @[cache.scala 18:24]
  reg [63:0] ram_1_58; // @[cache.scala 18:24]
  reg [63:0] ram_1_59; // @[cache.scala 18:24]
  reg [63:0] ram_1_60; // @[cache.scala 18:24]
  reg [63:0] ram_1_61; // @[cache.scala 18:24]
  reg [63:0] ram_1_62; // @[cache.scala 18:24]
  reg [63:0] ram_1_63; // @[cache.scala 18:24]
  reg [63:0] ram_1_64; // @[cache.scala 18:24]
  reg [63:0] ram_1_65; // @[cache.scala 18:24]
  reg [63:0] ram_1_66; // @[cache.scala 18:24]
  reg [63:0] ram_1_67; // @[cache.scala 18:24]
  reg [63:0] ram_1_68; // @[cache.scala 18:24]
  reg [63:0] ram_1_69; // @[cache.scala 18:24]
  reg [63:0] ram_1_70; // @[cache.scala 18:24]
  reg [63:0] ram_1_71; // @[cache.scala 18:24]
  reg [63:0] ram_1_72; // @[cache.scala 18:24]
  reg [63:0] ram_1_73; // @[cache.scala 18:24]
  reg [63:0] ram_1_74; // @[cache.scala 18:24]
  reg [63:0] ram_1_75; // @[cache.scala 18:24]
  reg [63:0] ram_1_76; // @[cache.scala 18:24]
  reg [63:0] ram_1_77; // @[cache.scala 18:24]
  reg [63:0] ram_1_78; // @[cache.scala 18:24]
  reg [63:0] ram_1_79; // @[cache.scala 18:24]
  reg [63:0] ram_1_80; // @[cache.scala 18:24]
  reg [63:0] ram_1_81; // @[cache.scala 18:24]
  reg [63:0] ram_1_82; // @[cache.scala 18:24]
  reg [63:0] ram_1_83; // @[cache.scala 18:24]
  reg [63:0] ram_1_84; // @[cache.scala 18:24]
  reg [63:0] ram_1_85; // @[cache.scala 18:24]
  reg [63:0] ram_1_86; // @[cache.scala 18:24]
  reg [63:0] ram_1_87; // @[cache.scala 18:24]
  reg [63:0] ram_1_88; // @[cache.scala 18:24]
  reg [63:0] ram_1_89; // @[cache.scala 18:24]
  reg [63:0] ram_1_90; // @[cache.scala 18:24]
  reg [63:0] ram_1_91; // @[cache.scala 18:24]
  reg [63:0] ram_1_92; // @[cache.scala 18:24]
  reg [63:0] ram_1_93; // @[cache.scala 18:24]
  reg [63:0] ram_1_94; // @[cache.scala 18:24]
  reg [63:0] ram_1_95; // @[cache.scala 18:24]
  reg [63:0] ram_1_96; // @[cache.scala 18:24]
  reg [63:0] ram_1_97; // @[cache.scala 18:24]
  reg [63:0] ram_1_98; // @[cache.scala 18:24]
  reg [63:0] ram_1_99; // @[cache.scala 18:24]
  reg [63:0] ram_1_100; // @[cache.scala 18:24]
  reg [63:0] ram_1_101; // @[cache.scala 18:24]
  reg [63:0] ram_1_102; // @[cache.scala 18:24]
  reg [63:0] ram_1_103; // @[cache.scala 18:24]
  reg [63:0] ram_1_104; // @[cache.scala 18:24]
  reg [63:0] ram_1_105; // @[cache.scala 18:24]
  reg [63:0] ram_1_106; // @[cache.scala 18:24]
  reg [63:0] ram_1_107; // @[cache.scala 18:24]
  reg [63:0] ram_1_108; // @[cache.scala 18:24]
  reg [63:0] ram_1_109; // @[cache.scala 18:24]
  reg [63:0] ram_1_110; // @[cache.scala 18:24]
  reg [63:0] ram_1_111; // @[cache.scala 18:24]
  reg [63:0] ram_1_112; // @[cache.scala 18:24]
  reg [63:0] ram_1_113; // @[cache.scala 18:24]
  reg [63:0] ram_1_114; // @[cache.scala 18:24]
  reg [63:0] ram_1_115; // @[cache.scala 18:24]
  reg [63:0] ram_1_116; // @[cache.scala 18:24]
  reg [63:0] ram_1_117; // @[cache.scala 18:24]
  reg [63:0] ram_1_118; // @[cache.scala 18:24]
  reg [63:0] ram_1_119; // @[cache.scala 18:24]
  reg [63:0] ram_1_120; // @[cache.scala 18:24]
  reg [63:0] ram_1_121; // @[cache.scala 18:24]
  reg [63:0] ram_1_122; // @[cache.scala 18:24]
  reg [63:0] ram_1_123; // @[cache.scala 18:24]
  reg [63:0] ram_1_124; // @[cache.scala 18:24]
  reg [63:0] ram_1_125; // @[cache.scala 18:24]
  reg [63:0] ram_1_126; // @[cache.scala 18:24]
  reg [63:0] ram_1_127; // @[cache.scala 18:24]
  reg [31:0] tag_0_0; // @[cache.scala 19:24]
  reg [31:0] tag_0_1; // @[cache.scala 19:24]
  reg [31:0] tag_0_2; // @[cache.scala 19:24]
  reg [31:0] tag_0_3; // @[cache.scala 19:24]
  reg [31:0] tag_0_4; // @[cache.scala 19:24]
  reg [31:0] tag_0_5; // @[cache.scala 19:24]
  reg [31:0] tag_0_6; // @[cache.scala 19:24]
  reg [31:0] tag_0_7; // @[cache.scala 19:24]
  reg [31:0] tag_0_8; // @[cache.scala 19:24]
  reg [31:0] tag_0_9; // @[cache.scala 19:24]
  reg [31:0] tag_0_10; // @[cache.scala 19:24]
  reg [31:0] tag_0_11; // @[cache.scala 19:24]
  reg [31:0] tag_0_12; // @[cache.scala 19:24]
  reg [31:0] tag_0_13; // @[cache.scala 19:24]
  reg [31:0] tag_0_14; // @[cache.scala 19:24]
  reg [31:0] tag_0_15; // @[cache.scala 19:24]
  reg [31:0] tag_0_16; // @[cache.scala 19:24]
  reg [31:0] tag_0_17; // @[cache.scala 19:24]
  reg [31:0] tag_0_18; // @[cache.scala 19:24]
  reg [31:0] tag_0_19; // @[cache.scala 19:24]
  reg [31:0] tag_0_20; // @[cache.scala 19:24]
  reg [31:0] tag_0_21; // @[cache.scala 19:24]
  reg [31:0] tag_0_22; // @[cache.scala 19:24]
  reg [31:0] tag_0_23; // @[cache.scala 19:24]
  reg [31:0] tag_0_24; // @[cache.scala 19:24]
  reg [31:0] tag_0_25; // @[cache.scala 19:24]
  reg [31:0] tag_0_26; // @[cache.scala 19:24]
  reg [31:0] tag_0_27; // @[cache.scala 19:24]
  reg [31:0] tag_0_28; // @[cache.scala 19:24]
  reg [31:0] tag_0_29; // @[cache.scala 19:24]
  reg [31:0] tag_0_30; // @[cache.scala 19:24]
  reg [31:0] tag_0_31; // @[cache.scala 19:24]
  reg [31:0] tag_0_32; // @[cache.scala 19:24]
  reg [31:0] tag_0_33; // @[cache.scala 19:24]
  reg [31:0] tag_0_34; // @[cache.scala 19:24]
  reg [31:0] tag_0_35; // @[cache.scala 19:24]
  reg [31:0] tag_0_36; // @[cache.scala 19:24]
  reg [31:0] tag_0_37; // @[cache.scala 19:24]
  reg [31:0] tag_0_38; // @[cache.scala 19:24]
  reg [31:0] tag_0_39; // @[cache.scala 19:24]
  reg [31:0] tag_0_40; // @[cache.scala 19:24]
  reg [31:0] tag_0_41; // @[cache.scala 19:24]
  reg [31:0] tag_0_42; // @[cache.scala 19:24]
  reg [31:0] tag_0_43; // @[cache.scala 19:24]
  reg [31:0] tag_0_44; // @[cache.scala 19:24]
  reg [31:0] tag_0_45; // @[cache.scala 19:24]
  reg [31:0] tag_0_46; // @[cache.scala 19:24]
  reg [31:0] tag_0_47; // @[cache.scala 19:24]
  reg [31:0] tag_0_48; // @[cache.scala 19:24]
  reg [31:0] tag_0_49; // @[cache.scala 19:24]
  reg [31:0] tag_0_50; // @[cache.scala 19:24]
  reg [31:0] tag_0_51; // @[cache.scala 19:24]
  reg [31:0] tag_0_52; // @[cache.scala 19:24]
  reg [31:0] tag_0_53; // @[cache.scala 19:24]
  reg [31:0] tag_0_54; // @[cache.scala 19:24]
  reg [31:0] tag_0_55; // @[cache.scala 19:24]
  reg [31:0] tag_0_56; // @[cache.scala 19:24]
  reg [31:0] tag_0_57; // @[cache.scala 19:24]
  reg [31:0] tag_0_58; // @[cache.scala 19:24]
  reg [31:0] tag_0_59; // @[cache.scala 19:24]
  reg [31:0] tag_0_60; // @[cache.scala 19:24]
  reg [31:0] tag_0_61; // @[cache.scala 19:24]
  reg [31:0] tag_0_62; // @[cache.scala 19:24]
  reg [31:0] tag_0_63; // @[cache.scala 19:24]
  reg [31:0] tag_0_64; // @[cache.scala 19:24]
  reg [31:0] tag_0_65; // @[cache.scala 19:24]
  reg [31:0] tag_0_66; // @[cache.scala 19:24]
  reg [31:0] tag_0_67; // @[cache.scala 19:24]
  reg [31:0] tag_0_68; // @[cache.scala 19:24]
  reg [31:0] tag_0_69; // @[cache.scala 19:24]
  reg [31:0] tag_0_70; // @[cache.scala 19:24]
  reg [31:0] tag_0_71; // @[cache.scala 19:24]
  reg [31:0] tag_0_72; // @[cache.scala 19:24]
  reg [31:0] tag_0_73; // @[cache.scala 19:24]
  reg [31:0] tag_0_74; // @[cache.scala 19:24]
  reg [31:0] tag_0_75; // @[cache.scala 19:24]
  reg [31:0] tag_0_76; // @[cache.scala 19:24]
  reg [31:0] tag_0_77; // @[cache.scala 19:24]
  reg [31:0] tag_0_78; // @[cache.scala 19:24]
  reg [31:0] tag_0_79; // @[cache.scala 19:24]
  reg [31:0] tag_0_80; // @[cache.scala 19:24]
  reg [31:0] tag_0_81; // @[cache.scala 19:24]
  reg [31:0] tag_0_82; // @[cache.scala 19:24]
  reg [31:0] tag_0_83; // @[cache.scala 19:24]
  reg [31:0] tag_0_84; // @[cache.scala 19:24]
  reg [31:0] tag_0_85; // @[cache.scala 19:24]
  reg [31:0] tag_0_86; // @[cache.scala 19:24]
  reg [31:0] tag_0_87; // @[cache.scala 19:24]
  reg [31:0] tag_0_88; // @[cache.scala 19:24]
  reg [31:0] tag_0_89; // @[cache.scala 19:24]
  reg [31:0] tag_0_90; // @[cache.scala 19:24]
  reg [31:0] tag_0_91; // @[cache.scala 19:24]
  reg [31:0] tag_0_92; // @[cache.scala 19:24]
  reg [31:0] tag_0_93; // @[cache.scala 19:24]
  reg [31:0] tag_0_94; // @[cache.scala 19:24]
  reg [31:0] tag_0_95; // @[cache.scala 19:24]
  reg [31:0] tag_0_96; // @[cache.scala 19:24]
  reg [31:0] tag_0_97; // @[cache.scala 19:24]
  reg [31:0] tag_0_98; // @[cache.scala 19:24]
  reg [31:0] tag_0_99; // @[cache.scala 19:24]
  reg [31:0] tag_0_100; // @[cache.scala 19:24]
  reg [31:0] tag_0_101; // @[cache.scala 19:24]
  reg [31:0] tag_0_102; // @[cache.scala 19:24]
  reg [31:0] tag_0_103; // @[cache.scala 19:24]
  reg [31:0] tag_0_104; // @[cache.scala 19:24]
  reg [31:0] tag_0_105; // @[cache.scala 19:24]
  reg [31:0] tag_0_106; // @[cache.scala 19:24]
  reg [31:0] tag_0_107; // @[cache.scala 19:24]
  reg [31:0] tag_0_108; // @[cache.scala 19:24]
  reg [31:0] tag_0_109; // @[cache.scala 19:24]
  reg [31:0] tag_0_110; // @[cache.scala 19:24]
  reg [31:0] tag_0_111; // @[cache.scala 19:24]
  reg [31:0] tag_0_112; // @[cache.scala 19:24]
  reg [31:0] tag_0_113; // @[cache.scala 19:24]
  reg [31:0] tag_0_114; // @[cache.scala 19:24]
  reg [31:0] tag_0_115; // @[cache.scala 19:24]
  reg [31:0] tag_0_116; // @[cache.scala 19:24]
  reg [31:0] tag_0_117; // @[cache.scala 19:24]
  reg [31:0] tag_0_118; // @[cache.scala 19:24]
  reg [31:0] tag_0_119; // @[cache.scala 19:24]
  reg [31:0] tag_0_120; // @[cache.scala 19:24]
  reg [31:0] tag_0_121; // @[cache.scala 19:24]
  reg [31:0] tag_0_122; // @[cache.scala 19:24]
  reg [31:0] tag_0_123; // @[cache.scala 19:24]
  reg [31:0] tag_0_124; // @[cache.scala 19:24]
  reg [31:0] tag_0_125; // @[cache.scala 19:24]
  reg [31:0] tag_0_126; // @[cache.scala 19:24]
  reg [31:0] tag_0_127; // @[cache.scala 19:24]
  reg [31:0] tag_1_0; // @[cache.scala 20:24]
  reg [31:0] tag_1_1; // @[cache.scala 20:24]
  reg [31:0] tag_1_2; // @[cache.scala 20:24]
  reg [31:0] tag_1_3; // @[cache.scala 20:24]
  reg [31:0] tag_1_4; // @[cache.scala 20:24]
  reg [31:0] tag_1_5; // @[cache.scala 20:24]
  reg [31:0] tag_1_6; // @[cache.scala 20:24]
  reg [31:0] tag_1_7; // @[cache.scala 20:24]
  reg [31:0] tag_1_8; // @[cache.scala 20:24]
  reg [31:0] tag_1_9; // @[cache.scala 20:24]
  reg [31:0] tag_1_10; // @[cache.scala 20:24]
  reg [31:0] tag_1_11; // @[cache.scala 20:24]
  reg [31:0] tag_1_12; // @[cache.scala 20:24]
  reg [31:0] tag_1_13; // @[cache.scala 20:24]
  reg [31:0] tag_1_14; // @[cache.scala 20:24]
  reg [31:0] tag_1_15; // @[cache.scala 20:24]
  reg [31:0] tag_1_16; // @[cache.scala 20:24]
  reg [31:0] tag_1_17; // @[cache.scala 20:24]
  reg [31:0] tag_1_18; // @[cache.scala 20:24]
  reg [31:0] tag_1_19; // @[cache.scala 20:24]
  reg [31:0] tag_1_20; // @[cache.scala 20:24]
  reg [31:0] tag_1_21; // @[cache.scala 20:24]
  reg [31:0] tag_1_22; // @[cache.scala 20:24]
  reg [31:0] tag_1_23; // @[cache.scala 20:24]
  reg [31:0] tag_1_24; // @[cache.scala 20:24]
  reg [31:0] tag_1_25; // @[cache.scala 20:24]
  reg [31:0] tag_1_26; // @[cache.scala 20:24]
  reg [31:0] tag_1_27; // @[cache.scala 20:24]
  reg [31:0] tag_1_28; // @[cache.scala 20:24]
  reg [31:0] tag_1_29; // @[cache.scala 20:24]
  reg [31:0] tag_1_30; // @[cache.scala 20:24]
  reg [31:0] tag_1_31; // @[cache.scala 20:24]
  reg [31:0] tag_1_32; // @[cache.scala 20:24]
  reg [31:0] tag_1_33; // @[cache.scala 20:24]
  reg [31:0] tag_1_34; // @[cache.scala 20:24]
  reg [31:0] tag_1_35; // @[cache.scala 20:24]
  reg [31:0] tag_1_36; // @[cache.scala 20:24]
  reg [31:0] tag_1_37; // @[cache.scala 20:24]
  reg [31:0] tag_1_38; // @[cache.scala 20:24]
  reg [31:0] tag_1_39; // @[cache.scala 20:24]
  reg [31:0] tag_1_40; // @[cache.scala 20:24]
  reg [31:0] tag_1_41; // @[cache.scala 20:24]
  reg [31:0] tag_1_42; // @[cache.scala 20:24]
  reg [31:0] tag_1_43; // @[cache.scala 20:24]
  reg [31:0] tag_1_44; // @[cache.scala 20:24]
  reg [31:0] tag_1_45; // @[cache.scala 20:24]
  reg [31:0] tag_1_46; // @[cache.scala 20:24]
  reg [31:0] tag_1_47; // @[cache.scala 20:24]
  reg [31:0] tag_1_48; // @[cache.scala 20:24]
  reg [31:0] tag_1_49; // @[cache.scala 20:24]
  reg [31:0] tag_1_50; // @[cache.scala 20:24]
  reg [31:0] tag_1_51; // @[cache.scala 20:24]
  reg [31:0] tag_1_52; // @[cache.scala 20:24]
  reg [31:0] tag_1_53; // @[cache.scala 20:24]
  reg [31:0] tag_1_54; // @[cache.scala 20:24]
  reg [31:0] tag_1_55; // @[cache.scala 20:24]
  reg [31:0] tag_1_56; // @[cache.scala 20:24]
  reg [31:0] tag_1_57; // @[cache.scala 20:24]
  reg [31:0] tag_1_58; // @[cache.scala 20:24]
  reg [31:0] tag_1_59; // @[cache.scala 20:24]
  reg [31:0] tag_1_60; // @[cache.scala 20:24]
  reg [31:0] tag_1_61; // @[cache.scala 20:24]
  reg [31:0] tag_1_62; // @[cache.scala 20:24]
  reg [31:0] tag_1_63; // @[cache.scala 20:24]
  reg [31:0] tag_1_64; // @[cache.scala 20:24]
  reg [31:0] tag_1_65; // @[cache.scala 20:24]
  reg [31:0] tag_1_66; // @[cache.scala 20:24]
  reg [31:0] tag_1_67; // @[cache.scala 20:24]
  reg [31:0] tag_1_68; // @[cache.scala 20:24]
  reg [31:0] tag_1_69; // @[cache.scala 20:24]
  reg [31:0] tag_1_70; // @[cache.scala 20:24]
  reg [31:0] tag_1_71; // @[cache.scala 20:24]
  reg [31:0] tag_1_72; // @[cache.scala 20:24]
  reg [31:0] tag_1_73; // @[cache.scala 20:24]
  reg [31:0] tag_1_74; // @[cache.scala 20:24]
  reg [31:0] tag_1_75; // @[cache.scala 20:24]
  reg [31:0] tag_1_76; // @[cache.scala 20:24]
  reg [31:0] tag_1_77; // @[cache.scala 20:24]
  reg [31:0] tag_1_78; // @[cache.scala 20:24]
  reg [31:0] tag_1_79; // @[cache.scala 20:24]
  reg [31:0] tag_1_80; // @[cache.scala 20:24]
  reg [31:0] tag_1_81; // @[cache.scala 20:24]
  reg [31:0] tag_1_82; // @[cache.scala 20:24]
  reg [31:0] tag_1_83; // @[cache.scala 20:24]
  reg [31:0] tag_1_84; // @[cache.scala 20:24]
  reg [31:0] tag_1_85; // @[cache.scala 20:24]
  reg [31:0] tag_1_86; // @[cache.scala 20:24]
  reg [31:0] tag_1_87; // @[cache.scala 20:24]
  reg [31:0] tag_1_88; // @[cache.scala 20:24]
  reg [31:0] tag_1_89; // @[cache.scala 20:24]
  reg [31:0] tag_1_90; // @[cache.scala 20:24]
  reg [31:0] tag_1_91; // @[cache.scala 20:24]
  reg [31:0] tag_1_92; // @[cache.scala 20:24]
  reg [31:0] tag_1_93; // @[cache.scala 20:24]
  reg [31:0] tag_1_94; // @[cache.scala 20:24]
  reg [31:0] tag_1_95; // @[cache.scala 20:24]
  reg [31:0] tag_1_96; // @[cache.scala 20:24]
  reg [31:0] tag_1_97; // @[cache.scala 20:24]
  reg [31:0] tag_1_98; // @[cache.scala 20:24]
  reg [31:0] tag_1_99; // @[cache.scala 20:24]
  reg [31:0] tag_1_100; // @[cache.scala 20:24]
  reg [31:0] tag_1_101; // @[cache.scala 20:24]
  reg [31:0] tag_1_102; // @[cache.scala 20:24]
  reg [31:0] tag_1_103; // @[cache.scala 20:24]
  reg [31:0] tag_1_104; // @[cache.scala 20:24]
  reg [31:0] tag_1_105; // @[cache.scala 20:24]
  reg [31:0] tag_1_106; // @[cache.scala 20:24]
  reg [31:0] tag_1_107; // @[cache.scala 20:24]
  reg [31:0] tag_1_108; // @[cache.scala 20:24]
  reg [31:0] tag_1_109; // @[cache.scala 20:24]
  reg [31:0] tag_1_110; // @[cache.scala 20:24]
  reg [31:0] tag_1_111; // @[cache.scala 20:24]
  reg [31:0] tag_1_112; // @[cache.scala 20:24]
  reg [31:0] tag_1_113; // @[cache.scala 20:24]
  reg [31:0] tag_1_114; // @[cache.scala 20:24]
  reg [31:0] tag_1_115; // @[cache.scala 20:24]
  reg [31:0] tag_1_116; // @[cache.scala 20:24]
  reg [31:0] tag_1_117; // @[cache.scala 20:24]
  reg [31:0] tag_1_118; // @[cache.scala 20:24]
  reg [31:0] tag_1_119; // @[cache.scala 20:24]
  reg [31:0] tag_1_120; // @[cache.scala 20:24]
  reg [31:0] tag_1_121; // @[cache.scala 20:24]
  reg [31:0] tag_1_122; // @[cache.scala 20:24]
  reg [31:0] tag_1_123; // @[cache.scala 20:24]
  reg [31:0] tag_1_124; // @[cache.scala 20:24]
  reg [31:0] tag_1_125; // @[cache.scala 20:24]
  reg [31:0] tag_1_126; // @[cache.scala 20:24]
  reg [31:0] tag_1_127; // @[cache.scala 20:24]
  reg  valid_0_0; // @[cache.scala 21:26]
  reg  valid_0_1; // @[cache.scala 21:26]
  reg  valid_0_2; // @[cache.scala 21:26]
  reg  valid_0_3; // @[cache.scala 21:26]
  reg  valid_0_4; // @[cache.scala 21:26]
  reg  valid_0_5; // @[cache.scala 21:26]
  reg  valid_0_6; // @[cache.scala 21:26]
  reg  valid_0_7; // @[cache.scala 21:26]
  reg  valid_0_8; // @[cache.scala 21:26]
  reg  valid_0_9; // @[cache.scala 21:26]
  reg  valid_0_10; // @[cache.scala 21:26]
  reg  valid_0_11; // @[cache.scala 21:26]
  reg  valid_0_12; // @[cache.scala 21:26]
  reg  valid_0_13; // @[cache.scala 21:26]
  reg  valid_0_14; // @[cache.scala 21:26]
  reg  valid_0_15; // @[cache.scala 21:26]
  reg  valid_0_16; // @[cache.scala 21:26]
  reg  valid_0_17; // @[cache.scala 21:26]
  reg  valid_0_18; // @[cache.scala 21:26]
  reg  valid_0_19; // @[cache.scala 21:26]
  reg  valid_0_20; // @[cache.scala 21:26]
  reg  valid_0_21; // @[cache.scala 21:26]
  reg  valid_0_22; // @[cache.scala 21:26]
  reg  valid_0_23; // @[cache.scala 21:26]
  reg  valid_0_24; // @[cache.scala 21:26]
  reg  valid_0_25; // @[cache.scala 21:26]
  reg  valid_0_26; // @[cache.scala 21:26]
  reg  valid_0_27; // @[cache.scala 21:26]
  reg  valid_0_28; // @[cache.scala 21:26]
  reg  valid_0_29; // @[cache.scala 21:26]
  reg  valid_0_30; // @[cache.scala 21:26]
  reg  valid_0_31; // @[cache.scala 21:26]
  reg  valid_0_32; // @[cache.scala 21:26]
  reg  valid_0_33; // @[cache.scala 21:26]
  reg  valid_0_34; // @[cache.scala 21:26]
  reg  valid_0_35; // @[cache.scala 21:26]
  reg  valid_0_36; // @[cache.scala 21:26]
  reg  valid_0_37; // @[cache.scala 21:26]
  reg  valid_0_38; // @[cache.scala 21:26]
  reg  valid_0_39; // @[cache.scala 21:26]
  reg  valid_0_40; // @[cache.scala 21:26]
  reg  valid_0_41; // @[cache.scala 21:26]
  reg  valid_0_42; // @[cache.scala 21:26]
  reg  valid_0_43; // @[cache.scala 21:26]
  reg  valid_0_44; // @[cache.scala 21:26]
  reg  valid_0_45; // @[cache.scala 21:26]
  reg  valid_0_46; // @[cache.scala 21:26]
  reg  valid_0_47; // @[cache.scala 21:26]
  reg  valid_0_48; // @[cache.scala 21:26]
  reg  valid_0_49; // @[cache.scala 21:26]
  reg  valid_0_50; // @[cache.scala 21:26]
  reg  valid_0_51; // @[cache.scala 21:26]
  reg  valid_0_52; // @[cache.scala 21:26]
  reg  valid_0_53; // @[cache.scala 21:26]
  reg  valid_0_54; // @[cache.scala 21:26]
  reg  valid_0_55; // @[cache.scala 21:26]
  reg  valid_0_56; // @[cache.scala 21:26]
  reg  valid_0_57; // @[cache.scala 21:26]
  reg  valid_0_58; // @[cache.scala 21:26]
  reg  valid_0_59; // @[cache.scala 21:26]
  reg  valid_0_60; // @[cache.scala 21:26]
  reg  valid_0_61; // @[cache.scala 21:26]
  reg  valid_0_62; // @[cache.scala 21:26]
  reg  valid_0_63; // @[cache.scala 21:26]
  reg  valid_0_64; // @[cache.scala 21:26]
  reg  valid_0_65; // @[cache.scala 21:26]
  reg  valid_0_66; // @[cache.scala 21:26]
  reg  valid_0_67; // @[cache.scala 21:26]
  reg  valid_0_68; // @[cache.scala 21:26]
  reg  valid_0_69; // @[cache.scala 21:26]
  reg  valid_0_70; // @[cache.scala 21:26]
  reg  valid_0_71; // @[cache.scala 21:26]
  reg  valid_0_72; // @[cache.scala 21:26]
  reg  valid_0_73; // @[cache.scala 21:26]
  reg  valid_0_74; // @[cache.scala 21:26]
  reg  valid_0_75; // @[cache.scala 21:26]
  reg  valid_0_76; // @[cache.scala 21:26]
  reg  valid_0_77; // @[cache.scala 21:26]
  reg  valid_0_78; // @[cache.scala 21:26]
  reg  valid_0_79; // @[cache.scala 21:26]
  reg  valid_0_80; // @[cache.scala 21:26]
  reg  valid_0_81; // @[cache.scala 21:26]
  reg  valid_0_82; // @[cache.scala 21:26]
  reg  valid_0_83; // @[cache.scala 21:26]
  reg  valid_0_84; // @[cache.scala 21:26]
  reg  valid_0_85; // @[cache.scala 21:26]
  reg  valid_0_86; // @[cache.scala 21:26]
  reg  valid_0_87; // @[cache.scala 21:26]
  reg  valid_0_88; // @[cache.scala 21:26]
  reg  valid_0_89; // @[cache.scala 21:26]
  reg  valid_0_90; // @[cache.scala 21:26]
  reg  valid_0_91; // @[cache.scala 21:26]
  reg  valid_0_92; // @[cache.scala 21:26]
  reg  valid_0_93; // @[cache.scala 21:26]
  reg  valid_0_94; // @[cache.scala 21:26]
  reg  valid_0_95; // @[cache.scala 21:26]
  reg  valid_0_96; // @[cache.scala 21:26]
  reg  valid_0_97; // @[cache.scala 21:26]
  reg  valid_0_98; // @[cache.scala 21:26]
  reg  valid_0_99; // @[cache.scala 21:26]
  reg  valid_0_100; // @[cache.scala 21:26]
  reg  valid_0_101; // @[cache.scala 21:26]
  reg  valid_0_102; // @[cache.scala 21:26]
  reg  valid_0_103; // @[cache.scala 21:26]
  reg  valid_0_104; // @[cache.scala 21:26]
  reg  valid_0_105; // @[cache.scala 21:26]
  reg  valid_0_106; // @[cache.scala 21:26]
  reg  valid_0_107; // @[cache.scala 21:26]
  reg  valid_0_108; // @[cache.scala 21:26]
  reg  valid_0_109; // @[cache.scala 21:26]
  reg  valid_0_110; // @[cache.scala 21:26]
  reg  valid_0_111; // @[cache.scala 21:26]
  reg  valid_0_112; // @[cache.scala 21:26]
  reg  valid_0_113; // @[cache.scala 21:26]
  reg  valid_0_114; // @[cache.scala 21:26]
  reg  valid_0_115; // @[cache.scala 21:26]
  reg  valid_0_116; // @[cache.scala 21:26]
  reg  valid_0_117; // @[cache.scala 21:26]
  reg  valid_0_118; // @[cache.scala 21:26]
  reg  valid_0_119; // @[cache.scala 21:26]
  reg  valid_0_120; // @[cache.scala 21:26]
  reg  valid_0_121; // @[cache.scala 21:26]
  reg  valid_0_122; // @[cache.scala 21:26]
  reg  valid_0_123; // @[cache.scala 21:26]
  reg  valid_0_124; // @[cache.scala 21:26]
  reg  valid_0_125; // @[cache.scala 21:26]
  reg  valid_0_126; // @[cache.scala 21:26]
  reg  valid_0_127; // @[cache.scala 21:26]
  reg  valid_1_0; // @[cache.scala 22:26]
  reg  valid_1_1; // @[cache.scala 22:26]
  reg  valid_1_2; // @[cache.scala 22:26]
  reg  valid_1_3; // @[cache.scala 22:26]
  reg  valid_1_4; // @[cache.scala 22:26]
  reg  valid_1_5; // @[cache.scala 22:26]
  reg  valid_1_6; // @[cache.scala 22:26]
  reg  valid_1_7; // @[cache.scala 22:26]
  reg  valid_1_8; // @[cache.scala 22:26]
  reg  valid_1_9; // @[cache.scala 22:26]
  reg  valid_1_10; // @[cache.scala 22:26]
  reg  valid_1_11; // @[cache.scala 22:26]
  reg  valid_1_12; // @[cache.scala 22:26]
  reg  valid_1_13; // @[cache.scala 22:26]
  reg  valid_1_14; // @[cache.scala 22:26]
  reg  valid_1_15; // @[cache.scala 22:26]
  reg  valid_1_16; // @[cache.scala 22:26]
  reg  valid_1_17; // @[cache.scala 22:26]
  reg  valid_1_18; // @[cache.scala 22:26]
  reg  valid_1_19; // @[cache.scala 22:26]
  reg  valid_1_20; // @[cache.scala 22:26]
  reg  valid_1_21; // @[cache.scala 22:26]
  reg  valid_1_22; // @[cache.scala 22:26]
  reg  valid_1_23; // @[cache.scala 22:26]
  reg  valid_1_24; // @[cache.scala 22:26]
  reg  valid_1_25; // @[cache.scala 22:26]
  reg  valid_1_26; // @[cache.scala 22:26]
  reg  valid_1_27; // @[cache.scala 22:26]
  reg  valid_1_28; // @[cache.scala 22:26]
  reg  valid_1_29; // @[cache.scala 22:26]
  reg  valid_1_30; // @[cache.scala 22:26]
  reg  valid_1_31; // @[cache.scala 22:26]
  reg  valid_1_32; // @[cache.scala 22:26]
  reg  valid_1_33; // @[cache.scala 22:26]
  reg  valid_1_34; // @[cache.scala 22:26]
  reg  valid_1_35; // @[cache.scala 22:26]
  reg  valid_1_36; // @[cache.scala 22:26]
  reg  valid_1_37; // @[cache.scala 22:26]
  reg  valid_1_38; // @[cache.scala 22:26]
  reg  valid_1_39; // @[cache.scala 22:26]
  reg  valid_1_40; // @[cache.scala 22:26]
  reg  valid_1_41; // @[cache.scala 22:26]
  reg  valid_1_42; // @[cache.scala 22:26]
  reg  valid_1_43; // @[cache.scala 22:26]
  reg  valid_1_44; // @[cache.scala 22:26]
  reg  valid_1_45; // @[cache.scala 22:26]
  reg  valid_1_46; // @[cache.scala 22:26]
  reg  valid_1_47; // @[cache.scala 22:26]
  reg  valid_1_48; // @[cache.scala 22:26]
  reg  valid_1_49; // @[cache.scala 22:26]
  reg  valid_1_50; // @[cache.scala 22:26]
  reg  valid_1_51; // @[cache.scala 22:26]
  reg  valid_1_52; // @[cache.scala 22:26]
  reg  valid_1_53; // @[cache.scala 22:26]
  reg  valid_1_54; // @[cache.scala 22:26]
  reg  valid_1_55; // @[cache.scala 22:26]
  reg  valid_1_56; // @[cache.scala 22:26]
  reg  valid_1_57; // @[cache.scala 22:26]
  reg  valid_1_58; // @[cache.scala 22:26]
  reg  valid_1_59; // @[cache.scala 22:26]
  reg  valid_1_60; // @[cache.scala 22:26]
  reg  valid_1_61; // @[cache.scala 22:26]
  reg  valid_1_62; // @[cache.scala 22:26]
  reg  valid_1_63; // @[cache.scala 22:26]
  reg  valid_1_64; // @[cache.scala 22:26]
  reg  valid_1_65; // @[cache.scala 22:26]
  reg  valid_1_66; // @[cache.scala 22:26]
  reg  valid_1_67; // @[cache.scala 22:26]
  reg  valid_1_68; // @[cache.scala 22:26]
  reg  valid_1_69; // @[cache.scala 22:26]
  reg  valid_1_70; // @[cache.scala 22:26]
  reg  valid_1_71; // @[cache.scala 22:26]
  reg  valid_1_72; // @[cache.scala 22:26]
  reg  valid_1_73; // @[cache.scala 22:26]
  reg  valid_1_74; // @[cache.scala 22:26]
  reg  valid_1_75; // @[cache.scala 22:26]
  reg  valid_1_76; // @[cache.scala 22:26]
  reg  valid_1_77; // @[cache.scala 22:26]
  reg  valid_1_78; // @[cache.scala 22:26]
  reg  valid_1_79; // @[cache.scala 22:26]
  reg  valid_1_80; // @[cache.scala 22:26]
  reg  valid_1_81; // @[cache.scala 22:26]
  reg  valid_1_82; // @[cache.scala 22:26]
  reg  valid_1_83; // @[cache.scala 22:26]
  reg  valid_1_84; // @[cache.scala 22:26]
  reg  valid_1_85; // @[cache.scala 22:26]
  reg  valid_1_86; // @[cache.scala 22:26]
  reg  valid_1_87; // @[cache.scala 22:26]
  reg  valid_1_88; // @[cache.scala 22:26]
  reg  valid_1_89; // @[cache.scala 22:26]
  reg  valid_1_90; // @[cache.scala 22:26]
  reg  valid_1_91; // @[cache.scala 22:26]
  reg  valid_1_92; // @[cache.scala 22:26]
  reg  valid_1_93; // @[cache.scala 22:26]
  reg  valid_1_94; // @[cache.scala 22:26]
  reg  valid_1_95; // @[cache.scala 22:26]
  reg  valid_1_96; // @[cache.scala 22:26]
  reg  valid_1_97; // @[cache.scala 22:26]
  reg  valid_1_98; // @[cache.scala 22:26]
  reg  valid_1_99; // @[cache.scala 22:26]
  reg  valid_1_100; // @[cache.scala 22:26]
  reg  valid_1_101; // @[cache.scala 22:26]
  reg  valid_1_102; // @[cache.scala 22:26]
  reg  valid_1_103; // @[cache.scala 22:26]
  reg  valid_1_104; // @[cache.scala 22:26]
  reg  valid_1_105; // @[cache.scala 22:26]
  reg  valid_1_106; // @[cache.scala 22:26]
  reg  valid_1_107; // @[cache.scala 22:26]
  reg  valid_1_108; // @[cache.scala 22:26]
  reg  valid_1_109; // @[cache.scala 22:26]
  reg  valid_1_110; // @[cache.scala 22:26]
  reg  valid_1_111; // @[cache.scala 22:26]
  reg  valid_1_112; // @[cache.scala 22:26]
  reg  valid_1_113; // @[cache.scala 22:26]
  reg  valid_1_114; // @[cache.scala 22:26]
  reg  valid_1_115; // @[cache.scala 22:26]
  reg  valid_1_116; // @[cache.scala 22:26]
  reg  valid_1_117; // @[cache.scala 22:26]
  reg  valid_1_118; // @[cache.scala 22:26]
  reg  valid_1_119; // @[cache.scala 22:26]
  reg  valid_1_120; // @[cache.scala 22:26]
  reg  valid_1_121; // @[cache.scala 22:26]
  reg  valid_1_122; // @[cache.scala 22:26]
  reg  valid_1_123; // @[cache.scala 22:26]
  reg  valid_1_124; // @[cache.scala 22:26]
  reg  valid_1_125; // @[cache.scala 22:26]
  reg  valid_1_126; // @[cache.scala 22:26]
  reg  valid_1_127; // @[cache.scala 22:26]
  reg  way0_hit; // @[cache.scala 23:27]
  reg  way1_hit; // @[cache.scala 24:27]
  reg [1:0] unuse_way; // @[cache.scala 26:28]
  reg [63:0] receive_data; // @[cache.scala 27:31]
  reg  quene; // @[cache.scala 28:24]
  wire [6:0] index = io_from_ifu_araddr[12:6]; // @[cache.scala 31:35]
  wire [18:0] tag = io_from_ifu_araddr[31:13]; // @[cache.scala 32:33]
  wire [31:0] _GEN_1 = 7'h1 == index ? tag_0_1 : tag_0_0; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_2 = 7'h2 == index ? tag_0_2 : _GEN_1; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_3 = 7'h3 == index ? tag_0_3 : _GEN_2; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_4 = 7'h4 == index ? tag_0_4 : _GEN_3; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_5 = 7'h5 == index ? tag_0_5 : _GEN_4; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_6 = 7'h6 == index ? tag_0_6 : _GEN_5; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_7 = 7'h7 == index ? tag_0_7 : _GEN_6; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_8 = 7'h8 == index ? tag_0_8 : _GEN_7; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_9 = 7'h9 == index ? tag_0_9 : _GEN_8; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_10 = 7'ha == index ? tag_0_10 : _GEN_9; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_11 = 7'hb == index ? tag_0_11 : _GEN_10; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_12 = 7'hc == index ? tag_0_12 : _GEN_11; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_13 = 7'hd == index ? tag_0_13 : _GEN_12; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_14 = 7'he == index ? tag_0_14 : _GEN_13; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_15 = 7'hf == index ? tag_0_15 : _GEN_14; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_16 = 7'h10 == index ? tag_0_16 : _GEN_15; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_17 = 7'h11 == index ? tag_0_17 : _GEN_16; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_18 = 7'h12 == index ? tag_0_18 : _GEN_17; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_19 = 7'h13 == index ? tag_0_19 : _GEN_18; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_20 = 7'h14 == index ? tag_0_20 : _GEN_19; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_21 = 7'h15 == index ? tag_0_21 : _GEN_20; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_22 = 7'h16 == index ? tag_0_22 : _GEN_21; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_23 = 7'h17 == index ? tag_0_23 : _GEN_22; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_24 = 7'h18 == index ? tag_0_24 : _GEN_23; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_25 = 7'h19 == index ? tag_0_25 : _GEN_24; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_26 = 7'h1a == index ? tag_0_26 : _GEN_25; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_27 = 7'h1b == index ? tag_0_27 : _GEN_26; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_28 = 7'h1c == index ? tag_0_28 : _GEN_27; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_29 = 7'h1d == index ? tag_0_29 : _GEN_28; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_30 = 7'h1e == index ? tag_0_30 : _GEN_29; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_31 = 7'h1f == index ? tag_0_31 : _GEN_30; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_32 = 7'h20 == index ? tag_0_32 : _GEN_31; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_33 = 7'h21 == index ? tag_0_33 : _GEN_32; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_34 = 7'h22 == index ? tag_0_34 : _GEN_33; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_35 = 7'h23 == index ? tag_0_35 : _GEN_34; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_36 = 7'h24 == index ? tag_0_36 : _GEN_35; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_37 = 7'h25 == index ? tag_0_37 : _GEN_36; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_38 = 7'h26 == index ? tag_0_38 : _GEN_37; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_39 = 7'h27 == index ? tag_0_39 : _GEN_38; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_40 = 7'h28 == index ? tag_0_40 : _GEN_39; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_41 = 7'h29 == index ? tag_0_41 : _GEN_40; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_42 = 7'h2a == index ? tag_0_42 : _GEN_41; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_43 = 7'h2b == index ? tag_0_43 : _GEN_42; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_44 = 7'h2c == index ? tag_0_44 : _GEN_43; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_45 = 7'h2d == index ? tag_0_45 : _GEN_44; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_46 = 7'h2e == index ? tag_0_46 : _GEN_45; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_47 = 7'h2f == index ? tag_0_47 : _GEN_46; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_48 = 7'h30 == index ? tag_0_48 : _GEN_47; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_49 = 7'h31 == index ? tag_0_49 : _GEN_48; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_50 = 7'h32 == index ? tag_0_50 : _GEN_49; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_51 = 7'h33 == index ? tag_0_51 : _GEN_50; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_52 = 7'h34 == index ? tag_0_52 : _GEN_51; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_53 = 7'h35 == index ? tag_0_53 : _GEN_52; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_54 = 7'h36 == index ? tag_0_54 : _GEN_53; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_55 = 7'h37 == index ? tag_0_55 : _GEN_54; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_56 = 7'h38 == index ? tag_0_56 : _GEN_55; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_57 = 7'h39 == index ? tag_0_57 : _GEN_56; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_58 = 7'h3a == index ? tag_0_58 : _GEN_57; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_59 = 7'h3b == index ? tag_0_59 : _GEN_58; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_60 = 7'h3c == index ? tag_0_60 : _GEN_59; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_61 = 7'h3d == index ? tag_0_61 : _GEN_60; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_62 = 7'h3e == index ? tag_0_62 : _GEN_61; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_63 = 7'h3f == index ? tag_0_63 : _GEN_62; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_64 = 7'h40 == index ? tag_0_64 : _GEN_63; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_65 = 7'h41 == index ? tag_0_65 : _GEN_64; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_66 = 7'h42 == index ? tag_0_66 : _GEN_65; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_67 = 7'h43 == index ? tag_0_67 : _GEN_66; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_68 = 7'h44 == index ? tag_0_68 : _GEN_67; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_69 = 7'h45 == index ? tag_0_69 : _GEN_68; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_70 = 7'h46 == index ? tag_0_70 : _GEN_69; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_71 = 7'h47 == index ? tag_0_71 : _GEN_70; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_72 = 7'h48 == index ? tag_0_72 : _GEN_71; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_73 = 7'h49 == index ? tag_0_73 : _GEN_72; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_74 = 7'h4a == index ? tag_0_74 : _GEN_73; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_75 = 7'h4b == index ? tag_0_75 : _GEN_74; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_76 = 7'h4c == index ? tag_0_76 : _GEN_75; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_77 = 7'h4d == index ? tag_0_77 : _GEN_76; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_78 = 7'h4e == index ? tag_0_78 : _GEN_77; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_79 = 7'h4f == index ? tag_0_79 : _GEN_78; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_80 = 7'h50 == index ? tag_0_80 : _GEN_79; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_81 = 7'h51 == index ? tag_0_81 : _GEN_80; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_82 = 7'h52 == index ? tag_0_82 : _GEN_81; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_83 = 7'h53 == index ? tag_0_83 : _GEN_82; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_84 = 7'h54 == index ? tag_0_84 : _GEN_83; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_85 = 7'h55 == index ? tag_0_85 : _GEN_84; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_86 = 7'h56 == index ? tag_0_86 : _GEN_85; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_87 = 7'h57 == index ? tag_0_87 : _GEN_86; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_88 = 7'h58 == index ? tag_0_88 : _GEN_87; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_89 = 7'h59 == index ? tag_0_89 : _GEN_88; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_90 = 7'h5a == index ? tag_0_90 : _GEN_89; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_91 = 7'h5b == index ? tag_0_91 : _GEN_90; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_92 = 7'h5c == index ? tag_0_92 : _GEN_91; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_93 = 7'h5d == index ? tag_0_93 : _GEN_92; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_94 = 7'h5e == index ? tag_0_94 : _GEN_93; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_95 = 7'h5f == index ? tag_0_95 : _GEN_94; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_96 = 7'h60 == index ? tag_0_96 : _GEN_95; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_97 = 7'h61 == index ? tag_0_97 : _GEN_96; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_98 = 7'h62 == index ? tag_0_98 : _GEN_97; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_99 = 7'h63 == index ? tag_0_99 : _GEN_98; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_100 = 7'h64 == index ? tag_0_100 : _GEN_99; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_101 = 7'h65 == index ? tag_0_101 : _GEN_100; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_102 = 7'h66 == index ? tag_0_102 : _GEN_101; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_103 = 7'h67 == index ? tag_0_103 : _GEN_102; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_104 = 7'h68 == index ? tag_0_104 : _GEN_103; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_105 = 7'h69 == index ? tag_0_105 : _GEN_104; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_106 = 7'h6a == index ? tag_0_106 : _GEN_105; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_107 = 7'h6b == index ? tag_0_107 : _GEN_106; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_108 = 7'h6c == index ? tag_0_108 : _GEN_107; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_109 = 7'h6d == index ? tag_0_109 : _GEN_108; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_110 = 7'h6e == index ? tag_0_110 : _GEN_109; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_111 = 7'h6f == index ? tag_0_111 : _GEN_110; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_112 = 7'h70 == index ? tag_0_112 : _GEN_111; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_113 = 7'h71 == index ? tag_0_113 : _GEN_112; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_114 = 7'h72 == index ? tag_0_114 : _GEN_113; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_115 = 7'h73 == index ? tag_0_115 : _GEN_114; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_116 = 7'h74 == index ? tag_0_116 : _GEN_115; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_117 = 7'h75 == index ? tag_0_117 : _GEN_116; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_118 = 7'h76 == index ? tag_0_118 : _GEN_117; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_119 = 7'h77 == index ? tag_0_119 : _GEN_118; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_120 = 7'h78 == index ? tag_0_120 : _GEN_119; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_121 = 7'h79 == index ? tag_0_121 : _GEN_120; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_122 = 7'h7a == index ? tag_0_122 : _GEN_121; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_123 = 7'h7b == index ? tag_0_123 : _GEN_122; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_124 = 7'h7c == index ? tag_0_124 : _GEN_123; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_125 = 7'h7d == index ? tag_0_125 : _GEN_124; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_126 = 7'h7e == index ? tag_0_126 : _GEN_125; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_127 = 7'h7f == index ? tag_0_127 : _GEN_126; // @[cache.scala 34:{24,24}]
  wire [31:0] _GEN_7705 = {{13'd0}, tag}; // @[cache.scala 34:24]
  wire  _GEN_129 = 7'h1 == index ? valid_0_1 : valid_0_0; // @[cache.scala 34:{50,50}]
  wire  _GEN_130 = 7'h2 == index ? valid_0_2 : _GEN_129; // @[cache.scala 34:{50,50}]
  wire  _GEN_131 = 7'h3 == index ? valid_0_3 : _GEN_130; // @[cache.scala 34:{50,50}]
  wire  _GEN_132 = 7'h4 == index ? valid_0_4 : _GEN_131; // @[cache.scala 34:{50,50}]
  wire  _GEN_133 = 7'h5 == index ? valid_0_5 : _GEN_132; // @[cache.scala 34:{50,50}]
  wire  _GEN_134 = 7'h6 == index ? valid_0_6 : _GEN_133; // @[cache.scala 34:{50,50}]
  wire  _GEN_135 = 7'h7 == index ? valid_0_7 : _GEN_134; // @[cache.scala 34:{50,50}]
  wire  _GEN_136 = 7'h8 == index ? valid_0_8 : _GEN_135; // @[cache.scala 34:{50,50}]
  wire  _GEN_137 = 7'h9 == index ? valid_0_9 : _GEN_136; // @[cache.scala 34:{50,50}]
  wire  _GEN_138 = 7'ha == index ? valid_0_10 : _GEN_137; // @[cache.scala 34:{50,50}]
  wire  _GEN_139 = 7'hb == index ? valid_0_11 : _GEN_138; // @[cache.scala 34:{50,50}]
  wire  _GEN_140 = 7'hc == index ? valid_0_12 : _GEN_139; // @[cache.scala 34:{50,50}]
  wire  _GEN_141 = 7'hd == index ? valid_0_13 : _GEN_140; // @[cache.scala 34:{50,50}]
  wire  _GEN_142 = 7'he == index ? valid_0_14 : _GEN_141; // @[cache.scala 34:{50,50}]
  wire  _GEN_143 = 7'hf == index ? valid_0_15 : _GEN_142; // @[cache.scala 34:{50,50}]
  wire  _GEN_144 = 7'h10 == index ? valid_0_16 : _GEN_143; // @[cache.scala 34:{50,50}]
  wire  _GEN_145 = 7'h11 == index ? valid_0_17 : _GEN_144; // @[cache.scala 34:{50,50}]
  wire  _GEN_146 = 7'h12 == index ? valid_0_18 : _GEN_145; // @[cache.scala 34:{50,50}]
  wire  _GEN_147 = 7'h13 == index ? valid_0_19 : _GEN_146; // @[cache.scala 34:{50,50}]
  wire  _GEN_148 = 7'h14 == index ? valid_0_20 : _GEN_147; // @[cache.scala 34:{50,50}]
  wire  _GEN_149 = 7'h15 == index ? valid_0_21 : _GEN_148; // @[cache.scala 34:{50,50}]
  wire  _GEN_150 = 7'h16 == index ? valid_0_22 : _GEN_149; // @[cache.scala 34:{50,50}]
  wire  _GEN_151 = 7'h17 == index ? valid_0_23 : _GEN_150; // @[cache.scala 34:{50,50}]
  wire  _GEN_152 = 7'h18 == index ? valid_0_24 : _GEN_151; // @[cache.scala 34:{50,50}]
  wire  _GEN_153 = 7'h19 == index ? valid_0_25 : _GEN_152; // @[cache.scala 34:{50,50}]
  wire  _GEN_154 = 7'h1a == index ? valid_0_26 : _GEN_153; // @[cache.scala 34:{50,50}]
  wire  _GEN_155 = 7'h1b == index ? valid_0_27 : _GEN_154; // @[cache.scala 34:{50,50}]
  wire  _GEN_156 = 7'h1c == index ? valid_0_28 : _GEN_155; // @[cache.scala 34:{50,50}]
  wire  _GEN_157 = 7'h1d == index ? valid_0_29 : _GEN_156; // @[cache.scala 34:{50,50}]
  wire  _GEN_158 = 7'h1e == index ? valid_0_30 : _GEN_157; // @[cache.scala 34:{50,50}]
  wire  _GEN_159 = 7'h1f == index ? valid_0_31 : _GEN_158; // @[cache.scala 34:{50,50}]
  wire  _GEN_160 = 7'h20 == index ? valid_0_32 : _GEN_159; // @[cache.scala 34:{50,50}]
  wire  _GEN_161 = 7'h21 == index ? valid_0_33 : _GEN_160; // @[cache.scala 34:{50,50}]
  wire  _GEN_162 = 7'h22 == index ? valid_0_34 : _GEN_161; // @[cache.scala 34:{50,50}]
  wire  _GEN_163 = 7'h23 == index ? valid_0_35 : _GEN_162; // @[cache.scala 34:{50,50}]
  wire  _GEN_164 = 7'h24 == index ? valid_0_36 : _GEN_163; // @[cache.scala 34:{50,50}]
  wire  _GEN_165 = 7'h25 == index ? valid_0_37 : _GEN_164; // @[cache.scala 34:{50,50}]
  wire  _GEN_166 = 7'h26 == index ? valid_0_38 : _GEN_165; // @[cache.scala 34:{50,50}]
  wire  _GEN_167 = 7'h27 == index ? valid_0_39 : _GEN_166; // @[cache.scala 34:{50,50}]
  wire  _GEN_168 = 7'h28 == index ? valid_0_40 : _GEN_167; // @[cache.scala 34:{50,50}]
  wire  _GEN_169 = 7'h29 == index ? valid_0_41 : _GEN_168; // @[cache.scala 34:{50,50}]
  wire  _GEN_170 = 7'h2a == index ? valid_0_42 : _GEN_169; // @[cache.scala 34:{50,50}]
  wire  _GEN_171 = 7'h2b == index ? valid_0_43 : _GEN_170; // @[cache.scala 34:{50,50}]
  wire  _GEN_172 = 7'h2c == index ? valid_0_44 : _GEN_171; // @[cache.scala 34:{50,50}]
  wire  _GEN_173 = 7'h2d == index ? valid_0_45 : _GEN_172; // @[cache.scala 34:{50,50}]
  wire  _GEN_174 = 7'h2e == index ? valid_0_46 : _GEN_173; // @[cache.scala 34:{50,50}]
  wire  _GEN_175 = 7'h2f == index ? valid_0_47 : _GEN_174; // @[cache.scala 34:{50,50}]
  wire  _GEN_176 = 7'h30 == index ? valid_0_48 : _GEN_175; // @[cache.scala 34:{50,50}]
  wire  _GEN_177 = 7'h31 == index ? valid_0_49 : _GEN_176; // @[cache.scala 34:{50,50}]
  wire  _GEN_178 = 7'h32 == index ? valid_0_50 : _GEN_177; // @[cache.scala 34:{50,50}]
  wire  _GEN_179 = 7'h33 == index ? valid_0_51 : _GEN_178; // @[cache.scala 34:{50,50}]
  wire  _GEN_180 = 7'h34 == index ? valid_0_52 : _GEN_179; // @[cache.scala 34:{50,50}]
  wire  _GEN_181 = 7'h35 == index ? valid_0_53 : _GEN_180; // @[cache.scala 34:{50,50}]
  wire  _GEN_182 = 7'h36 == index ? valid_0_54 : _GEN_181; // @[cache.scala 34:{50,50}]
  wire  _GEN_183 = 7'h37 == index ? valid_0_55 : _GEN_182; // @[cache.scala 34:{50,50}]
  wire  _GEN_184 = 7'h38 == index ? valid_0_56 : _GEN_183; // @[cache.scala 34:{50,50}]
  wire  _GEN_185 = 7'h39 == index ? valid_0_57 : _GEN_184; // @[cache.scala 34:{50,50}]
  wire  _GEN_186 = 7'h3a == index ? valid_0_58 : _GEN_185; // @[cache.scala 34:{50,50}]
  wire  _GEN_187 = 7'h3b == index ? valid_0_59 : _GEN_186; // @[cache.scala 34:{50,50}]
  wire  _GEN_188 = 7'h3c == index ? valid_0_60 : _GEN_187; // @[cache.scala 34:{50,50}]
  wire  _GEN_189 = 7'h3d == index ? valid_0_61 : _GEN_188; // @[cache.scala 34:{50,50}]
  wire  _GEN_190 = 7'h3e == index ? valid_0_62 : _GEN_189; // @[cache.scala 34:{50,50}]
  wire  _GEN_191 = 7'h3f == index ? valid_0_63 : _GEN_190; // @[cache.scala 34:{50,50}]
  wire  _GEN_192 = 7'h40 == index ? valid_0_64 : _GEN_191; // @[cache.scala 34:{50,50}]
  wire  _GEN_193 = 7'h41 == index ? valid_0_65 : _GEN_192; // @[cache.scala 34:{50,50}]
  wire  _GEN_194 = 7'h42 == index ? valid_0_66 : _GEN_193; // @[cache.scala 34:{50,50}]
  wire  _GEN_195 = 7'h43 == index ? valid_0_67 : _GEN_194; // @[cache.scala 34:{50,50}]
  wire  _GEN_196 = 7'h44 == index ? valid_0_68 : _GEN_195; // @[cache.scala 34:{50,50}]
  wire  _GEN_197 = 7'h45 == index ? valid_0_69 : _GEN_196; // @[cache.scala 34:{50,50}]
  wire  _GEN_198 = 7'h46 == index ? valid_0_70 : _GEN_197; // @[cache.scala 34:{50,50}]
  wire  _GEN_199 = 7'h47 == index ? valid_0_71 : _GEN_198; // @[cache.scala 34:{50,50}]
  wire  _GEN_200 = 7'h48 == index ? valid_0_72 : _GEN_199; // @[cache.scala 34:{50,50}]
  wire  _GEN_201 = 7'h49 == index ? valid_0_73 : _GEN_200; // @[cache.scala 34:{50,50}]
  wire  _GEN_202 = 7'h4a == index ? valid_0_74 : _GEN_201; // @[cache.scala 34:{50,50}]
  wire  _GEN_203 = 7'h4b == index ? valid_0_75 : _GEN_202; // @[cache.scala 34:{50,50}]
  wire  _GEN_204 = 7'h4c == index ? valid_0_76 : _GEN_203; // @[cache.scala 34:{50,50}]
  wire  _GEN_205 = 7'h4d == index ? valid_0_77 : _GEN_204; // @[cache.scala 34:{50,50}]
  wire  _GEN_206 = 7'h4e == index ? valid_0_78 : _GEN_205; // @[cache.scala 34:{50,50}]
  wire  _GEN_207 = 7'h4f == index ? valid_0_79 : _GEN_206; // @[cache.scala 34:{50,50}]
  wire  _GEN_208 = 7'h50 == index ? valid_0_80 : _GEN_207; // @[cache.scala 34:{50,50}]
  wire  _GEN_209 = 7'h51 == index ? valid_0_81 : _GEN_208; // @[cache.scala 34:{50,50}]
  wire  _GEN_210 = 7'h52 == index ? valid_0_82 : _GEN_209; // @[cache.scala 34:{50,50}]
  wire  _GEN_211 = 7'h53 == index ? valid_0_83 : _GEN_210; // @[cache.scala 34:{50,50}]
  wire  _GEN_212 = 7'h54 == index ? valid_0_84 : _GEN_211; // @[cache.scala 34:{50,50}]
  wire  _GEN_213 = 7'h55 == index ? valid_0_85 : _GEN_212; // @[cache.scala 34:{50,50}]
  wire  _GEN_214 = 7'h56 == index ? valid_0_86 : _GEN_213; // @[cache.scala 34:{50,50}]
  wire  _GEN_215 = 7'h57 == index ? valid_0_87 : _GEN_214; // @[cache.scala 34:{50,50}]
  wire  _GEN_216 = 7'h58 == index ? valid_0_88 : _GEN_215; // @[cache.scala 34:{50,50}]
  wire  _GEN_217 = 7'h59 == index ? valid_0_89 : _GEN_216; // @[cache.scala 34:{50,50}]
  wire  _GEN_218 = 7'h5a == index ? valid_0_90 : _GEN_217; // @[cache.scala 34:{50,50}]
  wire  _GEN_219 = 7'h5b == index ? valid_0_91 : _GEN_218; // @[cache.scala 34:{50,50}]
  wire  _GEN_220 = 7'h5c == index ? valid_0_92 : _GEN_219; // @[cache.scala 34:{50,50}]
  wire  _GEN_221 = 7'h5d == index ? valid_0_93 : _GEN_220; // @[cache.scala 34:{50,50}]
  wire  _GEN_222 = 7'h5e == index ? valid_0_94 : _GEN_221; // @[cache.scala 34:{50,50}]
  wire  _GEN_223 = 7'h5f == index ? valid_0_95 : _GEN_222; // @[cache.scala 34:{50,50}]
  wire  _GEN_224 = 7'h60 == index ? valid_0_96 : _GEN_223; // @[cache.scala 34:{50,50}]
  wire  _GEN_225 = 7'h61 == index ? valid_0_97 : _GEN_224; // @[cache.scala 34:{50,50}]
  wire  _GEN_226 = 7'h62 == index ? valid_0_98 : _GEN_225; // @[cache.scala 34:{50,50}]
  wire  _GEN_227 = 7'h63 == index ? valid_0_99 : _GEN_226; // @[cache.scala 34:{50,50}]
  wire  _GEN_228 = 7'h64 == index ? valid_0_100 : _GEN_227; // @[cache.scala 34:{50,50}]
  wire  _GEN_229 = 7'h65 == index ? valid_0_101 : _GEN_228; // @[cache.scala 34:{50,50}]
  wire  _GEN_230 = 7'h66 == index ? valid_0_102 : _GEN_229; // @[cache.scala 34:{50,50}]
  wire  _GEN_231 = 7'h67 == index ? valid_0_103 : _GEN_230; // @[cache.scala 34:{50,50}]
  wire  _GEN_232 = 7'h68 == index ? valid_0_104 : _GEN_231; // @[cache.scala 34:{50,50}]
  wire  _GEN_233 = 7'h69 == index ? valid_0_105 : _GEN_232; // @[cache.scala 34:{50,50}]
  wire  _GEN_234 = 7'h6a == index ? valid_0_106 : _GEN_233; // @[cache.scala 34:{50,50}]
  wire  _GEN_235 = 7'h6b == index ? valid_0_107 : _GEN_234; // @[cache.scala 34:{50,50}]
  wire  _GEN_236 = 7'h6c == index ? valid_0_108 : _GEN_235; // @[cache.scala 34:{50,50}]
  wire  _GEN_237 = 7'h6d == index ? valid_0_109 : _GEN_236; // @[cache.scala 34:{50,50}]
  wire  _GEN_238 = 7'h6e == index ? valid_0_110 : _GEN_237; // @[cache.scala 34:{50,50}]
  wire  _GEN_239 = 7'h6f == index ? valid_0_111 : _GEN_238; // @[cache.scala 34:{50,50}]
  wire  _GEN_240 = 7'h70 == index ? valid_0_112 : _GEN_239; // @[cache.scala 34:{50,50}]
  wire  _GEN_241 = 7'h71 == index ? valid_0_113 : _GEN_240; // @[cache.scala 34:{50,50}]
  wire  _GEN_242 = 7'h72 == index ? valid_0_114 : _GEN_241; // @[cache.scala 34:{50,50}]
  wire  _GEN_243 = 7'h73 == index ? valid_0_115 : _GEN_242; // @[cache.scala 34:{50,50}]
  wire  _GEN_244 = 7'h74 == index ? valid_0_116 : _GEN_243; // @[cache.scala 34:{50,50}]
  wire  _GEN_245 = 7'h75 == index ? valid_0_117 : _GEN_244; // @[cache.scala 34:{50,50}]
  wire  _GEN_246 = 7'h76 == index ? valid_0_118 : _GEN_245; // @[cache.scala 34:{50,50}]
  wire  _GEN_247 = 7'h77 == index ? valid_0_119 : _GEN_246; // @[cache.scala 34:{50,50}]
  wire  _GEN_248 = 7'h78 == index ? valid_0_120 : _GEN_247; // @[cache.scala 34:{50,50}]
  wire  _GEN_249 = 7'h79 == index ? valid_0_121 : _GEN_248; // @[cache.scala 34:{50,50}]
  wire  _GEN_250 = 7'h7a == index ? valid_0_122 : _GEN_249; // @[cache.scala 34:{50,50}]
  wire  _GEN_251 = 7'h7b == index ? valid_0_123 : _GEN_250; // @[cache.scala 34:{50,50}]
  wire  _GEN_252 = 7'h7c == index ? valid_0_124 : _GEN_251; // @[cache.scala 34:{50,50}]
  wire  _GEN_253 = 7'h7d == index ? valid_0_125 : _GEN_252; // @[cache.scala 34:{50,50}]
  wire  _GEN_254 = 7'h7e == index ? valid_0_126 : _GEN_253; // @[cache.scala 34:{50,50}]
  wire  _GEN_255 = 7'h7f == index ? valid_0_127 : _GEN_254; // @[cache.scala 34:{50,50}]
  wire  _GEN_256 = _GEN_127 == _GEN_7705 & _GEN_255 | way0_hit; // @[cache.scala 34:57 35:19 23:27]
  wire [31:0] _GEN_258 = 7'h1 == index ? tag_1_1 : tag_1_0; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_259 = 7'h2 == index ? tag_1_2 : _GEN_258; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_260 = 7'h3 == index ? tag_1_3 : _GEN_259; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_261 = 7'h4 == index ? tag_1_4 : _GEN_260; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_262 = 7'h5 == index ? tag_1_5 : _GEN_261; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_263 = 7'h6 == index ? tag_1_6 : _GEN_262; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_264 = 7'h7 == index ? tag_1_7 : _GEN_263; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_265 = 7'h8 == index ? tag_1_8 : _GEN_264; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_266 = 7'h9 == index ? tag_1_9 : _GEN_265; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_267 = 7'ha == index ? tag_1_10 : _GEN_266; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_268 = 7'hb == index ? tag_1_11 : _GEN_267; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_269 = 7'hc == index ? tag_1_12 : _GEN_268; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_270 = 7'hd == index ? tag_1_13 : _GEN_269; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_271 = 7'he == index ? tag_1_14 : _GEN_270; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_272 = 7'hf == index ? tag_1_15 : _GEN_271; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_273 = 7'h10 == index ? tag_1_16 : _GEN_272; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_274 = 7'h11 == index ? tag_1_17 : _GEN_273; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_275 = 7'h12 == index ? tag_1_18 : _GEN_274; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_276 = 7'h13 == index ? tag_1_19 : _GEN_275; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_277 = 7'h14 == index ? tag_1_20 : _GEN_276; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_278 = 7'h15 == index ? tag_1_21 : _GEN_277; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_279 = 7'h16 == index ? tag_1_22 : _GEN_278; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_280 = 7'h17 == index ? tag_1_23 : _GEN_279; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_281 = 7'h18 == index ? tag_1_24 : _GEN_280; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_282 = 7'h19 == index ? tag_1_25 : _GEN_281; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_283 = 7'h1a == index ? tag_1_26 : _GEN_282; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_284 = 7'h1b == index ? tag_1_27 : _GEN_283; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_285 = 7'h1c == index ? tag_1_28 : _GEN_284; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_286 = 7'h1d == index ? tag_1_29 : _GEN_285; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_287 = 7'h1e == index ? tag_1_30 : _GEN_286; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_288 = 7'h1f == index ? tag_1_31 : _GEN_287; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_289 = 7'h20 == index ? tag_1_32 : _GEN_288; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_290 = 7'h21 == index ? tag_1_33 : _GEN_289; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_291 = 7'h22 == index ? tag_1_34 : _GEN_290; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_292 = 7'h23 == index ? tag_1_35 : _GEN_291; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_293 = 7'h24 == index ? tag_1_36 : _GEN_292; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_294 = 7'h25 == index ? tag_1_37 : _GEN_293; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_295 = 7'h26 == index ? tag_1_38 : _GEN_294; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_296 = 7'h27 == index ? tag_1_39 : _GEN_295; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_297 = 7'h28 == index ? tag_1_40 : _GEN_296; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_298 = 7'h29 == index ? tag_1_41 : _GEN_297; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_299 = 7'h2a == index ? tag_1_42 : _GEN_298; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_300 = 7'h2b == index ? tag_1_43 : _GEN_299; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_301 = 7'h2c == index ? tag_1_44 : _GEN_300; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_302 = 7'h2d == index ? tag_1_45 : _GEN_301; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_303 = 7'h2e == index ? tag_1_46 : _GEN_302; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_304 = 7'h2f == index ? tag_1_47 : _GEN_303; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_305 = 7'h30 == index ? tag_1_48 : _GEN_304; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_306 = 7'h31 == index ? tag_1_49 : _GEN_305; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_307 = 7'h32 == index ? tag_1_50 : _GEN_306; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_308 = 7'h33 == index ? tag_1_51 : _GEN_307; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_309 = 7'h34 == index ? tag_1_52 : _GEN_308; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_310 = 7'h35 == index ? tag_1_53 : _GEN_309; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_311 = 7'h36 == index ? tag_1_54 : _GEN_310; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_312 = 7'h37 == index ? tag_1_55 : _GEN_311; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_313 = 7'h38 == index ? tag_1_56 : _GEN_312; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_314 = 7'h39 == index ? tag_1_57 : _GEN_313; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_315 = 7'h3a == index ? tag_1_58 : _GEN_314; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_316 = 7'h3b == index ? tag_1_59 : _GEN_315; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_317 = 7'h3c == index ? tag_1_60 : _GEN_316; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_318 = 7'h3d == index ? tag_1_61 : _GEN_317; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_319 = 7'h3e == index ? tag_1_62 : _GEN_318; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_320 = 7'h3f == index ? tag_1_63 : _GEN_319; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_321 = 7'h40 == index ? tag_1_64 : _GEN_320; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_322 = 7'h41 == index ? tag_1_65 : _GEN_321; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_323 = 7'h42 == index ? tag_1_66 : _GEN_322; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_324 = 7'h43 == index ? tag_1_67 : _GEN_323; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_325 = 7'h44 == index ? tag_1_68 : _GEN_324; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_326 = 7'h45 == index ? tag_1_69 : _GEN_325; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_327 = 7'h46 == index ? tag_1_70 : _GEN_326; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_328 = 7'h47 == index ? tag_1_71 : _GEN_327; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_329 = 7'h48 == index ? tag_1_72 : _GEN_328; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_330 = 7'h49 == index ? tag_1_73 : _GEN_329; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_331 = 7'h4a == index ? tag_1_74 : _GEN_330; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_332 = 7'h4b == index ? tag_1_75 : _GEN_331; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_333 = 7'h4c == index ? tag_1_76 : _GEN_332; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_334 = 7'h4d == index ? tag_1_77 : _GEN_333; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_335 = 7'h4e == index ? tag_1_78 : _GEN_334; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_336 = 7'h4f == index ? tag_1_79 : _GEN_335; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_337 = 7'h50 == index ? tag_1_80 : _GEN_336; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_338 = 7'h51 == index ? tag_1_81 : _GEN_337; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_339 = 7'h52 == index ? tag_1_82 : _GEN_338; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_340 = 7'h53 == index ? tag_1_83 : _GEN_339; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_341 = 7'h54 == index ? tag_1_84 : _GEN_340; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_342 = 7'h55 == index ? tag_1_85 : _GEN_341; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_343 = 7'h56 == index ? tag_1_86 : _GEN_342; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_344 = 7'h57 == index ? tag_1_87 : _GEN_343; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_345 = 7'h58 == index ? tag_1_88 : _GEN_344; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_346 = 7'h59 == index ? tag_1_89 : _GEN_345; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_347 = 7'h5a == index ? tag_1_90 : _GEN_346; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_348 = 7'h5b == index ? tag_1_91 : _GEN_347; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_349 = 7'h5c == index ? tag_1_92 : _GEN_348; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_350 = 7'h5d == index ? tag_1_93 : _GEN_349; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_351 = 7'h5e == index ? tag_1_94 : _GEN_350; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_352 = 7'h5f == index ? tag_1_95 : _GEN_351; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_353 = 7'h60 == index ? tag_1_96 : _GEN_352; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_354 = 7'h61 == index ? tag_1_97 : _GEN_353; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_355 = 7'h62 == index ? tag_1_98 : _GEN_354; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_356 = 7'h63 == index ? tag_1_99 : _GEN_355; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_357 = 7'h64 == index ? tag_1_100 : _GEN_356; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_358 = 7'h65 == index ? tag_1_101 : _GEN_357; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_359 = 7'h66 == index ? tag_1_102 : _GEN_358; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_360 = 7'h67 == index ? tag_1_103 : _GEN_359; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_361 = 7'h68 == index ? tag_1_104 : _GEN_360; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_362 = 7'h69 == index ? tag_1_105 : _GEN_361; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_363 = 7'h6a == index ? tag_1_106 : _GEN_362; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_364 = 7'h6b == index ? tag_1_107 : _GEN_363; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_365 = 7'h6c == index ? tag_1_108 : _GEN_364; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_366 = 7'h6d == index ? tag_1_109 : _GEN_365; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_367 = 7'h6e == index ? tag_1_110 : _GEN_366; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_368 = 7'h6f == index ? tag_1_111 : _GEN_367; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_369 = 7'h70 == index ? tag_1_112 : _GEN_368; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_370 = 7'h71 == index ? tag_1_113 : _GEN_369; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_371 = 7'h72 == index ? tag_1_114 : _GEN_370; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_372 = 7'h73 == index ? tag_1_115 : _GEN_371; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_373 = 7'h74 == index ? tag_1_116 : _GEN_372; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_374 = 7'h75 == index ? tag_1_117 : _GEN_373; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_375 = 7'h76 == index ? tag_1_118 : _GEN_374; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_376 = 7'h77 == index ? tag_1_119 : _GEN_375; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_377 = 7'h78 == index ? tag_1_120 : _GEN_376; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_378 = 7'h79 == index ? tag_1_121 : _GEN_377; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_379 = 7'h7a == index ? tag_1_122 : _GEN_378; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_380 = 7'h7b == index ? tag_1_123 : _GEN_379; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_381 = 7'h7c == index ? tag_1_124 : _GEN_380; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_382 = 7'h7d == index ? tag_1_125 : _GEN_381; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_383 = 7'h7e == index ? tag_1_126 : _GEN_382; // @[cache.scala 37:{24,24}]
  wire [31:0] _GEN_384 = 7'h7f == index ? tag_1_127 : _GEN_383; // @[cache.scala 37:{24,24}]
  wire  _GEN_386 = 7'h1 == index ? valid_1_1 : valid_1_0; // @[cache.scala 37:{50,50}]
  wire  _GEN_387 = 7'h2 == index ? valid_1_2 : _GEN_386; // @[cache.scala 37:{50,50}]
  wire  _GEN_388 = 7'h3 == index ? valid_1_3 : _GEN_387; // @[cache.scala 37:{50,50}]
  wire  _GEN_389 = 7'h4 == index ? valid_1_4 : _GEN_388; // @[cache.scala 37:{50,50}]
  wire  _GEN_390 = 7'h5 == index ? valid_1_5 : _GEN_389; // @[cache.scala 37:{50,50}]
  wire  _GEN_391 = 7'h6 == index ? valid_1_6 : _GEN_390; // @[cache.scala 37:{50,50}]
  wire  _GEN_392 = 7'h7 == index ? valid_1_7 : _GEN_391; // @[cache.scala 37:{50,50}]
  wire  _GEN_393 = 7'h8 == index ? valid_1_8 : _GEN_392; // @[cache.scala 37:{50,50}]
  wire  _GEN_394 = 7'h9 == index ? valid_1_9 : _GEN_393; // @[cache.scala 37:{50,50}]
  wire  _GEN_395 = 7'ha == index ? valid_1_10 : _GEN_394; // @[cache.scala 37:{50,50}]
  wire  _GEN_396 = 7'hb == index ? valid_1_11 : _GEN_395; // @[cache.scala 37:{50,50}]
  wire  _GEN_397 = 7'hc == index ? valid_1_12 : _GEN_396; // @[cache.scala 37:{50,50}]
  wire  _GEN_398 = 7'hd == index ? valid_1_13 : _GEN_397; // @[cache.scala 37:{50,50}]
  wire  _GEN_399 = 7'he == index ? valid_1_14 : _GEN_398; // @[cache.scala 37:{50,50}]
  wire  _GEN_400 = 7'hf == index ? valid_1_15 : _GEN_399; // @[cache.scala 37:{50,50}]
  wire  _GEN_401 = 7'h10 == index ? valid_1_16 : _GEN_400; // @[cache.scala 37:{50,50}]
  wire  _GEN_402 = 7'h11 == index ? valid_1_17 : _GEN_401; // @[cache.scala 37:{50,50}]
  wire  _GEN_403 = 7'h12 == index ? valid_1_18 : _GEN_402; // @[cache.scala 37:{50,50}]
  wire  _GEN_404 = 7'h13 == index ? valid_1_19 : _GEN_403; // @[cache.scala 37:{50,50}]
  wire  _GEN_405 = 7'h14 == index ? valid_1_20 : _GEN_404; // @[cache.scala 37:{50,50}]
  wire  _GEN_406 = 7'h15 == index ? valid_1_21 : _GEN_405; // @[cache.scala 37:{50,50}]
  wire  _GEN_407 = 7'h16 == index ? valid_1_22 : _GEN_406; // @[cache.scala 37:{50,50}]
  wire  _GEN_408 = 7'h17 == index ? valid_1_23 : _GEN_407; // @[cache.scala 37:{50,50}]
  wire  _GEN_409 = 7'h18 == index ? valid_1_24 : _GEN_408; // @[cache.scala 37:{50,50}]
  wire  _GEN_410 = 7'h19 == index ? valid_1_25 : _GEN_409; // @[cache.scala 37:{50,50}]
  wire  _GEN_411 = 7'h1a == index ? valid_1_26 : _GEN_410; // @[cache.scala 37:{50,50}]
  wire  _GEN_412 = 7'h1b == index ? valid_1_27 : _GEN_411; // @[cache.scala 37:{50,50}]
  wire  _GEN_413 = 7'h1c == index ? valid_1_28 : _GEN_412; // @[cache.scala 37:{50,50}]
  wire  _GEN_414 = 7'h1d == index ? valid_1_29 : _GEN_413; // @[cache.scala 37:{50,50}]
  wire  _GEN_415 = 7'h1e == index ? valid_1_30 : _GEN_414; // @[cache.scala 37:{50,50}]
  wire  _GEN_416 = 7'h1f == index ? valid_1_31 : _GEN_415; // @[cache.scala 37:{50,50}]
  wire  _GEN_417 = 7'h20 == index ? valid_1_32 : _GEN_416; // @[cache.scala 37:{50,50}]
  wire  _GEN_418 = 7'h21 == index ? valid_1_33 : _GEN_417; // @[cache.scala 37:{50,50}]
  wire  _GEN_419 = 7'h22 == index ? valid_1_34 : _GEN_418; // @[cache.scala 37:{50,50}]
  wire  _GEN_420 = 7'h23 == index ? valid_1_35 : _GEN_419; // @[cache.scala 37:{50,50}]
  wire  _GEN_421 = 7'h24 == index ? valid_1_36 : _GEN_420; // @[cache.scala 37:{50,50}]
  wire  _GEN_422 = 7'h25 == index ? valid_1_37 : _GEN_421; // @[cache.scala 37:{50,50}]
  wire  _GEN_423 = 7'h26 == index ? valid_1_38 : _GEN_422; // @[cache.scala 37:{50,50}]
  wire  _GEN_424 = 7'h27 == index ? valid_1_39 : _GEN_423; // @[cache.scala 37:{50,50}]
  wire  _GEN_425 = 7'h28 == index ? valid_1_40 : _GEN_424; // @[cache.scala 37:{50,50}]
  wire  _GEN_426 = 7'h29 == index ? valid_1_41 : _GEN_425; // @[cache.scala 37:{50,50}]
  wire  _GEN_427 = 7'h2a == index ? valid_1_42 : _GEN_426; // @[cache.scala 37:{50,50}]
  wire  _GEN_428 = 7'h2b == index ? valid_1_43 : _GEN_427; // @[cache.scala 37:{50,50}]
  wire  _GEN_429 = 7'h2c == index ? valid_1_44 : _GEN_428; // @[cache.scala 37:{50,50}]
  wire  _GEN_430 = 7'h2d == index ? valid_1_45 : _GEN_429; // @[cache.scala 37:{50,50}]
  wire  _GEN_431 = 7'h2e == index ? valid_1_46 : _GEN_430; // @[cache.scala 37:{50,50}]
  wire  _GEN_432 = 7'h2f == index ? valid_1_47 : _GEN_431; // @[cache.scala 37:{50,50}]
  wire  _GEN_433 = 7'h30 == index ? valid_1_48 : _GEN_432; // @[cache.scala 37:{50,50}]
  wire  _GEN_434 = 7'h31 == index ? valid_1_49 : _GEN_433; // @[cache.scala 37:{50,50}]
  wire  _GEN_435 = 7'h32 == index ? valid_1_50 : _GEN_434; // @[cache.scala 37:{50,50}]
  wire  _GEN_436 = 7'h33 == index ? valid_1_51 : _GEN_435; // @[cache.scala 37:{50,50}]
  wire  _GEN_437 = 7'h34 == index ? valid_1_52 : _GEN_436; // @[cache.scala 37:{50,50}]
  wire  _GEN_438 = 7'h35 == index ? valid_1_53 : _GEN_437; // @[cache.scala 37:{50,50}]
  wire  _GEN_439 = 7'h36 == index ? valid_1_54 : _GEN_438; // @[cache.scala 37:{50,50}]
  wire  _GEN_440 = 7'h37 == index ? valid_1_55 : _GEN_439; // @[cache.scala 37:{50,50}]
  wire  _GEN_441 = 7'h38 == index ? valid_1_56 : _GEN_440; // @[cache.scala 37:{50,50}]
  wire  _GEN_442 = 7'h39 == index ? valid_1_57 : _GEN_441; // @[cache.scala 37:{50,50}]
  wire  _GEN_443 = 7'h3a == index ? valid_1_58 : _GEN_442; // @[cache.scala 37:{50,50}]
  wire  _GEN_444 = 7'h3b == index ? valid_1_59 : _GEN_443; // @[cache.scala 37:{50,50}]
  wire  _GEN_445 = 7'h3c == index ? valid_1_60 : _GEN_444; // @[cache.scala 37:{50,50}]
  wire  _GEN_446 = 7'h3d == index ? valid_1_61 : _GEN_445; // @[cache.scala 37:{50,50}]
  wire  _GEN_447 = 7'h3e == index ? valid_1_62 : _GEN_446; // @[cache.scala 37:{50,50}]
  wire  _GEN_448 = 7'h3f == index ? valid_1_63 : _GEN_447; // @[cache.scala 37:{50,50}]
  wire  _GEN_449 = 7'h40 == index ? valid_1_64 : _GEN_448; // @[cache.scala 37:{50,50}]
  wire  _GEN_450 = 7'h41 == index ? valid_1_65 : _GEN_449; // @[cache.scala 37:{50,50}]
  wire  _GEN_451 = 7'h42 == index ? valid_1_66 : _GEN_450; // @[cache.scala 37:{50,50}]
  wire  _GEN_452 = 7'h43 == index ? valid_1_67 : _GEN_451; // @[cache.scala 37:{50,50}]
  wire  _GEN_453 = 7'h44 == index ? valid_1_68 : _GEN_452; // @[cache.scala 37:{50,50}]
  wire  _GEN_454 = 7'h45 == index ? valid_1_69 : _GEN_453; // @[cache.scala 37:{50,50}]
  wire  _GEN_455 = 7'h46 == index ? valid_1_70 : _GEN_454; // @[cache.scala 37:{50,50}]
  wire  _GEN_456 = 7'h47 == index ? valid_1_71 : _GEN_455; // @[cache.scala 37:{50,50}]
  wire  _GEN_457 = 7'h48 == index ? valid_1_72 : _GEN_456; // @[cache.scala 37:{50,50}]
  wire  _GEN_458 = 7'h49 == index ? valid_1_73 : _GEN_457; // @[cache.scala 37:{50,50}]
  wire  _GEN_459 = 7'h4a == index ? valid_1_74 : _GEN_458; // @[cache.scala 37:{50,50}]
  wire  _GEN_460 = 7'h4b == index ? valid_1_75 : _GEN_459; // @[cache.scala 37:{50,50}]
  wire  _GEN_461 = 7'h4c == index ? valid_1_76 : _GEN_460; // @[cache.scala 37:{50,50}]
  wire  _GEN_462 = 7'h4d == index ? valid_1_77 : _GEN_461; // @[cache.scala 37:{50,50}]
  wire  _GEN_463 = 7'h4e == index ? valid_1_78 : _GEN_462; // @[cache.scala 37:{50,50}]
  wire  _GEN_464 = 7'h4f == index ? valid_1_79 : _GEN_463; // @[cache.scala 37:{50,50}]
  wire  _GEN_465 = 7'h50 == index ? valid_1_80 : _GEN_464; // @[cache.scala 37:{50,50}]
  wire  _GEN_466 = 7'h51 == index ? valid_1_81 : _GEN_465; // @[cache.scala 37:{50,50}]
  wire  _GEN_467 = 7'h52 == index ? valid_1_82 : _GEN_466; // @[cache.scala 37:{50,50}]
  wire  _GEN_468 = 7'h53 == index ? valid_1_83 : _GEN_467; // @[cache.scala 37:{50,50}]
  wire  _GEN_469 = 7'h54 == index ? valid_1_84 : _GEN_468; // @[cache.scala 37:{50,50}]
  wire  _GEN_470 = 7'h55 == index ? valid_1_85 : _GEN_469; // @[cache.scala 37:{50,50}]
  wire  _GEN_471 = 7'h56 == index ? valid_1_86 : _GEN_470; // @[cache.scala 37:{50,50}]
  wire  _GEN_472 = 7'h57 == index ? valid_1_87 : _GEN_471; // @[cache.scala 37:{50,50}]
  wire  _GEN_473 = 7'h58 == index ? valid_1_88 : _GEN_472; // @[cache.scala 37:{50,50}]
  wire  _GEN_474 = 7'h59 == index ? valid_1_89 : _GEN_473; // @[cache.scala 37:{50,50}]
  wire  _GEN_475 = 7'h5a == index ? valid_1_90 : _GEN_474; // @[cache.scala 37:{50,50}]
  wire  _GEN_476 = 7'h5b == index ? valid_1_91 : _GEN_475; // @[cache.scala 37:{50,50}]
  wire  _GEN_477 = 7'h5c == index ? valid_1_92 : _GEN_476; // @[cache.scala 37:{50,50}]
  wire  _GEN_478 = 7'h5d == index ? valid_1_93 : _GEN_477; // @[cache.scala 37:{50,50}]
  wire  _GEN_479 = 7'h5e == index ? valid_1_94 : _GEN_478; // @[cache.scala 37:{50,50}]
  wire  _GEN_480 = 7'h5f == index ? valid_1_95 : _GEN_479; // @[cache.scala 37:{50,50}]
  wire  _GEN_481 = 7'h60 == index ? valid_1_96 : _GEN_480; // @[cache.scala 37:{50,50}]
  wire  _GEN_482 = 7'h61 == index ? valid_1_97 : _GEN_481; // @[cache.scala 37:{50,50}]
  wire  _GEN_483 = 7'h62 == index ? valid_1_98 : _GEN_482; // @[cache.scala 37:{50,50}]
  wire  _GEN_484 = 7'h63 == index ? valid_1_99 : _GEN_483; // @[cache.scala 37:{50,50}]
  wire  _GEN_485 = 7'h64 == index ? valid_1_100 : _GEN_484; // @[cache.scala 37:{50,50}]
  wire  _GEN_486 = 7'h65 == index ? valid_1_101 : _GEN_485; // @[cache.scala 37:{50,50}]
  wire  _GEN_487 = 7'h66 == index ? valid_1_102 : _GEN_486; // @[cache.scala 37:{50,50}]
  wire  _GEN_488 = 7'h67 == index ? valid_1_103 : _GEN_487; // @[cache.scala 37:{50,50}]
  wire  _GEN_489 = 7'h68 == index ? valid_1_104 : _GEN_488; // @[cache.scala 37:{50,50}]
  wire  _GEN_490 = 7'h69 == index ? valid_1_105 : _GEN_489; // @[cache.scala 37:{50,50}]
  wire  _GEN_491 = 7'h6a == index ? valid_1_106 : _GEN_490; // @[cache.scala 37:{50,50}]
  wire  _GEN_492 = 7'h6b == index ? valid_1_107 : _GEN_491; // @[cache.scala 37:{50,50}]
  wire  _GEN_493 = 7'h6c == index ? valid_1_108 : _GEN_492; // @[cache.scala 37:{50,50}]
  wire  _GEN_494 = 7'h6d == index ? valid_1_109 : _GEN_493; // @[cache.scala 37:{50,50}]
  wire  _GEN_495 = 7'h6e == index ? valid_1_110 : _GEN_494; // @[cache.scala 37:{50,50}]
  wire  _GEN_496 = 7'h6f == index ? valid_1_111 : _GEN_495; // @[cache.scala 37:{50,50}]
  wire  _GEN_497 = 7'h70 == index ? valid_1_112 : _GEN_496; // @[cache.scala 37:{50,50}]
  wire  _GEN_498 = 7'h71 == index ? valid_1_113 : _GEN_497; // @[cache.scala 37:{50,50}]
  wire  _GEN_499 = 7'h72 == index ? valid_1_114 : _GEN_498; // @[cache.scala 37:{50,50}]
  wire  _GEN_500 = 7'h73 == index ? valid_1_115 : _GEN_499; // @[cache.scala 37:{50,50}]
  wire  _GEN_501 = 7'h74 == index ? valid_1_116 : _GEN_500; // @[cache.scala 37:{50,50}]
  wire  _GEN_502 = 7'h75 == index ? valid_1_117 : _GEN_501; // @[cache.scala 37:{50,50}]
  wire  _GEN_503 = 7'h76 == index ? valid_1_118 : _GEN_502; // @[cache.scala 37:{50,50}]
  wire  _GEN_504 = 7'h77 == index ? valid_1_119 : _GEN_503; // @[cache.scala 37:{50,50}]
  wire  _GEN_505 = 7'h78 == index ? valid_1_120 : _GEN_504; // @[cache.scala 37:{50,50}]
  wire  _GEN_506 = 7'h79 == index ? valid_1_121 : _GEN_505; // @[cache.scala 37:{50,50}]
  wire  _GEN_507 = 7'h7a == index ? valid_1_122 : _GEN_506; // @[cache.scala 37:{50,50}]
  wire  _GEN_508 = 7'h7b == index ? valid_1_123 : _GEN_507; // @[cache.scala 37:{50,50}]
  wire  _GEN_509 = 7'h7c == index ? valid_1_124 : _GEN_508; // @[cache.scala 37:{50,50}]
  wire  _GEN_510 = 7'h7d == index ? valid_1_125 : _GEN_509; // @[cache.scala 37:{50,50}]
  wire  _GEN_511 = 7'h7e == index ? valid_1_126 : _GEN_510; // @[cache.scala 37:{50,50}]
  wire  _GEN_512 = 7'h7f == index ? valid_1_127 : _GEN_511; // @[cache.scala 37:{50,50}]
  wire  _GEN_513 = _GEN_384 == _GEN_7705 & _GEN_512 | way1_hit; // @[cache.scala 37:57 38:18 24:27]
  reg [1:0] state; // @[cache.scala 49:24]
  wire [1:0] _GEN_517 = io_from_ifu_rready ? 2'h0 : state; // @[cache.scala 49:24 60:41 61:27]
  wire [1:0] _GEN_518 = way1_hit ? _GEN_517 : 2'h2; // @[cache.scala 64:33 69:23]
  wire [1:0] _GEN_520 = io_from_axi_rvalid ? 2'h3 : state; // @[cache.scala 73:37 74:23 49:24]
  wire [63:0] _GEN_521 = io_from_axi_rvalid ? io_from_axi_rdata : receive_data; // @[cache.scala 76:37 77:30 27:31]
  wire [63:0] _GEN_522 = 7'h0 == index ? receive_data : ram_0_0; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_523 = 7'h1 == index ? receive_data : ram_0_1; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_524 = 7'h2 == index ? receive_data : ram_0_2; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_525 = 7'h3 == index ? receive_data : ram_0_3; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_526 = 7'h4 == index ? receive_data : ram_0_4; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_527 = 7'h5 == index ? receive_data : ram_0_5; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_528 = 7'h6 == index ? receive_data : ram_0_6; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_529 = 7'h7 == index ? receive_data : ram_0_7; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_530 = 7'h8 == index ? receive_data : ram_0_8; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_531 = 7'h9 == index ? receive_data : ram_0_9; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_532 = 7'ha == index ? receive_data : ram_0_10; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_533 = 7'hb == index ? receive_data : ram_0_11; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_534 = 7'hc == index ? receive_data : ram_0_12; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_535 = 7'hd == index ? receive_data : ram_0_13; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_536 = 7'he == index ? receive_data : ram_0_14; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_537 = 7'hf == index ? receive_data : ram_0_15; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_538 = 7'h10 == index ? receive_data : ram_0_16; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_539 = 7'h11 == index ? receive_data : ram_0_17; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_540 = 7'h12 == index ? receive_data : ram_0_18; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_541 = 7'h13 == index ? receive_data : ram_0_19; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_542 = 7'h14 == index ? receive_data : ram_0_20; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_543 = 7'h15 == index ? receive_data : ram_0_21; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_544 = 7'h16 == index ? receive_data : ram_0_22; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_545 = 7'h17 == index ? receive_data : ram_0_23; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_546 = 7'h18 == index ? receive_data : ram_0_24; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_547 = 7'h19 == index ? receive_data : ram_0_25; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_548 = 7'h1a == index ? receive_data : ram_0_26; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_549 = 7'h1b == index ? receive_data : ram_0_27; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_550 = 7'h1c == index ? receive_data : ram_0_28; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_551 = 7'h1d == index ? receive_data : ram_0_29; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_552 = 7'h1e == index ? receive_data : ram_0_30; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_553 = 7'h1f == index ? receive_data : ram_0_31; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_554 = 7'h20 == index ? receive_data : ram_0_32; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_555 = 7'h21 == index ? receive_data : ram_0_33; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_556 = 7'h22 == index ? receive_data : ram_0_34; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_557 = 7'h23 == index ? receive_data : ram_0_35; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_558 = 7'h24 == index ? receive_data : ram_0_36; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_559 = 7'h25 == index ? receive_data : ram_0_37; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_560 = 7'h26 == index ? receive_data : ram_0_38; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_561 = 7'h27 == index ? receive_data : ram_0_39; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_562 = 7'h28 == index ? receive_data : ram_0_40; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_563 = 7'h29 == index ? receive_data : ram_0_41; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_564 = 7'h2a == index ? receive_data : ram_0_42; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_565 = 7'h2b == index ? receive_data : ram_0_43; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_566 = 7'h2c == index ? receive_data : ram_0_44; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_567 = 7'h2d == index ? receive_data : ram_0_45; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_568 = 7'h2e == index ? receive_data : ram_0_46; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_569 = 7'h2f == index ? receive_data : ram_0_47; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_570 = 7'h30 == index ? receive_data : ram_0_48; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_571 = 7'h31 == index ? receive_data : ram_0_49; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_572 = 7'h32 == index ? receive_data : ram_0_50; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_573 = 7'h33 == index ? receive_data : ram_0_51; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_574 = 7'h34 == index ? receive_data : ram_0_52; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_575 = 7'h35 == index ? receive_data : ram_0_53; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_576 = 7'h36 == index ? receive_data : ram_0_54; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_577 = 7'h37 == index ? receive_data : ram_0_55; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_578 = 7'h38 == index ? receive_data : ram_0_56; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_579 = 7'h39 == index ? receive_data : ram_0_57; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_580 = 7'h3a == index ? receive_data : ram_0_58; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_581 = 7'h3b == index ? receive_data : ram_0_59; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_582 = 7'h3c == index ? receive_data : ram_0_60; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_583 = 7'h3d == index ? receive_data : ram_0_61; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_584 = 7'h3e == index ? receive_data : ram_0_62; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_585 = 7'h3f == index ? receive_data : ram_0_63; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_586 = 7'h40 == index ? receive_data : ram_0_64; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_587 = 7'h41 == index ? receive_data : ram_0_65; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_588 = 7'h42 == index ? receive_data : ram_0_66; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_589 = 7'h43 == index ? receive_data : ram_0_67; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_590 = 7'h44 == index ? receive_data : ram_0_68; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_591 = 7'h45 == index ? receive_data : ram_0_69; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_592 = 7'h46 == index ? receive_data : ram_0_70; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_593 = 7'h47 == index ? receive_data : ram_0_71; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_594 = 7'h48 == index ? receive_data : ram_0_72; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_595 = 7'h49 == index ? receive_data : ram_0_73; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_596 = 7'h4a == index ? receive_data : ram_0_74; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_597 = 7'h4b == index ? receive_data : ram_0_75; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_598 = 7'h4c == index ? receive_data : ram_0_76; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_599 = 7'h4d == index ? receive_data : ram_0_77; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_600 = 7'h4e == index ? receive_data : ram_0_78; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_601 = 7'h4f == index ? receive_data : ram_0_79; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_602 = 7'h50 == index ? receive_data : ram_0_80; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_603 = 7'h51 == index ? receive_data : ram_0_81; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_604 = 7'h52 == index ? receive_data : ram_0_82; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_605 = 7'h53 == index ? receive_data : ram_0_83; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_606 = 7'h54 == index ? receive_data : ram_0_84; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_607 = 7'h55 == index ? receive_data : ram_0_85; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_608 = 7'h56 == index ? receive_data : ram_0_86; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_609 = 7'h57 == index ? receive_data : ram_0_87; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_610 = 7'h58 == index ? receive_data : ram_0_88; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_611 = 7'h59 == index ? receive_data : ram_0_89; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_612 = 7'h5a == index ? receive_data : ram_0_90; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_613 = 7'h5b == index ? receive_data : ram_0_91; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_614 = 7'h5c == index ? receive_data : ram_0_92; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_615 = 7'h5d == index ? receive_data : ram_0_93; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_616 = 7'h5e == index ? receive_data : ram_0_94; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_617 = 7'h5f == index ? receive_data : ram_0_95; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_618 = 7'h60 == index ? receive_data : ram_0_96; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_619 = 7'h61 == index ? receive_data : ram_0_97; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_620 = 7'h62 == index ? receive_data : ram_0_98; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_621 = 7'h63 == index ? receive_data : ram_0_99; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_622 = 7'h64 == index ? receive_data : ram_0_100; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_623 = 7'h65 == index ? receive_data : ram_0_101; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_624 = 7'h66 == index ? receive_data : ram_0_102; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_625 = 7'h67 == index ? receive_data : ram_0_103; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_626 = 7'h68 == index ? receive_data : ram_0_104; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_627 = 7'h69 == index ? receive_data : ram_0_105; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_628 = 7'h6a == index ? receive_data : ram_0_106; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_629 = 7'h6b == index ? receive_data : ram_0_107; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_630 = 7'h6c == index ? receive_data : ram_0_108; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_631 = 7'h6d == index ? receive_data : ram_0_109; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_632 = 7'h6e == index ? receive_data : ram_0_110; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_633 = 7'h6f == index ? receive_data : ram_0_111; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_634 = 7'h70 == index ? receive_data : ram_0_112; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_635 = 7'h71 == index ? receive_data : ram_0_113; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_636 = 7'h72 == index ? receive_data : ram_0_114; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_637 = 7'h73 == index ? receive_data : ram_0_115; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_638 = 7'h74 == index ? receive_data : ram_0_116; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_639 = 7'h75 == index ? receive_data : ram_0_117; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_640 = 7'h76 == index ? receive_data : ram_0_118; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_641 = 7'h77 == index ? receive_data : ram_0_119; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_642 = 7'h78 == index ? receive_data : ram_0_120; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_643 = 7'h79 == index ? receive_data : ram_0_121; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_644 = 7'h7a == index ? receive_data : ram_0_122; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_645 = 7'h7b == index ? receive_data : ram_0_123; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_646 = 7'h7c == index ? receive_data : ram_0_124; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_647 = 7'h7d == index ? receive_data : ram_0_125; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_648 = 7'h7e == index ? receive_data : ram_0_126; // @[cache.scala 17:24 83:{30,30}]
  wire [63:0] _GEN_649 = 7'h7f == index ? receive_data : ram_0_127; // @[cache.scala 17:24 83:{30,30}]
  wire [31:0] _GEN_650 = 7'h0 == index ? _GEN_7705 : tag_0_0; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_651 = 7'h1 == index ? _GEN_7705 : tag_0_1; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_652 = 7'h2 == index ? _GEN_7705 : tag_0_2; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_653 = 7'h3 == index ? _GEN_7705 : tag_0_3; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_654 = 7'h4 == index ? _GEN_7705 : tag_0_4; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_655 = 7'h5 == index ? _GEN_7705 : tag_0_5; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_656 = 7'h6 == index ? _GEN_7705 : tag_0_6; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_657 = 7'h7 == index ? _GEN_7705 : tag_0_7; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_658 = 7'h8 == index ? _GEN_7705 : tag_0_8; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_659 = 7'h9 == index ? _GEN_7705 : tag_0_9; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_660 = 7'ha == index ? _GEN_7705 : tag_0_10; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_661 = 7'hb == index ? _GEN_7705 : tag_0_11; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_662 = 7'hc == index ? _GEN_7705 : tag_0_12; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_663 = 7'hd == index ? _GEN_7705 : tag_0_13; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_664 = 7'he == index ? _GEN_7705 : tag_0_14; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_665 = 7'hf == index ? _GEN_7705 : tag_0_15; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_666 = 7'h10 == index ? _GEN_7705 : tag_0_16; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_667 = 7'h11 == index ? _GEN_7705 : tag_0_17; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_668 = 7'h12 == index ? _GEN_7705 : tag_0_18; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_669 = 7'h13 == index ? _GEN_7705 : tag_0_19; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_670 = 7'h14 == index ? _GEN_7705 : tag_0_20; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_671 = 7'h15 == index ? _GEN_7705 : tag_0_21; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_672 = 7'h16 == index ? _GEN_7705 : tag_0_22; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_673 = 7'h17 == index ? _GEN_7705 : tag_0_23; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_674 = 7'h18 == index ? _GEN_7705 : tag_0_24; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_675 = 7'h19 == index ? _GEN_7705 : tag_0_25; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_676 = 7'h1a == index ? _GEN_7705 : tag_0_26; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_677 = 7'h1b == index ? _GEN_7705 : tag_0_27; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_678 = 7'h1c == index ? _GEN_7705 : tag_0_28; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_679 = 7'h1d == index ? _GEN_7705 : tag_0_29; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_680 = 7'h1e == index ? _GEN_7705 : tag_0_30; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_681 = 7'h1f == index ? _GEN_7705 : tag_0_31; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_682 = 7'h20 == index ? _GEN_7705 : tag_0_32; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_683 = 7'h21 == index ? _GEN_7705 : tag_0_33; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_684 = 7'h22 == index ? _GEN_7705 : tag_0_34; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_685 = 7'h23 == index ? _GEN_7705 : tag_0_35; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_686 = 7'h24 == index ? _GEN_7705 : tag_0_36; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_687 = 7'h25 == index ? _GEN_7705 : tag_0_37; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_688 = 7'h26 == index ? _GEN_7705 : tag_0_38; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_689 = 7'h27 == index ? _GEN_7705 : tag_0_39; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_690 = 7'h28 == index ? _GEN_7705 : tag_0_40; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_691 = 7'h29 == index ? _GEN_7705 : tag_0_41; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_692 = 7'h2a == index ? _GEN_7705 : tag_0_42; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_693 = 7'h2b == index ? _GEN_7705 : tag_0_43; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_694 = 7'h2c == index ? _GEN_7705 : tag_0_44; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_695 = 7'h2d == index ? _GEN_7705 : tag_0_45; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_696 = 7'h2e == index ? _GEN_7705 : tag_0_46; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_697 = 7'h2f == index ? _GEN_7705 : tag_0_47; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_698 = 7'h30 == index ? _GEN_7705 : tag_0_48; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_699 = 7'h31 == index ? _GEN_7705 : tag_0_49; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_700 = 7'h32 == index ? _GEN_7705 : tag_0_50; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_701 = 7'h33 == index ? _GEN_7705 : tag_0_51; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_702 = 7'h34 == index ? _GEN_7705 : tag_0_52; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_703 = 7'h35 == index ? _GEN_7705 : tag_0_53; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_704 = 7'h36 == index ? _GEN_7705 : tag_0_54; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_705 = 7'h37 == index ? _GEN_7705 : tag_0_55; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_706 = 7'h38 == index ? _GEN_7705 : tag_0_56; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_707 = 7'h39 == index ? _GEN_7705 : tag_0_57; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_708 = 7'h3a == index ? _GEN_7705 : tag_0_58; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_709 = 7'h3b == index ? _GEN_7705 : tag_0_59; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_710 = 7'h3c == index ? _GEN_7705 : tag_0_60; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_711 = 7'h3d == index ? _GEN_7705 : tag_0_61; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_712 = 7'h3e == index ? _GEN_7705 : tag_0_62; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_713 = 7'h3f == index ? _GEN_7705 : tag_0_63; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_714 = 7'h40 == index ? _GEN_7705 : tag_0_64; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_715 = 7'h41 == index ? _GEN_7705 : tag_0_65; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_716 = 7'h42 == index ? _GEN_7705 : tag_0_66; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_717 = 7'h43 == index ? _GEN_7705 : tag_0_67; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_718 = 7'h44 == index ? _GEN_7705 : tag_0_68; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_719 = 7'h45 == index ? _GEN_7705 : tag_0_69; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_720 = 7'h46 == index ? _GEN_7705 : tag_0_70; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_721 = 7'h47 == index ? _GEN_7705 : tag_0_71; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_722 = 7'h48 == index ? _GEN_7705 : tag_0_72; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_723 = 7'h49 == index ? _GEN_7705 : tag_0_73; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_724 = 7'h4a == index ? _GEN_7705 : tag_0_74; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_725 = 7'h4b == index ? _GEN_7705 : tag_0_75; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_726 = 7'h4c == index ? _GEN_7705 : tag_0_76; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_727 = 7'h4d == index ? _GEN_7705 : tag_0_77; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_728 = 7'h4e == index ? _GEN_7705 : tag_0_78; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_729 = 7'h4f == index ? _GEN_7705 : tag_0_79; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_730 = 7'h50 == index ? _GEN_7705 : tag_0_80; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_731 = 7'h51 == index ? _GEN_7705 : tag_0_81; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_732 = 7'h52 == index ? _GEN_7705 : tag_0_82; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_733 = 7'h53 == index ? _GEN_7705 : tag_0_83; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_734 = 7'h54 == index ? _GEN_7705 : tag_0_84; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_735 = 7'h55 == index ? _GEN_7705 : tag_0_85; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_736 = 7'h56 == index ? _GEN_7705 : tag_0_86; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_737 = 7'h57 == index ? _GEN_7705 : tag_0_87; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_738 = 7'h58 == index ? _GEN_7705 : tag_0_88; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_739 = 7'h59 == index ? _GEN_7705 : tag_0_89; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_740 = 7'h5a == index ? _GEN_7705 : tag_0_90; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_741 = 7'h5b == index ? _GEN_7705 : tag_0_91; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_742 = 7'h5c == index ? _GEN_7705 : tag_0_92; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_743 = 7'h5d == index ? _GEN_7705 : tag_0_93; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_744 = 7'h5e == index ? _GEN_7705 : tag_0_94; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_745 = 7'h5f == index ? _GEN_7705 : tag_0_95; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_746 = 7'h60 == index ? _GEN_7705 : tag_0_96; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_747 = 7'h61 == index ? _GEN_7705 : tag_0_97; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_748 = 7'h62 == index ? _GEN_7705 : tag_0_98; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_749 = 7'h63 == index ? _GEN_7705 : tag_0_99; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_750 = 7'h64 == index ? _GEN_7705 : tag_0_100; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_751 = 7'h65 == index ? _GEN_7705 : tag_0_101; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_752 = 7'h66 == index ? _GEN_7705 : tag_0_102; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_753 = 7'h67 == index ? _GEN_7705 : tag_0_103; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_754 = 7'h68 == index ? _GEN_7705 : tag_0_104; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_755 = 7'h69 == index ? _GEN_7705 : tag_0_105; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_756 = 7'h6a == index ? _GEN_7705 : tag_0_106; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_757 = 7'h6b == index ? _GEN_7705 : tag_0_107; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_758 = 7'h6c == index ? _GEN_7705 : tag_0_108; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_759 = 7'h6d == index ? _GEN_7705 : tag_0_109; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_760 = 7'h6e == index ? _GEN_7705 : tag_0_110; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_761 = 7'h6f == index ? _GEN_7705 : tag_0_111; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_762 = 7'h70 == index ? _GEN_7705 : tag_0_112; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_763 = 7'h71 == index ? _GEN_7705 : tag_0_113; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_764 = 7'h72 == index ? _GEN_7705 : tag_0_114; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_765 = 7'h73 == index ? _GEN_7705 : tag_0_115; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_766 = 7'h74 == index ? _GEN_7705 : tag_0_116; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_767 = 7'h75 == index ? _GEN_7705 : tag_0_117; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_768 = 7'h76 == index ? _GEN_7705 : tag_0_118; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_769 = 7'h77 == index ? _GEN_7705 : tag_0_119; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_770 = 7'h78 == index ? _GEN_7705 : tag_0_120; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_771 = 7'h79 == index ? _GEN_7705 : tag_0_121; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_772 = 7'h7a == index ? _GEN_7705 : tag_0_122; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_773 = 7'h7b == index ? _GEN_7705 : tag_0_123; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_774 = 7'h7c == index ? _GEN_7705 : tag_0_124; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_775 = 7'h7d == index ? _GEN_7705 : tag_0_125; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_776 = 7'h7e == index ? _GEN_7705 : tag_0_126; // @[cache.scala 19:24 84:{30,30}]
  wire [31:0] _GEN_777 = 7'h7f == index ? _GEN_7705 : tag_0_127; // @[cache.scala 19:24 84:{30,30}]
  wire  _GEN_7709 = 7'h0 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_778 = 7'h0 == index | valid_0_0; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7711 = 7'h1 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_779 = 7'h1 == index | valid_0_1; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7713 = 7'h2 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_780 = 7'h2 == index | valid_0_2; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7717 = 7'h3 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_781 = 7'h3 == index | valid_0_3; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7726 = 7'h4 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_782 = 7'h4 == index | valid_0_4; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7728 = 7'h5 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_783 = 7'h5 == index | valid_0_5; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7730 = 7'h6 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_784 = 7'h6 == index | valid_0_6; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7732 = 7'h7 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_785 = 7'h7 == index | valid_0_7; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7737 = 7'h8 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_786 = 7'h8 == index | valid_0_8; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7738 = 7'h9 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_787 = 7'h9 == index | valid_0_9; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7739 = 7'ha == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_788 = 7'ha == index | valid_0_10; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7740 = 7'hb == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_789 = 7'hb == index | valid_0_11; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7741 = 7'hc == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_790 = 7'hc == index | valid_0_12; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7742 = 7'hd == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_791 = 7'hd == index | valid_0_13; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7743 = 7'he == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_792 = 7'he == index | valid_0_14; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7744 = 7'hf == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_793 = 7'hf == index | valid_0_15; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7745 = 7'h10 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_794 = 7'h10 == index | valid_0_16; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7746 = 7'h11 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_795 = 7'h11 == index | valid_0_17; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7747 = 7'h12 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_796 = 7'h12 == index | valid_0_18; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7748 = 7'h13 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_797 = 7'h13 == index | valid_0_19; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7749 = 7'h14 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_798 = 7'h14 == index | valid_0_20; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7750 = 7'h15 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_799 = 7'h15 == index | valid_0_21; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7751 = 7'h16 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_800 = 7'h16 == index | valid_0_22; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7752 = 7'h17 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_801 = 7'h17 == index | valid_0_23; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7753 = 7'h18 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_802 = 7'h18 == index | valid_0_24; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7754 = 7'h19 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_803 = 7'h19 == index | valid_0_25; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7755 = 7'h1a == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_804 = 7'h1a == index | valid_0_26; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7756 = 7'h1b == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_805 = 7'h1b == index | valid_0_27; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7757 = 7'h1c == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_806 = 7'h1c == index | valid_0_28; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7758 = 7'h1d == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_807 = 7'h1d == index | valid_0_29; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7759 = 7'h1e == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_808 = 7'h1e == index | valid_0_30; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7760 = 7'h1f == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_809 = 7'h1f == index | valid_0_31; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7761 = 7'h20 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_810 = 7'h20 == index | valid_0_32; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7762 = 7'h21 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_811 = 7'h21 == index | valid_0_33; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7763 = 7'h22 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_812 = 7'h22 == index | valid_0_34; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7764 = 7'h23 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_813 = 7'h23 == index | valid_0_35; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7765 = 7'h24 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_814 = 7'h24 == index | valid_0_36; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7766 = 7'h25 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_815 = 7'h25 == index | valid_0_37; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7767 = 7'h26 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_816 = 7'h26 == index | valid_0_38; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7768 = 7'h27 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_817 = 7'h27 == index | valid_0_39; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7769 = 7'h28 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_818 = 7'h28 == index | valid_0_40; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7770 = 7'h29 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_819 = 7'h29 == index | valid_0_41; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7771 = 7'h2a == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_820 = 7'h2a == index | valid_0_42; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7772 = 7'h2b == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_821 = 7'h2b == index | valid_0_43; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7773 = 7'h2c == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_822 = 7'h2c == index | valid_0_44; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7774 = 7'h2d == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_823 = 7'h2d == index | valid_0_45; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7775 = 7'h2e == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_824 = 7'h2e == index | valid_0_46; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7776 = 7'h2f == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_825 = 7'h2f == index | valid_0_47; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7777 = 7'h30 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_826 = 7'h30 == index | valid_0_48; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7778 = 7'h31 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_827 = 7'h31 == index | valid_0_49; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7779 = 7'h32 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_828 = 7'h32 == index | valid_0_50; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7780 = 7'h33 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_829 = 7'h33 == index | valid_0_51; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7781 = 7'h34 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_830 = 7'h34 == index | valid_0_52; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7782 = 7'h35 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_831 = 7'h35 == index | valid_0_53; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7783 = 7'h36 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_832 = 7'h36 == index | valid_0_54; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7784 = 7'h37 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_833 = 7'h37 == index | valid_0_55; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7785 = 7'h38 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_834 = 7'h38 == index | valid_0_56; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7786 = 7'h39 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_835 = 7'h39 == index | valid_0_57; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7787 = 7'h3a == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_836 = 7'h3a == index | valid_0_58; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7788 = 7'h3b == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_837 = 7'h3b == index | valid_0_59; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7789 = 7'h3c == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_838 = 7'h3c == index | valid_0_60; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7790 = 7'h3d == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_839 = 7'h3d == index | valid_0_61; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7791 = 7'h3e == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_840 = 7'h3e == index | valid_0_62; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7792 = 7'h3f == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_841 = 7'h3f == index | valid_0_63; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7793 = 7'h40 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_842 = 7'h40 == index | valid_0_64; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7794 = 7'h41 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_843 = 7'h41 == index | valid_0_65; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7795 = 7'h42 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_844 = 7'h42 == index | valid_0_66; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7796 = 7'h43 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_845 = 7'h43 == index | valid_0_67; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7797 = 7'h44 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_846 = 7'h44 == index | valid_0_68; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7798 = 7'h45 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_847 = 7'h45 == index | valid_0_69; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7799 = 7'h46 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_848 = 7'h46 == index | valid_0_70; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7800 = 7'h47 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_849 = 7'h47 == index | valid_0_71; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7801 = 7'h48 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_850 = 7'h48 == index | valid_0_72; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7802 = 7'h49 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_851 = 7'h49 == index | valid_0_73; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7803 = 7'h4a == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_852 = 7'h4a == index | valid_0_74; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7804 = 7'h4b == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_853 = 7'h4b == index | valid_0_75; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7805 = 7'h4c == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_854 = 7'h4c == index | valid_0_76; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7806 = 7'h4d == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_855 = 7'h4d == index | valid_0_77; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7807 = 7'h4e == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_856 = 7'h4e == index | valid_0_78; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7808 = 7'h4f == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_857 = 7'h4f == index | valid_0_79; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7809 = 7'h50 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_858 = 7'h50 == index | valid_0_80; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7810 = 7'h51 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_859 = 7'h51 == index | valid_0_81; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7811 = 7'h52 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_860 = 7'h52 == index | valid_0_82; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7812 = 7'h53 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_861 = 7'h53 == index | valid_0_83; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7813 = 7'h54 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_862 = 7'h54 == index | valid_0_84; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7814 = 7'h55 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_863 = 7'h55 == index | valid_0_85; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7815 = 7'h56 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_864 = 7'h56 == index | valid_0_86; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7816 = 7'h57 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_865 = 7'h57 == index | valid_0_87; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7817 = 7'h58 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_866 = 7'h58 == index | valid_0_88; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7818 = 7'h59 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_867 = 7'h59 == index | valid_0_89; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7819 = 7'h5a == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_868 = 7'h5a == index | valid_0_90; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7820 = 7'h5b == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_869 = 7'h5b == index | valid_0_91; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7821 = 7'h5c == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_870 = 7'h5c == index | valid_0_92; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7822 = 7'h5d == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_871 = 7'h5d == index | valid_0_93; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7823 = 7'h5e == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_872 = 7'h5e == index | valid_0_94; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7824 = 7'h5f == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_873 = 7'h5f == index | valid_0_95; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7825 = 7'h60 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_874 = 7'h60 == index | valid_0_96; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7826 = 7'h61 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_875 = 7'h61 == index | valid_0_97; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7827 = 7'h62 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_876 = 7'h62 == index | valid_0_98; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7828 = 7'h63 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_877 = 7'h63 == index | valid_0_99; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7829 = 7'h64 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_878 = 7'h64 == index | valid_0_100; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7830 = 7'h65 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_879 = 7'h65 == index | valid_0_101; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7831 = 7'h66 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_880 = 7'h66 == index | valid_0_102; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7832 = 7'h67 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_881 = 7'h67 == index | valid_0_103; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7833 = 7'h68 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_882 = 7'h68 == index | valid_0_104; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7834 = 7'h69 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_883 = 7'h69 == index | valid_0_105; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7835 = 7'h6a == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_884 = 7'h6a == index | valid_0_106; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7836 = 7'h6b == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_885 = 7'h6b == index | valid_0_107; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7837 = 7'h6c == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_886 = 7'h6c == index | valid_0_108; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7838 = 7'h6d == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_887 = 7'h6d == index | valid_0_109; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7839 = 7'h6e == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_888 = 7'h6e == index | valid_0_110; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7840 = 7'h6f == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_889 = 7'h6f == index | valid_0_111; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7841 = 7'h70 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_890 = 7'h70 == index | valid_0_112; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7842 = 7'h71 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_891 = 7'h71 == index | valid_0_113; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7843 = 7'h72 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_892 = 7'h72 == index | valid_0_114; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7844 = 7'h73 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_893 = 7'h73 == index | valid_0_115; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7845 = 7'h74 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_894 = 7'h74 == index | valid_0_116; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7846 = 7'h75 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_895 = 7'h75 == index | valid_0_117; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7847 = 7'h76 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_896 = 7'h76 == index | valid_0_118; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7848 = 7'h77 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_897 = 7'h77 == index | valid_0_119; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7849 = 7'h78 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_898 = 7'h78 == index | valid_0_120; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7850 = 7'h79 == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_899 = 7'h79 == index | valid_0_121; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7851 = 7'h7a == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_900 = 7'h7a == index | valid_0_122; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7852 = 7'h7b == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_901 = 7'h7b == index | valid_0_123; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7853 = 7'h7c == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_902 = 7'h7c == index | valid_0_124; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7854 = 7'h7d == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_903 = 7'h7d == index | valid_0_125; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7855 = 7'h7e == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_904 = 7'h7e == index | valid_0_126; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_7856 = 7'h7f == index; // @[cache.scala 21:26 85:{32,32}]
  wire  _GEN_905 = 7'h7f == index | valid_0_127; // @[cache.scala 21:26 85:{32,32}]
  wire [63:0] _GEN_906 = 7'h0 == index ? receive_data : ram_1_0; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_907 = 7'h1 == index ? receive_data : ram_1_1; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_908 = 7'h2 == index ? receive_data : ram_1_2; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_909 = 7'h3 == index ? receive_data : ram_1_3; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_910 = 7'h4 == index ? receive_data : ram_1_4; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_911 = 7'h5 == index ? receive_data : ram_1_5; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_912 = 7'h6 == index ? receive_data : ram_1_6; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_913 = 7'h7 == index ? receive_data : ram_1_7; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_914 = 7'h8 == index ? receive_data : ram_1_8; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_915 = 7'h9 == index ? receive_data : ram_1_9; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_916 = 7'ha == index ? receive_data : ram_1_10; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_917 = 7'hb == index ? receive_data : ram_1_11; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_918 = 7'hc == index ? receive_data : ram_1_12; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_919 = 7'hd == index ? receive_data : ram_1_13; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_920 = 7'he == index ? receive_data : ram_1_14; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_921 = 7'hf == index ? receive_data : ram_1_15; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_922 = 7'h10 == index ? receive_data : ram_1_16; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_923 = 7'h11 == index ? receive_data : ram_1_17; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_924 = 7'h12 == index ? receive_data : ram_1_18; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_925 = 7'h13 == index ? receive_data : ram_1_19; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_926 = 7'h14 == index ? receive_data : ram_1_20; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_927 = 7'h15 == index ? receive_data : ram_1_21; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_928 = 7'h16 == index ? receive_data : ram_1_22; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_929 = 7'h17 == index ? receive_data : ram_1_23; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_930 = 7'h18 == index ? receive_data : ram_1_24; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_931 = 7'h19 == index ? receive_data : ram_1_25; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_932 = 7'h1a == index ? receive_data : ram_1_26; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_933 = 7'h1b == index ? receive_data : ram_1_27; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_934 = 7'h1c == index ? receive_data : ram_1_28; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_935 = 7'h1d == index ? receive_data : ram_1_29; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_936 = 7'h1e == index ? receive_data : ram_1_30; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_937 = 7'h1f == index ? receive_data : ram_1_31; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_938 = 7'h20 == index ? receive_data : ram_1_32; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_939 = 7'h21 == index ? receive_data : ram_1_33; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_940 = 7'h22 == index ? receive_data : ram_1_34; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_941 = 7'h23 == index ? receive_data : ram_1_35; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_942 = 7'h24 == index ? receive_data : ram_1_36; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_943 = 7'h25 == index ? receive_data : ram_1_37; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_944 = 7'h26 == index ? receive_data : ram_1_38; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_945 = 7'h27 == index ? receive_data : ram_1_39; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_946 = 7'h28 == index ? receive_data : ram_1_40; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_947 = 7'h29 == index ? receive_data : ram_1_41; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_948 = 7'h2a == index ? receive_data : ram_1_42; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_949 = 7'h2b == index ? receive_data : ram_1_43; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_950 = 7'h2c == index ? receive_data : ram_1_44; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_951 = 7'h2d == index ? receive_data : ram_1_45; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_952 = 7'h2e == index ? receive_data : ram_1_46; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_953 = 7'h2f == index ? receive_data : ram_1_47; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_954 = 7'h30 == index ? receive_data : ram_1_48; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_955 = 7'h31 == index ? receive_data : ram_1_49; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_956 = 7'h32 == index ? receive_data : ram_1_50; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_957 = 7'h33 == index ? receive_data : ram_1_51; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_958 = 7'h34 == index ? receive_data : ram_1_52; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_959 = 7'h35 == index ? receive_data : ram_1_53; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_960 = 7'h36 == index ? receive_data : ram_1_54; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_961 = 7'h37 == index ? receive_data : ram_1_55; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_962 = 7'h38 == index ? receive_data : ram_1_56; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_963 = 7'h39 == index ? receive_data : ram_1_57; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_964 = 7'h3a == index ? receive_data : ram_1_58; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_965 = 7'h3b == index ? receive_data : ram_1_59; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_966 = 7'h3c == index ? receive_data : ram_1_60; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_967 = 7'h3d == index ? receive_data : ram_1_61; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_968 = 7'h3e == index ? receive_data : ram_1_62; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_969 = 7'h3f == index ? receive_data : ram_1_63; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_970 = 7'h40 == index ? receive_data : ram_1_64; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_971 = 7'h41 == index ? receive_data : ram_1_65; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_972 = 7'h42 == index ? receive_data : ram_1_66; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_973 = 7'h43 == index ? receive_data : ram_1_67; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_974 = 7'h44 == index ? receive_data : ram_1_68; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_975 = 7'h45 == index ? receive_data : ram_1_69; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_976 = 7'h46 == index ? receive_data : ram_1_70; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_977 = 7'h47 == index ? receive_data : ram_1_71; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_978 = 7'h48 == index ? receive_data : ram_1_72; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_979 = 7'h49 == index ? receive_data : ram_1_73; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_980 = 7'h4a == index ? receive_data : ram_1_74; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_981 = 7'h4b == index ? receive_data : ram_1_75; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_982 = 7'h4c == index ? receive_data : ram_1_76; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_983 = 7'h4d == index ? receive_data : ram_1_77; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_984 = 7'h4e == index ? receive_data : ram_1_78; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_985 = 7'h4f == index ? receive_data : ram_1_79; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_986 = 7'h50 == index ? receive_data : ram_1_80; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_987 = 7'h51 == index ? receive_data : ram_1_81; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_988 = 7'h52 == index ? receive_data : ram_1_82; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_989 = 7'h53 == index ? receive_data : ram_1_83; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_990 = 7'h54 == index ? receive_data : ram_1_84; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_991 = 7'h55 == index ? receive_data : ram_1_85; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_992 = 7'h56 == index ? receive_data : ram_1_86; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_993 = 7'h57 == index ? receive_data : ram_1_87; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_994 = 7'h58 == index ? receive_data : ram_1_88; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_995 = 7'h59 == index ? receive_data : ram_1_89; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_996 = 7'h5a == index ? receive_data : ram_1_90; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_997 = 7'h5b == index ? receive_data : ram_1_91; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_998 = 7'h5c == index ? receive_data : ram_1_92; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_999 = 7'h5d == index ? receive_data : ram_1_93; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1000 = 7'h5e == index ? receive_data : ram_1_94; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1001 = 7'h5f == index ? receive_data : ram_1_95; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1002 = 7'h60 == index ? receive_data : ram_1_96; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1003 = 7'h61 == index ? receive_data : ram_1_97; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1004 = 7'h62 == index ? receive_data : ram_1_98; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1005 = 7'h63 == index ? receive_data : ram_1_99; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1006 = 7'h64 == index ? receive_data : ram_1_100; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1007 = 7'h65 == index ? receive_data : ram_1_101; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1008 = 7'h66 == index ? receive_data : ram_1_102; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1009 = 7'h67 == index ? receive_data : ram_1_103; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1010 = 7'h68 == index ? receive_data : ram_1_104; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1011 = 7'h69 == index ? receive_data : ram_1_105; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1012 = 7'h6a == index ? receive_data : ram_1_106; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1013 = 7'h6b == index ? receive_data : ram_1_107; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1014 = 7'h6c == index ? receive_data : ram_1_108; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1015 = 7'h6d == index ? receive_data : ram_1_109; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1016 = 7'h6e == index ? receive_data : ram_1_110; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1017 = 7'h6f == index ? receive_data : ram_1_111; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1018 = 7'h70 == index ? receive_data : ram_1_112; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1019 = 7'h71 == index ? receive_data : ram_1_113; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1020 = 7'h72 == index ? receive_data : ram_1_114; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1021 = 7'h73 == index ? receive_data : ram_1_115; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1022 = 7'h74 == index ? receive_data : ram_1_116; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1023 = 7'h75 == index ? receive_data : ram_1_117; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1024 = 7'h76 == index ? receive_data : ram_1_118; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1025 = 7'h77 == index ? receive_data : ram_1_119; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1026 = 7'h78 == index ? receive_data : ram_1_120; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1027 = 7'h79 == index ? receive_data : ram_1_121; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1028 = 7'h7a == index ? receive_data : ram_1_122; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1029 = 7'h7b == index ? receive_data : ram_1_123; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1030 = 7'h7c == index ? receive_data : ram_1_124; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1031 = 7'h7d == index ? receive_data : ram_1_125; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1032 = 7'h7e == index ? receive_data : ram_1_126; // @[cache.scala 18:24 88:{30,30}]
  wire [63:0] _GEN_1033 = 7'h7f == index ? receive_data : ram_1_127; // @[cache.scala 18:24 88:{30,30}]
  wire [31:0] _GEN_1034 = 7'h0 == index ? _GEN_7705 : tag_1_0; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1035 = 7'h1 == index ? _GEN_7705 : tag_1_1; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1036 = 7'h2 == index ? _GEN_7705 : tag_1_2; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1037 = 7'h3 == index ? _GEN_7705 : tag_1_3; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1038 = 7'h4 == index ? _GEN_7705 : tag_1_4; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1039 = 7'h5 == index ? _GEN_7705 : tag_1_5; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1040 = 7'h6 == index ? _GEN_7705 : tag_1_6; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1041 = 7'h7 == index ? _GEN_7705 : tag_1_7; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1042 = 7'h8 == index ? _GEN_7705 : tag_1_8; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1043 = 7'h9 == index ? _GEN_7705 : tag_1_9; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1044 = 7'ha == index ? _GEN_7705 : tag_1_10; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1045 = 7'hb == index ? _GEN_7705 : tag_1_11; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1046 = 7'hc == index ? _GEN_7705 : tag_1_12; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1047 = 7'hd == index ? _GEN_7705 : tag_1_13; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1048 = 7'he == index ? _GEN_7705 : tag_1_14; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1049 = 7'hf == index ? _GEN_7705 : tag_1_15; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1050 = 7'h10 == index ? _GEN_7705 : tag_1_16; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1051 = 7'h11 == index ? _GEN_7705 : tag_1_17; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1052 = 7'h12 == index ? _GEN_7705 : tag_1_18; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1053 = 7'h13 == index ? _GEN_7705 : tag_1_19; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1054 = 7'h14 == index ? _GEN_7705 : tag_1_20; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1055 = 7'h15 == index ? _GEN_7705 : tag_1_21; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1056 = 7'h16 == index ? _GEN_7705 : tag_1_22; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1057 = 7'h17 == index ? _GEN_7705 : tag_1_23; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1058 = 7'h18 == index ? _GEN_7705 : tag_1_24; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1059 = 7'h19 == index ? _GEN_7705 : tag_1_25; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1060 = 7'h1a == index ? _GEN_7705 : tag_1_26; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1061 = 7'h1b == index ? _GEN_7705 : tag_1_27; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1062 = 7'h1c == index ? _GEN_7705 : tag_1_28; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1063 = 7'h1d == index ? _GEN_7705 : tag_1_29; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1064 = 7'h1e == index ? _GEN_7705 : tag_1_30; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1065 = 7'h1f == index ? _GEN_7705 : tag_1_31; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1066 = 7'h20 == index ? _GEN_7705 : tag_1_32; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1067 = 7'h21 == index ? _GEN_7705 : tag_1_33; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1068 = 7'h22 == index ? _GEN_7705 : tag_1_34; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1069 = 7'h23 == index ? _GEN_7705 : tag_1_35; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1070 = 7'h24 == index ? _GEN_7705 : tag_1_36; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1071 = 7'h25 == index ? _GEN_7705 : tag_1_37; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1072 = 7'h26 == index ? _GEN_7705 : tag_1_38; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1073 = 7'h27 == index ? _GEN_7705 : tag_1_39; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1074 = 7'h28 == index ? _GEN_7705 : tag_1_40; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1075 = 7'h29 == index ? _GEN_7705 : tag_1_41; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1076 = 7'h2a == index ? _GEN_7705 : tag_1_42; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1077 = 7'h2b == index ? _GEN_7705 : tag_1_43; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1078 = 7'h2c == index ? _GEN_7705 : tag_1_44; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1079 = 7'h2d == index ? _GEN_7705 : tag_1_45; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1080 = 7'h2e == index ? _GEN_7705 : tag_1_46; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1081 = 7'h2f == index ? _GEN_7705 : tag_1_47; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1082 = 7'h30 == index ? _GEN_7705 : tag_1_48; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1083 = 7'h31 == index ? _GEN_7705 : tag_1_49; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1084 = 7'h32 == index ? _GEN_7705 : tag_1_50; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1085 = 7'h33 == index ? _GEN_7705 : tag_1_51; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1086 = 7'h34 == index ? _GEN_7705 : tag_1_52; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1087 = 7'h35 == index ? _GEN_7705 : tag_1_53; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1088 = 7'h36 == index ? _GEN_7705 : tag_1_54; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1089 = 7'h37 == index ? _GEN_7705 : tag_1_55; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1090 = 7'h38 == index ? _GEN_7705 : tag_1_56; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1091 = 7'h39 == index ? _GEN_7705 : tag_1_57; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1092 = 7'h3a == index ? _GEN_7705 : tag_1_58; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1093 = 7'h3b == index ? _GEN_7705 : tag_1_59; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1094 = 7'h3c == index ? _GEN_7705 : tag_1_60; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1095 = 7'h3d == index ? _GEN_7705 : tag_1_61; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1096 = 7'h3e == index ? _GEN_7705 : tag_1_62; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1097 = 7'h3f == index ? _GEN_7705 : tag_1_63; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1098 = 7'h40 == index ? _GEN_7705 : tag_1_64; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1099 = 7'h41 == index ? _GEN_7705 : tag_1_65; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1100 = 7'h42 == index ? _GEN_7705 : tag_1_66; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1101 = 7'h43 == index ? _GEN_7705 : tag_1_67; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1102 = 7'h44 == index ? _GEN_7705 : tag_1_68; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1103 = 7'h45 == index ? _GEN_7705 : tag_1_69; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1104 = 7'h46 == index ? _GEN_7705 : tag_1_70; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1105 = 7'h47 == index ? _GEN_7705 : tag_1_71; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1106 = 7'h48 == index ? _GEN_7705 : tag_1_72; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1107 = 7'h49 == index ? _GEN_7705 : tag_1_73; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1108 = 7'h4a == index ? _GEN_7705 : tag_1_74; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1109 = 7'h4b == index ? _GEN_7705 : tag_1_75; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1110 = 7'h4c == index ? _GEN_7705 : tag_1_76; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1111 = 7'h4d == index ? _GEN_7705 : tag_1_77; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1112 = 7'h4e == index ? _GEN_7705 : tag_1_78; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1113 = 7'h4f == index ? _GEN_7705 : tag_1_79; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1114 = 7'h50 == index ? _GEN_7705 : tag_1_80; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1115 = 7'h51 == index ? _GEN_7705 : tag_1_81; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1116 = 7'h52 == index ? _GEN_7705 : tag_1_82; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1117 = 7'h53 == index ? _GEN_7705 : tag_1_83; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1118 = 7'h54 == index ? _GEN_7705 : tag_1_84; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1119 = 7'h55 == index ? _GEN_7705 : tag_1_85; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1120 = 7'h56 == index ? _GEN_7705 : tag_1_86; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1121 = 7'h57 == index ? _GEN_7705 : tag_1_87; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1122 = 7'h58 == index ? _GEN_7705 : tag_1_88; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1123 = 7'h59 == index ? _GEN_7705 : tag_1_89; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1124 = 7'h5a == index ? _GEN_7705 : tag_1_90; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1125 = 7'h5b == index ? _GEN_7705 : tag_1_91; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1126 = 7'h5c == index ? _GEN_7705 : tag_1_92; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1127 = 7'h5d == index ? _GEN_7705 : tag_1_93; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1128 = 7'h5e == index ? _GEN_7705 : tag_1_94; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1129 = 7'h5f == index ? _GEN_7705 : tag_1_95; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1130 = 7'h60 == index ? _GEN_7705 : tag_1_96; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1131 = 7'h61 == index ? _GEN_7705 : tag_1_97; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1132 = 7'h62 == index ? _GEN_7705 : tag_1_98; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1133 = 7'h63 == index ? _GEN_7705 : tag_1_99; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1134 = 7'h64 == index ? _GEN_7705 : tag_1_100; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1135 = 7'h65 == index ? _GEN_7705 : tag_1_101; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1136 = 7'h66 == index ? _GEN_7705 : tag_1_102; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1137 = 7'h67 == index ? _GEN_7705 : tag_1_103; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1138 = 7'h68 == index ? _GEN_7705 : tag_1_104; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1139 = 7'h69 == index ? _GEN_7705 : tag_1_105; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1140 = 7'h6a == index ? _GEN_7705 : tag_1_106; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1141 = 7'h6b == index ? _GEN_7705 : tag_1_107; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1142 = 7'h6c == index ? _GEN_7705 : tag_1_108; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1143 = 7'h6d == index ? _GEN_7705 : tag_1_109; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1144 = 7'h6e == index ? _GEN_7705 : tag_1_110; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1145 = 7'h6f == index ? _GEN_7705 : tag_1_111; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1146 = 7'h70 == index ? _GEN_7705 : tag_1_112; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1147 = 7'h71 == index ? _GEN_7705 : tag_1_113; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1148 = 7'h72 == index ? _GEN_7705 : tag_1_114; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1149 = 7'h73 == index ? _GEN_7705 : tag_1_115; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1150 = 7'h74 == index ? _GEN_7705 : tag_1_116; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1151 = 7'h75 == index ? _GEN_7705 : tag_1_117; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1152 = 7'h76 == index ? _GEN_7705 : tag_1_118; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1153 = 7'h77 == index ? _GEN_7705 : tag_1_119; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1154 = 7'h78 == index ? _GEN_7705 : tag_1_120; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1155 = 7'h79 == index ? _GEN_7705 : tag_1_121; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1156 = 7'h7a == index ? _GEN_7705 : tag_1_122; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1157 = 7'h7b == index ? _GEN_7705 : tag_1_123; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1158 = 7'h7c == index ? _GEN_7705 : tag_1_124; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1159 = 7'h7d == index ? _GEN_7705 : tag_1_125; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1160 = 7'h7e == index ? _GEN_7705 : tag_1_126; // @[cache.scala 20:24 89:{30,30}]
  wire [31:0] _GEN_1161 = 7'h7f == index ? _GEN_7705 : tag_1_127; // @[cache.scala 20:24 89:{30,30}]
  wire  _GEN_1162 = _GEN_7709 | valid_1_0; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1163 = _GEN_7711 | valid_1_1; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1164 = _GEN_7713 | valid_1_2; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1165 = _GEN_7717 | valid_1_3; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1166 = _GEN_7726 | valid_1_4; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1167 = _GEN_7728 | valid_1_5; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1168 = _GEN_7730 | valid_1_6; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1169 = _GEN_7732 | valid_1_7; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1170 = _GEN_7737 | valid_1_8; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1171 = _GEN_7738 | valid_1_9; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1172 = _GEN_7739 | valid_1_10; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1173 = _GEN_7740 | valid_1_11; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1174 = _GEN_7741 | valid_1_12; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1175 = _GEN_7742 | valid_1_13; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1176 = _GEN_7743 | valid_1_14; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1177 = _GEN_7744 | valid_1_15; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1178 = _GEN_7745 | valid_1_16; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1179 = _GEN_7746 | valid_1_17; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1180 = _GEN_7747 | valid_1_18; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1181 = _GEN_7748 | valid_1_19; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1182 = _GEN_7749 | valid_1_20; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1183 = _GEN_7750 | valid_1_21; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1184 = _GEN_7751 | valid_1_22; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1185 = _GEN_7752 | valid_1_23; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1186 = _GEN_7753 | valid_1_24; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1187 = _GEN_7754 | valid_1_25; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1188 = _GEN_7755 | valid_1_26; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1189 = _GEN_7756 | valid_1_27; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1190 = _GEN_7757 | valid_1_28; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1191 = _GEN_7758 | valid_1_29; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1192 = _GEN_7759 | valid_1_30; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1193 = _GEN_7760 | valid_1_31; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1194 = _GEN_7761 | valid_1_32; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1195 = _GEN_7762 | valid_1_33; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1196 = _GEN_7763 | valid_1_34; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1197 = _GEN_7764 | valid_1_35; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1198 = _GEN_7765 | valid_1_36; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1199 = _GEN_7766 | valid_1_37; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1200 = _GEN_7767 | valid_1_38; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1201 = _GEN_7768 | valid_1_39; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1202 = _GEN_7769 | valid_1_40; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1203 = _GEN_7770 | valid_1_41; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1204 = _GEN_7771 | valid_1_42; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1205 = _GEN_7772 | valid_1_43; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1206 = _GEN_7773 | valid_1_44; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1207 = _GEN_7774 | valid_1_45; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1208 = _GEN_7775 | valid_1_46; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1209 = _GEN_7776 | valid_1_47; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1210 = _GEN_7777 | valid_1_48; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1211 = _GEN_7778 | valid_1_49; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1212 = _GEN_7779 | valid_1_50; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1213 = _GEN_7780 | valid_1_51; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1214 = _GEN_7781 | valid_1_52; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1215 = _GEN_7782 | valid_1_53; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1216 = _GEN_7783 | valid_1_54; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1217 = _GEN_7784 | valid_1_55; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1218 = _GEN_7785 | valid_1_56; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1219 = _GEN_7786 | valid_1_57; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1220 = _GEN_7787 | valid_1_58; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1221 = _GEN_7788 | valid_1_59; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1222 = _GEN_7789 | valid_1_60; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1223 = _GEN_7790 | valid_1_61; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1224 = _GEN_7791 | valid_1_62; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1225 = _GEN_7792 | valid_1_63; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1226 = _GEN_7793 | valid_1_64; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1227 = _GEN_7794 | valid_1_65; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1228 = _GEN_7795 | valid_1_66; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1229 = _GEN_7796 | valid_1_67; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1230 = _GEN_7797 | valid_1_68; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1231 = _GEN_7798 | valid_1_69; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1232 = _GEN_7799 | valid_1_70; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1233 = _GEN_7800 | valid_1_71; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1234 = _GEN_7801 | valid_1_72; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1235 = _GEN_7802 | valid_1_73; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1236 = _GEN_7803 | valid_1_74; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1237 = _GEN_7804 | valid_1_75; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1238 = _GEN_7805 | valid_1_76; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1239 = _GEN_7806 | valid_1_77; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1240 = _GEN_7807 | valid_1_78; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1241 = _GEN_7808 | valid_1_79; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1242 = _GEN_7809 | valid_1_80; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1243 = _GEN_7810 | valid_1_81; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1244 = _GEN_7811 | valid_1_82; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1245 = _GEN_7812 | valid_1_83; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1246 = _GEN_7813 | valid_1_84; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1247 = _GEN_7814 | valid_1_85; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1248 = _GEN_7815 | valid_1_86; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1249 = _GEN_7816 | valid_1_87; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1250 = _GEN_7817 | valid_1_88; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1251 = _GEN_7818 | valid_1_89; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1252 = _GEN_7819 | valid_1_90; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1253 = _GEN_7820 | valid_1_91; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1254 = _GEN_7821 | valid_1_92; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1255 = _GEN_7822 | valid_1_93; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1256 = _GEN_7823 | valid_1_94; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1257 = _GEN_7824 | valid_1_95; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1258 = _GEN_7825 | valid_1_96; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1259 = _GEN_7826 | valid_1_97; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1260 = _GEN_7827 | valid_1_98; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1261 = _GEN_7828 | valid_1_99; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1262 = _GEN_7829 | valid_1_100; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1263 = _GEN_7830 | valid_1_101; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1264 = _GEN_7831 | valid_1_102; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1265 = _GEN_7832 | valid_1_103; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1266 = _GEN_7833 | valid_1_104; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1267 = _GEN_7834 | valid_1_105; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1268 = _GEN_7835 | valid_1_106; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1269 = _GEN_7836 | valid_1_107; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1270 = _GEN_7837 | valid_1_108; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1271 = _GEN_7838 | valid_1_109; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1272 = _GEN_7839 | valid_1_110; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1273 = _GEN_7840 | valid_1_111; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1274 = _GEN_7841 | valid_1_112; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1275 = _GEN_7842 | valid_1_113; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1276 = _GEN_7843 | valid_1_114; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1277 = _GEN_7844 | valid_1_115; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1278 = _GEN_7845 | valid_1_116; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1279 = _GEN_7846 | valid_1_117; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1280 = _GEN_7847 | valid_1_118; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1281 = _GEN_7848 | valid_1_119; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1282 = _GEN_7849 | valid_1_120; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1283 = _GEN_7850 | valid_1_121; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1284 = _GEN_7851 | valid_1_122; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1285 = _GEN_7852 | valid_1_123; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1286 = _GEN_7853 | valid_1_124; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1287 = _GEN_7854 | valid_1_125; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1288 = _GEN_7855 | valid_1_126; // @[cache.scala 22:26 90:{32,32}]
  wire  _GEN_1289 = _GEN_7856 | valid_1_127; // @[cache.scala 22:26 90:{32,32}]
  wire  _T_18 = ~quene; // @[cache.scala 93:27]
  wire [63:0] _GEN_2058 = ~quene ? _GEN_522 : ram_0_0; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2059 = ~quene ? _GEN_523 : ram_0_1; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2060 = ~quene ? _GEN_524 : ram_0_2; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2061 = ~quene ? _GEN_525 : ram_0_3; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2062 = ~quene ? _GEN_526 : ram_0_4; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2063 = ~quene ? _GEN_527 : ram_0_5; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2064 = ~quene ? _GEN_528 : ram_0_6; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2065 = ~quene ? _GEN_529 : ram_0_7; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2066 = ~quene ? _GEN_530 : ram_0_8; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2067 = ~quene ? _GEN_531 : ram_0_9; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2068 = ~quene ? _GEN_532 : ram_0_10; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2069 = ~quene ? _GEN_533 : ram_0_11; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2070 = ~quene ? _GEN_534 : ram_0_12; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2071 = ~quene ? _GEN_535 : ram_0_13; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2072 = ~quene ? _GEN_536 : ram_0_14; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2073 = ~quene ? _GEN_537 : ram_0_15; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2074 = ~quene ? _GEN_538 : ram_0_16; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2075 = ~quene ? _GEN_539 : ram_0_17; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2076 = ~quene ? _GEN_540 : ram_0_18; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2077 = ~quene ? _GEN_541 : ram_0_19; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2078 = ~quene ? _GEN_542 : ram_0_20; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2079 = ~quene ? _GEN_543 : ram_0_21; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2080 = ~quene ? _GEN_544 : ram_0_22; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2081 = ~quene ? _GEN_545 : ram_0_23; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2082 = ~quene ? _GEN_546 : ram_0_24; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2083 = ~quene ? _GEN_547 : ram_0_25; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2084 = ~quene ? _GEN_548 : ram_0_26; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2085 = ~quene ? _GEN_549 : ram_0_27; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2086 = ~quene ? _GEN_550 : ram_0_28; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2087 = ~quene ? _GEN_551 : ram_0_29; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2088 = ~quene ? _GEN_552 : ram_0_30; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2089 = ~quene ? _GEN_553 : ram_0_31; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2090 = ~quene ? _GEN_554 : ram_0_32; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2091 = ~quene ? _GEN_555 : ram_0_33; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2092 = ~quene ? _GEN_556 : ram_0_34; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2093 = ~quene ? _GEN_557 : ram_0_35; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2094 = ~quene ? _GEN_558 : ram_0_36; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2095 = ~quene ? _GEN_559 : ram_0_37; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2096 = ~quene ? _GEN_560 : ram_0_38; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2097 = ~quene ? _GEN_561 : ram_0_39; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2098 = ~quene ? _GEN_562 : ram_0_40; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2099 = ~quene ? _GEN_563 : ram_0_41; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2100 = ~quene ? _GEN_564 : ram_0_42; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2101 = ~quene ? _GEN_565 : ram_0_43; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2102 = ~quene ? _GEN_566 : ram_0_44; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2103 = ~quene ? _GEN_567 : ram_0_45; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2104 = ~quene ? _GEN_568 : ram_0_46; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2105 = ~quene ? _GEN_569 : ram_0_47; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2106 = ~quene ? _GEN_570 : ram_0_48; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2107 = ~quene ? _GEN_571 : ram_0_49; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2108 = ~quene ? _GEN_572 : ram_0_50; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2109 = ~quene ? _GEN_573 : ram_0_51; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2110 = ~quene ? _GEN_574 : ram_0_52; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2111 = ~quene ? _GEN_575 : ram_0_53; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2112 = ~quene ? _GEN_576 : ram_0_54; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2113 = ~quene ? _GEN_577 : ram_0_55; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2114 = ~quene ? _GEN_578 : ram_0_56; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2115 = ~quene ? _GEN_579 : ram_0_57; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2116 = ~quene ? _GEN_580 : ram_0_58; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2117 = ~quene ? _GEN_581 : ram_0_59; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2118 = ~quene ? _GEN_582 : ram_0_60; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2119 = ~quene ? _GEN_583 : ram_0_61; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2120 = ~quene ? _GEN_584 : ram_0_62; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2121 = ~quene ? _GEN_585 : ram_0_63; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2122 = ~quene ? _GEN_586 : ram_0_64; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2123 = ~quene ? _GEN_587 : ram_0_65; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2124 = ~quene ? _GEN_588 : ram_0_66; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2125 = ~quene ? _GEN_589 : ram_0_67; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2126 = ~quene ? _GEN_590 : ram_0_68; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2127 = ~quene ? _GEN_591 : ram_0_69; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2128 = ~quene ? _GEN_592 : ram_0_70; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2129 = ~quene ? _GEN_593 : ram_0_71; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2130 = ~quene ? _GEN_594 : ram_0_72; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2131 = ~quene ? _GEN_595 : ram_0_73; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2132 = ~quene ? _GEN_596 : ram_0_74; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2133 = ~quene ? _GEN_597 : ram_0_75; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2134 = ~quene ? _GEN_598 : ram_0_76; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2135 = ~quene ? _GEN_599 : ram_0_77; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2136 = ~quene ? _GEN_600 : ram_0_78; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2137 = ~quene ? _GEN_601 : ram_0_79; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2138 = ~quene ? _GEN_602 : ram_0_80; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2139 = ~quene ? _GEN_603 : ram_0_81; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2140 = ~quene ? _GEN_604 : ram_0_82; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2141 = ~quene ? _GEN_605 : ram_0_83; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2142 = ~quene ? _GEN_606 : ram_0_84; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2143 = ~quene ? _GEN_607 : ram_0_85; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2144 = ~quene ? _GEN_608 : ram_0_86; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2145 = ~quene ? _GEN_609 : ram_0_87; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2146 = ~quene ? _GEN_610 : ram_0_88; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2147 = ~quene ? _GEN_611 : ram_0_89; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2148 = ~quene ? _GEN_612 : ram_0_90; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2149 = ~quene ? _GEN_613 : ram_0_91; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2150 = ~quene ? _GEN_614 : ram_0_92; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2151 = ~quene ? _GEN_615 : ram_0_93; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2152 = ~quene ? _GEN_616 : ram_0_94; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2153 = ~quene ? _GEN_617 : ram_0_95; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2154 = ~quene ? _GEN_618 : ram_0_96; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2155 = ~quene ? _GEN_619 : ram_0_97; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2156 = ~quene ? _GEN_620 : ram_0_98; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2157 = ~quene ? _GEN_621 : ram_0_99; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2158 = ~quene ? _GEN_622 : ram_0_100; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2159 = ~quene ? _GEN_623 : ram_0_101; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2160 = ~quene ? _GEN_624 : ram_0_102; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2161 = ~quene ? _GEN_625 : ram_0_103; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2162 = ~quene ? _GEN_626 : ram_0_104; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2163 = ~quene ? _GEN_627 : ram_0_105; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2164 = ~quene ? _GEN_628 : ram_0_106; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2165 = ~quene ? _GEN_629 : ram_0_107; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2166 = ~quene ? _GEN_630 : ram_0_108; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2167 = ~quene ? _GEN_631 : ram_0_109; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2168 = ~quene ? _GEN_632 : ram_0_110; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2169 = ~quene ? _GEN_633 : ram_0_111; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2170 = ~quene ? _GEN_634 : ram_0_112; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2171 = ~quene ? _GEN_635 : ram_0_113; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2172 = ~quene ? _GEN_636 : ram_0_114; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2173 = ~quene ? _GEN_637 : ram_0_115; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2174 = ~quene ? _GEN_638 : ram_0_116; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2175 = ~quene ? _GEN_639 : ram_0_117; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2176 = ~quene ? _GEN_640 : ram_0_118; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2177 = ~quene ? _GEN_641 : ram_0_119; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2178 = ~quene ? _GEN_642 : ram_0_120; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2179 = ~quene ? _GEN_643 : ram_0_121; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2180 = ~quene ? _GEN_644 : ram_0_122; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2181 = ~quene ? _GEN_645 : ram_0_123; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2182 = ~quene ? _GEN_646 : ram_0_124; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2183 = ~quene ? _GEN_647 : ram_0_125; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2184 = ~quene ? _GEN_648 : ram_0_126; // @[cache.scala 17:24 93:34]
  wire [63:0] _GEN_2185 = ~quene ? _GEN_649 : ram_0_127; // @[cache.scala 17:24 93:34]
  wire [31:0] _GEN_2186 = ~quene ? _GEN_650 : tag_0_0; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2187 = ~quene ? _GEN_651 : tag_0_1; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2188 = ~quene ? _GEN_652 : tag_0_2; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2189 = ~quene ? _GEN_653 : tag_0_3; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2190 = ~quene ? _GEN_654 : tag_0_4; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2191 = ~quene ? _GEN_655 : tag_0_5; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2192 = ~quene ? _GEN_656 : tag_0_6; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2193 = ~quene ? _GEN_657 : tag_0_7; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2194 = ~quene ? _GEN_658 : tag_0_8; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2195 = ~quene ? _GEN_659 : tag_0_9; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2196 = ~quene ? _GEN_660 : tag_0_10; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2197 = ~quene ? _GEN_661 : tag_0_11; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2198 = ~quene ? _GEN_662 : tag_0_12; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2199 = ~quene ? _GEN_663 : tag_0_13; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2200 = ~quene ? _GEN_664 : tag_0_14; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2201 = ~quene ? _GEN_665 : tag_0_15; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2202 = ~quene ? _GEN_666 : tag_0_16; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2203 = ~quene ? _GEN_667 : tag_0_17; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2204 = ~quene ? _GEN_668 : tag_0_18; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2205 = ~quene ? _GEN_669 : tag_0_19; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2206 = ~quene ? _GEN_670 : tag_0_20; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2207 = ~quene ? _GEN_671 : tag_0_21; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2208 = ~quene ? _GEN_672 : tag_0_22; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2209 = ~quene ? _GEN_673 : tag_0_23; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2210 = ~quene ? _GEN_674 : tag_0_24; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2211 = ~quene ? _GEN_675 : tag_0_25; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2212 = ~quene ? _GEN_676 : tag_0_26; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2213 = ~quene ? _GEN_677 : tag_0_27; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2214 = ~quene ? _GEN_678 : tag_0_28; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2215 = ~quene ? _GEN_679 : tag_0_29; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2216 = ~quene ? _GEN_680 : tag_0_30; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2217 = ~quene ? _GEN_681 : tag_0_31; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2218 = ~quene ? _GEN_682 : tag_0_32; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2219 = ~quene ? _GEN_683 : tag_0_33; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2220 = ~quene ? _GEN_684 : tag_0_34; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2221 = ~quene ? _GEN_685 : tag_0_35; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2222 = ~quene ? _GEN_686 : tag_0_36; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2223 = ~quene ? _GEN_687 : tag_0_37; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2224 = ~quene ? _GEN_688 : tag_0_38; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2225 = ~quene ? _GEN_689 : tag_0_39; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2226 = ~quene ? _GEN_690 : tag_0_40; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2227 = ~quene ? _GEN_691 : tag_0_41; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2228 = ~quene ? _GEN_692 : tag_0_42; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2229 = ~quene ? _GEN_693 : tag_0_43; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2230 = ~quene ? _GEN_694 : tag_0_44; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2231 = ~quene ? _GEN_695 : tag_0_45; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2232 = ~quene ? _GEN_696 : tag_0_46; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2233 = ~quene ? _GEN_697 : tag_0_47; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2234 = ~quene ? _GEN_698 : tag_0_48; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2235 = ~quene ? _GEN_699 : tag_0_49; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2236 = ~quene ? _GEN_700 : tag_0_50; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2237 = ~quene ? _GEN_701 : tag_0_51; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2238 = ~quene ? _GEN_702 : tag_0_52; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2239 = ~quene ? _GEN_703 : tag_0_53; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2240 = ~quene ? _GEN_704 : tag_0_54; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2241 = ~quene ? _GEN_705 : tag_0_55; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2242 = ~quene ? _GEN_706 : tag_0_56; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2243 = ~quene ? _GEN_707 : tag_0_57; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2244 = ~quene ? _GEN_708 : tag_0_58; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2245 = ~quene ? _GEN_709 : tag_0_59; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2246 = ~quene ? _GEN_710 : tag_0_60; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2247 = ~quene ? _GEN_711 : tag_0_61; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2248 = ~quene ? _GEN_712 : tag_0_62; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2249 = ~quene ? _GEN_713 : tag_0_63; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2250 = ~quene ? _GEN_714 : tag_0_64; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2251 = ~quene ? _GEN_715 : tag_0_65; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2252 = ~quene ? _GEN_716 : tag_0_66; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2253 = ~quene ? _GEN_717 : tag_0_67; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2254 = ~quene ? _GEN_718 : tag_0_68; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2255 = ~quene ? _GEN_719 : tag_0_69; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2256 = ~quene ? _GEN_720 : tag_0_70; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2257 = ~quene ? _GEN_721 : tag_0_71; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2258 = ~quene ? _GEN_722 : tag_0_72; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2259 = ~quene ? _GEN_723 : tag_0_73; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2260 = ~quene ? _GEN_724 : tag_0_74; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2261 = ~quene ? _GEN_725 : tag_0_75; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2262 = ~quene ? _GEN_726 : tag_0_76; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2263 = ~quene ? _GEN_727 : tag_0_77; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2264 = ~quene ? _GEN_728 : tag_0_78; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2265 = ~quene ? _GEN_729 : tag_0_79; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2266 = ~quene ? _GEN_730 : tag_0_80; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2267 = ~quene ? _GEN_731 : tag_0_81; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2268 = ~quene ? _GEN_732 : tag_0_82; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2269 = ~quene ? _GEN_733 : tag_0_83; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2270 = ~quene ? _GEN_734 : tag_0_84; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2271 = ~quene ? _GEN_735 : tag_0_85; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2272 = ~quene ? _GEN_736 : tag_0_86; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2273 = ~quene ? _GEN_737 : tag_0_87; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2274 = ~quene ? _GEN_738 : tag_0_88; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2275 = ~quene ? _GEN_739 : tag_0_89; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2276 = ~quene ? _GEN_740 : tag_0_90; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2277 = ~quene ? _GEN_741 : tag_0_91; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2278 = ~quene ? _GEN_742 : tag_0_92; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2279 = ~quene ? _GEN_743 : tag_0_93; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2280 = ~quene ? _GEN_744 : tag_0_94; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2281 = ~quene ? _GEN_745 : tag_0_95; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2282 = ~quene ? _GEN_746 : tag_0_96; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2283 = ~quene ? _GEN_747 : tag_0_97; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2284 = ~quene ? _GEN_748 : tag_0_98; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2285 = ~quene ? _GEN_749 : tag_0_99; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2286 = ~quene ? _GEN_750 : tag_0_100; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2287 = ~quene ? _GEN_751 : tag_0_101; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2288 = ~quene ? _GEN_752 : tag_0_102; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2289 = ~quene ? _GEN_753 : tag_0_103; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2290 = ~quene ? _GEN_754 : tag_0_104; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2291 = ~quene ? _GEN_755 : tag_0_105; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2292 = ~quene ? _GEN_756 : tag_0_106; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2293 = ~quene ? _GEN_757 : tag_0_107; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2294 = ~quene ? _GEN_758 : tag_0_108; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2295 = ~quene ? _GEN_759 : tag_0_109; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2296 = ~quene ? _GEN_760 : tag_0_110; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2297 = ~quene ? _GEN_761 : tag_0_111; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2298 = ~quene ? _GEN_762 : tag_0_112; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2299 = ~quene ? _GEN_763 : tag_0_113; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2300 = ~quene ? _GEN_764 : tag_0_114; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2301 = ~quene ? _GEN_765 : tag_0_115; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2302 = ~quene ? _GEN_766 : tag_0_116; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2303 = ~quene ? _GEN_767 : tag_0_117; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2304 = ~quene ? _GEN_768 : tag_0_118; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2305 = ~quene ? _GEN_769 : tag_0_119; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2306 = ~quene ? _GEN_770 : tag_0_120; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2307 = ~quene ? _GEN_771 : tag_0_121; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2308 = ~quene ? _GEN_772 : tag_0_122; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2309 = ~quene ? _GEN_773 : tag_0_123; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2310 = ~quene ? _GEN_774 : tag_0_124; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2311 = ~quene ? _GEN_775 : tag_0_125; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2312 = ~quene ? _GEN_776 : tag_0_126; // @[cache.scala 19:24 93:34]
  wire [31:0] _GEN_2313 = ~quene ? _GEN_777 : tag_0_127; // @[cache.scala 19:24 93:34]
  wire  _GEN_2314 = ~quene ? _GEN_778 : valid_0_0; // @[cache.scala 21:26 93:34]
  wire  _GEN_2315 = ~quene ? _GEN_779 : valid_0_1; // @[cache.scala 21:26 93:34]
  wire  _GEN_2316 = ~quene ? _GEN_780 : valid_0_2; // @[cache.scala 21:26 93:34]
  wire  _GEN_2317 = ~quene ? _GEN_781 : valid_0_3; // @[cache.scala 21:26 93:34]
  wire  _GEN_2318 = ~quene ? _GEN_782 : valid_0_4; // @[cache.scala 21:26 93:34]
  wire  _GEN_2319 = ~quene ? _GEN_783 : valid_0_5; // @[cache.scala 21:26 93:34]
  wire  _GEN_2320 = ~quene ? _GEN_784 : valid_0_6; // @[cache.scala 21:26 93:34]
  wire  _GEN_2321 = ~quene ? _GEN_785 : valid_0_7; // @[cache.scala 21:26 93:34]
  wire  _GEN_2322 = ~quene ? _GEN_786 : valid_0_8; // @[cache.scala 21:26 93:34]
  wire  _GEN_2323 = ~quene ? _GEN_787 : valid_0_9; // @[cache.scala 21:26 93:34]
  wire  _GEN_2324 = ~quene ? _GEN_788 : valid_0_10; // @[cache.scala 21:26 93:34]
  wire  _GEN_2325 = ~quene ? _GEN_789 : valid_0_11; // @[cache.scala 21:26 93:34]
  wire  _GEN_2326 = ~quene ? _GEN_790 : valid_0_12; // @[cache.scala 21:26 93:34]
  wire  _GEN_2327 = ~quene ? _GEN_791 : valid_0_13; // @[cache.scala 21:26 93:34]
  wire  _GEN_2328 = ~quene ? _GEN_792 : valid_0_14; // @[cache.scala 21:26 93:34]
  wire  _GEN_2329 = ~quene ? _GEN_793 : valid_0_15; // @[cache.scala 21:26 93:34]
  wire  _GEN_2330 = ~quene ? _GEN_794 : valid_0_16; // @[cache.scala 21:26 93:34]
  wire  _GEN_2331 = ~quene ? _GEN_795 : valid_0_17; // @[cache.scala 21:26 93:34]
  wire  _GEN_2332 = ~quene ? _GEN_796 : valid_0_18; // @[cache.scala 21:26 93:34]
  wire  _GEN_2333 = ~quene ? _GEN_797 : valid_0_19; // @[cache.scala 21:26 93:34]
  wire  _GEN_2334 = ~quene ? _GEN_798 : valid_0_20; // @[cache.scala 21:26 93:34]
  wire  _GEN_2335 = ~quene ? _GEN_799 : valid_0_21; // @[cache.scala 21:26 93:34]
  wire  _GEN_2336 = ~quene ? _GEN_800 : valid_0_22; // @[cache.scala 21:26 93:34]
  wire  _GEN_2337 = ~quene ? _GEN_801 : valid_0_23; // @[cache.scala 21:26 93:34]
  wire  _GEN_2338 = ~quene ? _GEN_802 : valid_0_24; // @[cache.scala 21:26 93:34]
  wire  _GEN_2339 = ~quene ? _GEN_803 : valid_0_25; // @[cache.scala 21:26 93:34]
  wire  _GEN_2340 = ~quene ? _GEN_804 : valid_0_26; // @[cache.scala 21:26 93:34]
  wire  _GEN_2341 = ~quene ? _GEN_805 : valid_0_27; // @[cache.scala 21:26 93:34]
  wire  _GEN_2342 = ~quene ? _GEN_806 : valid_0_28; // @[cache.scala 21:26 93:34]
  wire  _GEN_2343 = ~quene ? _GEN_807 : valid_0_29; // @[cache.scala 21:26 93:34]
  wire  _GEN_2344 = ~quene ? _GEN_808 : valid_0_30; // @[cache.scala 21:26 93:34]
  wire  _GEN_2345 = ~quene ? _GEN_809 : valid_0_31; // @[cache.scala 21:26 93:34]
  wire  _GEN_2346 = ~quene ? _GEN_810 : valid_0_32; // @[cache.scala 21:26 93:34]
  wire  _GEN_2347 = ~quene ? _GEN_811 : valid_0_33; // @[cache.scala 21:26 93:34]
  wire  _GEN_2348 = ~quene ? _GEN_812 : valid_0_34; // @[cache.scala 21:26 93:34]
  wire  _GEN_2349 = ~quene ? _GEN_813 : valid_0_35; // @[cache.scala 21:26 93:34]
  wire  _GEN_2350 = ~quene ? _GEN_814 : valid_0_36; // @[cache.scala 21:26 93:34]
  wire  _GEN_2351 = ~quene ? _GEN_815 : valid_0_37; // @[cache.scala 21:26 93:34]
  wire  _GEN_2352 = ~quene ? _GEN_816 : valid_0_38; // @[cache.scala 21:26 93:34]
  wire  _GEN_2353 = ~quene ? _GEN_817 : valid_0_39; // @[cache.scala 21:26 93:34]
  wire  _GEN_2354 = ~quene ? _GEN_818 : valid_0_40; // @[cache.scala 21:26 93:34]
  wire  _GEN_2355 = ~quene ? _GEN_819 : valid_0_41; // @[cache.scala 21:26 93:34]
  wire  _GEN_2356 = ~quene ? _GEN_820 : valid_0_42; // @[cache.scala 21:26 93:34]
  wire  _GEN_2357 = ~quene ? _GEN_821 : valid_0_43; // @[cache.scala 21:26 93:34]
  wire  _GEN_2358 = ~quene ? _GEN_822 : valid_0_44; // @[cache.scala 21:26 93:34]
  wire  _GEN_2359 = ~quene ? _GEN_823 : valid_0_45; // @[cache.scala 21:26 93:34]
  wire  _GEN_2360 = ~quene ? _GEN_824 : valid_0_46; // @[cache.scala 21:26 93:34]
  wire  _GEN_2361 = ~quene ? _GEN_825 : valid_0_47; // @[cache.scala 21:26 93:34]
  wire  _GEN_2362 = ~quene ? _GEN_826 : valid_0_48; // @[cache.scala 21:26 93:34]
  wire  _GEN_2363 = ~quene ? _GEN_827 : valid_0_49; // @[cache.scala 21:26 93:34]
  wire  _GEN_2364 = ~quene ? _GEN_828 : valid_0_50; // @[cache.scala 21:26 93:34]
  wire  _GEN_2365 = ~quene ? _GEN_829 : valid_0_51; // @[cache.scala 21:26 93:34]
  wire  _GEN_2366 = ~quene ? _GEN_830 : valid_0_52; // @[cache.scala 21:26 93:34]
  wire  _GEN_2367 = ~quene ? _GEN_831 : valid_0_53; // @[cache.scala 21:26 93:34]
  wire  _GEN_2368 = ~quene ? _GEN_832 : valid_0_54; // @[cache.scala 21:26 93:34]
  wire  _GEN_2369 = ~quene ? _GEN_833 : valid_0_55; // @[cache.scala 21:26 93:34]
  wire  _GEN_2370 = ~quene ? _GEN_834 : valid_0_56; // @[cache.scala 21:26 93:34]
  wire  _GEN_2371 = ~quene ? _GEN_835 : valid_0_57; // @[cache.scala 21:26 93:34]
  wire  _GEN_2372 = ~quene ? _GEN_836 : valid_0_58; // @[cache.scala 21:26 93:34]
  wire  _GEN_2373 = ~quene ? _GEN_837 : valid_0_59; // @[cache.scala 21:26 93:34]
  wire  _GEN_2374 = ~quene ? _GEN_838 : valid_0_60; // @[cache.scala 21:26 93:34]
  wire  _GEN_2375 = ~quene ? _GEN_839 : valid_0_61; // @[cache.scala 21:26 93:34]
  wire  _GEN_2376 = ~quene ? _GEN_840 : valid_0_62; // @[cache.scala 21:26 93:34]
  wire  _GEN_2377 = ~quene ? _GEN_841 : valid_0_63; // @[cache.scala 21:26 93:34]
  wire  _GEN_2378 = ~quene ? _GEN_842 : valid_0_64; // @[cache.scala 21:26 93:34]
  wire  _GEN_2379 = ~quene ? _GEN_843 : valid_0_65; // @[cache.scala 21:26 93:34]
  wire  _GEN_2380 = ~quene ? _GEN_844 : valid_0_66; // @[cache.scala 21:26 93:34]
  wire  _GEN_2381 = ~quene ? _GEN_845 : valid_0_67; // @[cache.scala 21:26 93:34]
  wire  _GEN_2382 = ~quene ? _GEN_846 : valid_0_68; // @[cache.scala 21:26 93:34]
  wire  _GEN_2383 = ~quene ? _GEN_847 : valid_0_69; // @[cache.scala 21:26 93:34]
  wire  _GEN_2384 = ~quene ? _GEN_848 : valid_0_70; // @[cache.scala 21:26 93:34]
  wire  _GEN_2385 = ~quene ? _GEN_849 : valid_0_71; // @[cache.scala 21:26 93:34]
  wire  _GEN_2386 = ~quene ? _GEN_850 : valid_0_72; // @[cache.scala 21:26 93:34]
  wire  _GEN_2387 = ~quene ? _GEN_851 : valid_0_73; // @[cache.scala 21:26 93:34]
  wire  _GEN_2388 = ~quene ? _GEN_852 : valid_0_74; // @[cache.scala 21:26 93:34]
  wire  _GEN_2389 = ~quene ? _GEN_853 : valid_0_75; // @[cache.scala 21:26 93:34]
  wire  _GEN_2390 = ~quene ? _GEN_854 : valid_0_76; // @[cache.scala 21:26 93:34]
  wire  _GEN_2391 = ~quene ? _GEN_855 : valid_0_77; // @[cache.scala 21:26 93:34]
  wire  _GEN_2392 = ~quene ? _GEN_856 : valid_0_78; // @[cache.scala 21:26 93:34]
  wire  _GEN_2393 = ~quene ? _GEN_857 : valid_0_79; // @[cache.scala 21:26 93:34]
  wire  _GEN_2394 = ~quene ? _GEN_858 : valid_0_80; // @[cache.scala 21:26 93:34]
  wire  _GEN_2395 = ~quene ? _GEN_859 : valid_0_81; // @[cache.scala 21:26 93:34]
  wire  _GEN_2396 = ~quene ? _GEN_860 : valid_0_82; // @[cache.scala 21:26 93:34]
  wire  _GEN_2397 = ~quene ? _GEN_861 : valid_0_83; // @[cache.scala 21:26 93:34]
  wire  _GEN_2398 = ~quene ? _GEN_862 : valid_0_84; // @[cache.scala 21:26 93:34]
  wire  _GEN_2399 = ~quene ? _GEN_863 : valid_0_85; // @[cache.scala 21:26 93:34]
  wire  _GEN_2400 = ~quene ? _GEN_864 : valid_0_86; // @[cache.scala 21:26 93:34]
  wire  _GEN_2401 = ~quene ? _GEN_865 : valid_0_87; // @[cache.scala 21:26 93:34]
  wire  _GEN_2402 = ~quene ? _GEN_866 : valid_0_88; // @[cache.scala 21:26 93:34]
  wire  _GEN_2403 = ~quene ? _GEN_867 : valid_0_89; // @[cache.scala 21:26 93:34]
  wire  _GEN_2404 = ~quene ? _GEN_868 : valid_0_90; // @[cache.scala 21:26 93:34]
  wire  _GEN_2405 = ~quene ? _GEN_869 : valid_0_91; // @[cache.scala 21:26 93:34]
  wire  _GEN_2406 = ~quene ? _GEN_870 : valid_0_92; // @[cache.scala 21:26 93:34]
  wire  _GEN_2407 = ~quene ? _GEN_871 : valid_0_93; // @[cache.scala 21:26 93:34]
  wire  _GEN_2408 = ~quene ? _GEN_872 : valid_0_94; // @[cache.scala 21:26 93:34]
  wire  _GEN_2409 = ~quene ? _GEN_873 : valid_0_95; // @[cache.scala 21:26 93:34]
  wire  _GEN_2410 = ~quene ? _GEN_874 : valid_0_96; // @[cache.scala 21:26 93:34]
  wire  _GEN_2411 = ~quene ? _GEN_875 : valid_0_97; // @[cache.scala 21:26 93:34]
  wire  _GEN_2412 = ~quene ? _GEN_876 : valid_0_98; // @[cache.scala 21:26 93:34]
  wire  _GEN_2413 = ~quene ? _GEN_877 : valid_0_99; // @[cache.scala 21:26 93:34]
  wire  _GEN_2414 = ~quene ? _GEN_878 : valid_0_100; // @[cache.scala 21:26 93:34]
  wire  _GEN_2415 = ~quene ? _GEN_879 : valid_0_101; // @[cache.scala 21:26 93:34]
  wire  _GEN_2416 = ~quene ? _GEN_880 : valid_0_102; // @[cache.scala 21:26 93:34]
  wire  _GEN_2417 = ~quene ? _GEN_881 : valid_0_103; // @[cache.scala 21:26 93:34]
  wire  _GEN_2418 = ~quene ? _GEN_882 : valid_0_104; // @[cache.scala 21:26 93:34]
  wire  _GEN_2419 = ~quene ? _GEN_883 : valid_0_105; // @[cache.scala 21:26 93:34]
  wire  _GEN_2420 = ~quene ? _GEN_884 : valid_0_106; // @[cache.scala 21:26 93:34]
  wire  _GEN_2421 = ~quene ? _GEN_885 : valid_0_107; // @[cache.scala 21:26 93:34]
  wire  _GEN_2422 = ~quene ? _GEN_886 : valid_0_108; // @[cache.scala 21:26 93:34]
  wire  _GEN_2423 = ~quene ? _GEN_887 : valid_0_109; // @[cache.scala 21:26 93:34]
  wire  _GEN_2424 = ~quene ? _GEN_888 : valid_0_110; // @[cache.scala 21:26 93:34]
  wire  _GEN_2425 = ~quene ? _GEN_889 : valid_0_111; // @[cache.scala 21:26 93:34]
  wire  _GEN_2426 = ~quene ? _GEN_890 : valid_0_112; // @[cache.scala 21:26 93:34]
  wire  _GEN_2427 = ~quene ? _GEN_891 : valid_0_113; // @[cache.scala 21:26 93:34]
  wire  _GEN_2428 = ~quene ? _GEN_892 : valid_0_114; // @[cache.scala 21:26 93:34]
  wire  _GEN_2429 = ~quene ? _GEN_893 : valid_0_115; // @[cache.scala 21:26 93:34]
  wire  _GEN_2430 = ~quene ? _GEN_894 : valid_0_116; // @[cache.scala 21:26 93:34]
  wire  _GEN_2431 = ~quene ? _GEN_895 : valid_0_117; // @[cache.scala 21:26 93:34]
  wire  _GEN_2432 = ~quene ? _GEN_896 : valid_0_118; // @[cache.scala 21:26 93:34]
  wire  _GEN_2433 = ~quene ? _GEN_897 : valid_0_119; // @[cache.scala 21:26 93:34]
  wire  _GEN_2434 = ~quene ? _GEN_898 : valid_0_120; // @[cache.scala 21:26 93:34]
  wire  _GEN_2435 = ~quene ? _GEN_899 : valid_0_121; // @[cache.scala 21:26 93:34]
  wire  _GEN_2436 = ~quene ? _GEN_900 : valid_0_122; // @[cache.scala 21:26 93:34]
  wire  _GEN_2437 = ~quene ? _GEN_901 : valid_0_123; // @[cache.scala 21:26 93:34]
  wire  _GEN_2438 = ~quene ? _GEN_902 : valid_0_124; // @[cache.scala 21:26 93:34]
  wire  _GEN_2439 = ~quene ? _GEN_903 : valid_0_125; // @[cache.scala 21:26 93:34]
  wire  _GEN_2440 = ~quene ? _GEN_904 : valid_0_126; // @[cache.scala 21:26 93:34]
  wire  _GEN_2441 = ~quene ? _GEN_905 : valid_0_127; // @[cache.scala 21:26 93:34]
  wire [63:0] _GEN_2443 = ~quene ? ram_1_0 : _GEN_906; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2444 = ~quene ? ram_1_1 : _GEN_907; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2445 = ~quene ? ram_1_2 : _GEN_908; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2446 = ~quene ? ram_1_3 : _GEN_909; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2447 = ~quene ? ram_1_4 : _GEN_910; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2448 = ~quene ? ram_1_5 : _GEN_911; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2449 = ~quene ? ram_1_6 : _GEN_912; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2450 = ~quene ? ram_1_7 : _GEN_913; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2451 = ~quene ? ram_1_8 : _GEN_914; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2452 = ~quene ? ram_1_9 : _GEN_915; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2453 = ~quene ? ram_1_10 : _GEN_916; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2454 = ~quene ? ram_1_11 : _GEN_917; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2455 = ~quene ? ram_1_12 : _GEN_918; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2456 = ~quene ? ram_1_13 : _GEN_919; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2457 = ~quene ? ram_1_14 : _GEN_920; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2458 = ~quene ? ram_1_15 : _GEN_921; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2459 = ~quene ? ram_1_16 : _GEN_922; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2460 = ~quene ? ram_1_17 : _GEN_923; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2461 = ~quene ? ram_1_18 : _GEN_924; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2462 = ~quene ? ram_1_19 : _GEN_925; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2463 = ~quene ? ram_1_20 : _GEN_926; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2464 = ~quene ? ram_1_21 : _GEN_927; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2465 = ~quene ? ram_1_22 : _GEN_928; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2466 = ~quene ? ram_1_23 : _GEN_929; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2467 = ~quene ? ram_1_24 : _GEN_930; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2468 = ~quene ? ram_1_25 : _GEN_931; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2469 = ~quene ? ram_1_26 : _GEN_932; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2470 = ~quene ? ram_1_27 : _GEN_933; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2471 = ~quene ? ram_1_28 : _GEN_934; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2472 = ~quene ? ram_1_29 : _GEN_935; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2473 = ~quene ? ram_1_30 : _GEN_936; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2474 = ~quene ? ram_1_31 : _GEN_937; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2475 = ~quene ? ram_1_32 : _GEN_938; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2476 = ~quene ? ram_1_33 : _GEN_939; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2477 = ~quene ? ram_1_34 : _GEN_940; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2478 = ~quene ? ram_1_35 : _GEN_941; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2479 = ~quene ? ram_1_36 : _GEN_942; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2480 = ~quene ? ram_1_37 : _GEN_943; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2481 = ~quene ? ram_1_38 : _GEN_944; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2482 = ~quene ? ram_1_39 : _GEN_945; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2483 = ~quene ? ram_1_40 : _GEN_946; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2484 = ~quene ? ram_1_41 : _GEN_947; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2485 = ~quene ? ram_1_42 : _GEN_948; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2486 = ~quene ? ram_1_43 : _GEN_949; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2487 = ~quene ? ram_1_44 : _GEN_950; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2488 = ~quene ? ram_1_45 : _GEN_951; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2489 = ~quene ? ram_1_46 : _GEN_952; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2490 = ~quene ? ram_1_47 : _GEN_953; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2491 = ~quene ? ram_1_48 : _GEN_954; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2492 = ~quene ? ram_1_49 : _GEN_955; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2493 = ~quene ? ram_1_50 : _GEN_956; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2494 = ~quene ? ram_1_51 : _GEN_957; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2495 = ~quene ? ram_1_52 : _GEN_958; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2496 = ~quene ? ram_1_53 : _GEN_959; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2497 = ~quene ? ram_1_54 : _GEN_960; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2498 = ~quene ? ram_1_55 : _GEN_961; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2499 = ~quene ? ram_1_56 : _GEN_962; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2500 = ~quene ? ram_1_57 : _GEN_963; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2501 = ~quene ? ram_1_58 : _GEN_964; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2502 = ~quene ? ram_1_59 : _GEN_965; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2503 = ~quene ? ram_1_60 : _GEN_966; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2504 = ~quene ? ram_1_61 : _GEN_967; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2505 = ~quene ? ram_1_62 : _GEN_968; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2506 = ~quene ? ram_1_63 : _GEN_969; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2507 = ~quene ? ram_1_64 : _GEN_970; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2508 = ~quene ? ram_1_65 : _GEN_971; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2509 = ~quene ? ram_1_66 : _GEN_972; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2510 = ~quene ? ram_1_67 : _GEN_973; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2511 = ~quene ? ram_1_68 : _GEN_974; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2512 = ~quene ? ram_1_69 : _GEN_975; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2513 = ~quene ? ram_1_70 : _GEN_976; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2514 = ~quene ? ram_1_71 : _GEN_977; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2515 = ~quene ? ram_1_72 : _GEN_978; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2516 = ~quene ? ram_1_73 : _GEN_979; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2517 = ~quene ? ram_1_74 : _GEN_980; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2518 = ~quene ? ram_1_75 : _GEN_981; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2519 = ~quene ? ram_1_76 : _GEN_982; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2520 = ~quene ? ram_1_77 : _GEN_983; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2521 = ~quene ? ram_1_78 : _GEN_984; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2522 = ~quene ? ram_1_79 : _GEN_985; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2523 = ~quene ? ram_1_80 : _GEN_986; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2524 = ~quene ? ram_1_81 : _GEN_987; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2525 = ~quene ? ram_1_82 : _GEN_988; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2526 = ~quene ? ram_1_83 : _GEN_989; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2527 = ~quene ? ram_1_84 : _GEN_990; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2528 = ~quene ? ram_1_85 : _GEN_991; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2529 = ~quene ? ram_1_86 : _GEN_992; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2530 = ~quene ? ram_1_87 : _GEN_993; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2531 = ~quene ? ram_1_88 : _GEN_994; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2532 = ~quene ? ram_1_89 : _GEN_995; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2533 = ~quene ? ram_1_90 : _GEN_996; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2534 = ~quene ? ram_1_91 : _GEN_997; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2535 = ~quene ? ram_1_92 : _GEN_998; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2536 = ~quene ? ram_1_93 : _GEN_999; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2537 = ~quene ? ram_1_94 : _GEN_1000; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2538 = ~quene ? ram_1_95 : _GEN_1001; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2539 = ~quene ? ram_1_96 : _GEN_1002; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2540 = ~quene ? ram_1_97 : _GEN_1003; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2541 = ~quene ? ram_1_98 : _GEN_1004; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2542 = ~quene ? ram_1_99 : _GEN_1005; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2543 = ~quene ? ram_1_100 : _GEN_1006; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2544 = ~quene ? ram_1_101 : _GEN_1007; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2545 = ~quene ? ram_1_102 : _GEN_1008; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2546 = ~quene ? ram_1_103 : _GEN_1009; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2547 = ~quene ? ram_1_104 : _GEN_1010; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2548 = ~quene ? ram_1_105 : _GEN_1011; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2549 = ~quene ? ram_1_106 : _GEN_1012; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2550 = ~quene ? ram_1_107 : _GEN_1013; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2551 = ~quene ? ram_1_108 : _GEN_1014; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2552 = ~quene ? ram_1_109 : _GEN_1015; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2553 = ~quene ? ram_1_110 : _GEN_1016; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2554 = ~quene ? ram_1_111 : _GEN_1017; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2555 = ~quene ? ram_1_112 : _GEN_1018; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2556 = ~quene ? ram_1_113 : _GEN_1019; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2557 = ~quene ? ram_1_114 : _GEN_1020; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2558 = ~quene ? ram_1_115 : _GEN_1021; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2559 = ~quene ? ram_1_116 : _GEN_1022; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2560 = ~quene ? ram_1_117 : _GEN_1023; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2561 = ~quene ? ram_1_118 : _GEN_1024; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2562 = ~quene ? ram_1_119 : _GEN_1025; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2563 = ~quene ? ram_1_120 : _GEN_1026; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2564 = ~quene ? ram_1_121 : _GEN_1027; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2565 = ~quene ? ram_1_122 : _GEN_1028; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2566 = ~quene ? ram_1_123 : _GEN_1029; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2567 = ~quene ? ram_1_124 : _GEN_1030; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2568 = ~quene ? ram_1_125 : _GEN_1031; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2569 = ~quene ? ram_1_126 : _GEN_1032; // @[cache.scala 18:24 93:34]
  wire [63:0] _GEN_2570 = ~quene ? ram_1_127 : _GEN_1033; // @[cache.scala 18:24 93:34]
  wire [31:0] _GEN_2571 = ~quene ? tag_1_0 : _GEN_1034; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2572 = ~quene ? tag_1_1 : _GEN_1035; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2573 = ~quene ? tag_1_2 : _GEN_1036; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2574 = ~quene ? tag_1_3 : _GEN_1037; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2575 = ~quene ? tag_1_4 : _GEN_1038; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2576 = ~quene ? tag_1_5 : _GEN_1039; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2577 = ~quene ? tag_1_6 : _GEN_1040; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2578 = ~quene ? tag_1_7 : _GEN_1041; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2579 = ~quene ? tag_1_8 : _GEN_1042; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2580 = ~quene ? tag_1_9 : _GEN_1043; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2581 = ~quene ? tag_1_10 : _GEN_1044; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2582 = ~quene ? tag_1_11 : _GEN_1045; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2583 = ~quene ? tag_1_12 : _GEN_1046; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2584 = ~quene ? tag_1_13 : _GEN_1047; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2585 = ~quene ? tag_1_14 : _GEN_1048; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2586 = ~quene ? tag_1_15 : _GEN_1049; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2587 = ~quene ? tag_1_16 : _GEN_1050; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2588 = ~quene ? tag_1_17 : _GEN_1051; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2589 = ~quene ? tag_1_18 : _GEN_1052; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2590 = ~quene ? tag_1_19 : _GEN_1053; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2591 = ~quene ? tag_1_20 : _GEN_1054; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2592 = ~quene ? tag_1_21 : _GEN_1055; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2593 = ~quene ? tag_1_22 : _GEN_1056; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2594 = ~quene ? tag_1_23 : _GEN_1057; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2595 = ~quene ? tag_1_24 : _GEN_1058; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2596 = ~quene ? tag_1_25 : _GEN_1059; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2597 = ~quene ? tag_1_26 : _GEN_1060; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2598 = ~quene ? tag_1_27 : _GEN_1061; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2599 = ~quene ? tag_1_28 : _GEN_1062; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2600 = ~quene ? tag_1_29 : _GEN_1063; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2601 = ~quene ? tag_1_30 : _GEN_1064; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2602 = ~quene ? tag_1_31 : _GEN_1065; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2603 = ~quene ? tag_1_32 : _GEN_1066; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2604 = ~quene ? tag_1_33 : _GEN_1067; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2605 = ~quene ? tag_1_34 : _GEN_1068; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2606 = ~quene ? tag_1_35 : _GEN_1069; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2607 = ~quene ? tag_1_36 : _GEN_1070; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2608 = ~quene ? tag_1_37 : _GEN_1071; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2609 = ~quene ? tag_1_38 : _GEN_1072; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2610 = ~quene ? tag_1_39 : _GEN_1073; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2611 = ~quene ? tag_1_40 : _GEN_1074; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2612 = ~quene ? tag_1_41 : _GEN_1075; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2613 = ~quene ? tag_1_42 : _GEN_1076; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2614 = ~quene ? tag_1_43 : _GEN_1077; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2615 = ~quene ? tag_1_44 : _GEN_1078; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2616 = ~quene ? tag_1_45 : _GEN_1079; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2617 = ~quene ? tag_1_46 : _GEN_1080; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2618 = ~quene ? tag_1_47 : _GEN_1081; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2619 = ~quene ? tag_1_48 : _GEN_1082; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2620 = ~quene ? tag_1_49 : _GEN_1083; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2621 = ~quene ? tag_1_50 : _GEN_1084; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2622 = ~quene ? tag_1_51 : _GEN_1085; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2623 = ~quene ? tag_1_52 : _GEN_1086; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2624 = ~quene ? tag_1_53 : _GEN_1087; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2625 = ~quene ? tag_1_54 : _GEN_1088; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2626 = ~quene ? tag_1_55 : _GEN_1089; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2627 = ~quene ? tag_1_56 : _GEN_1090; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2628 = ~quene ? tag_1_57 : _GEN_1091; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2629 = ~quene ? tag_1_58 : _GEN_1092; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2630 = ~quene ? tag_1_59 : _GEN_1093; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2631 = ~quene ? tag_1_60 : _GEN_1094; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2632 = ~quene ? tag_1_61 : _GEN_1095; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2633 = ~quene ? tag_1_62 : _GEN_1096; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2634 = ~quene ? tag_1_63 : _GEN_1097; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2635 = ~quene ? tag_1_64 : _GEN_1098; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2636 = ~quene ? tag_1_65 : _GEN_1099; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2637 = ~quene ? tag_1_66 : _GEN_1100; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2638 = ~quene ? tag_1_67 : _GEN_1101; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2639 = ~quene ? tag_1_68 : _GEN_1102; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2640 = ~quene ? tag_1_69 : _GEN_1103; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2641 = ~quene ? tag_1_70 : _GEN_1104; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2642 = ~quene ? tag_1_71 : _GEN_1105; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2643 = ~quene ? tag_1_72 : _GEN_1106; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2644 = ~quene ? tag_1_73 : _GEN_1107; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2645 = ~quene ? tag_1_74 : _GEN_1108; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2646 = ~quene ? tag_1_75 : _GEN_1109; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2647 = ~quene ? tag_1_76 : _GEN_1110; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2648 = ~quene ? tag_1_77 : _GEN_1111; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2649 = ~quene ? tag_1_78 : _GEN_1112; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2650 = ~quene ? tag_1_79 : _GEN_1113; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2651 = ~quene ? tag_1_80 : _GEN_1114; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2652 = ~quene ? tag_1_81 : _GEN_1115; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2653 = ~quene ? tag_1_82 : _GEN_1116; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2654 = ~quene ? tag_1_83 : _GEN_1117; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2655 = ~quene ? tag_1_84 : _GEN_1118; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2656 = ~quene ? tag_1_85 : _GEN_1119; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2657 = ~quene ? tag_1_86 : _GEN_1120; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2658 = ~quene ? tag_1_87 : _GEN_1121; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2659 = ~quene ? tag_1_88 : _GEN_1122; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2660 = ~quene ? tag_1_89 : _GEN_1123; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2661 = ~quene ? tag_1_90 : _GEN_1124; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2662 = ~quene ? tag_1_91 : _GEN_1125; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2663 = ~quene ? tag_1_92 : _GEN_1126; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2664 = ~quene ? tag_1_93 : _GEN_1127; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2665 = ~quene ? tag_1_94 : _GEN_1128; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2666 = ~quene ? tag_1_95 : _GEN_1129; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2667 = ~quene ? tag_1_96 : _GEN_1130; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2668 = ~quene ? tag_1_97 : _GEN_1131; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2669 = ~quene ? tag_1_98 : _GEN_1132; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2670 = ~quene ? tag_1_99 : _GEN_1133; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2671 = ~quene ? tag_1_100 : _GEN_1134; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2672 = ~quene ? tag_1_101 : _GEN_1135; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2673 = ~quene ? tag_1_102 : _GEN_1136; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2674 = ~quene ? tag_1_103 : _GEN_1137; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2675 = ~quene ? tag_1_104 : _GEN_1138; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2676 = ~quene ? tag_1_105 : _GEN_1139; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2677 = ~quene ? tag_1_106 : _GEN_1140; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2678 = ~quene ? tag_1_107 : _GEN_1141; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2679 = ~quene ? tag_1_108 : _GEN_1142; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2680 = ~quene ? tag_1_109 : _GEN_1143; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2681 = ~quene ? tag_1_110 : _GEN_1144; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2682 = ~quene ? tag_1_111 : _GEN_1145; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2683 = ~quene ? tag_1_112 : _GEN_1146; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2684 = ~quene ? tag_1_113 : _GEN_1147; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2685 = ~quene ? tag_1_114 : _GEN_1148; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2686 = ~quene ? tag_1_115 : _GEN_1149; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2687 = ~quene ? tag_1_116 : _GEN_1150; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2688 = ~quene ? tag_1_117 : _GEN_1151; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2689 = ~quene ? tag_1_118 : _GEN_1152; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2690 = ~quene ? tag_1_119 : _GEN_1153; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2691 = ~quene ? tag_1_120 : _GEN_1154; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2692 = ~quene ? tag_1_121 : _GEN_1155; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2693 = ~quene ? tag_1_122 : _GEN_1156; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2694 = ~quene ? tag_1_123 : _GEN_1157; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2695 = ~quene ? tag_1_124 : _GEN_1158; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2696 = ~quene ? tag_1_125 : _GEN_1159; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2697 = ~quene ? tag_1_126 : _GEN_1160; // @[cache.scala 20:24 93:34]
  wire [31:0] _GEN_2698 = ~quene ? tag_1_127 : _GEN_1161; // @[cache.scala 20:24 93:34]
  wire  _GEN_2699 = ~quene ? valid_1_0 : _GEN_1162; // @[cache.scala 22:26 93:34]
  wire  _GEN_2700 = ~quene ? valid_1_1 : _GEN_1163; // @[cache.scala 22:26 93:34]
  wire  _GEN_2701 = ~quene ? valid_1_2 : _GEN_1164; // @[cache.scala 22:26 93:34]
  wire  _GEN_2702 = ~quene ? valid_1_3 : _GEN_1165; // @[cache.scala 22:26 93:34]
  wire  _GEN_2703 = ~quene ? valid_1_4 : _GEN_1166; // @[cache.scala 22:26 93:34]
  wire  _GEN_2704 = ~quene ? valid_1_5 : _GEN_1167; // @[cache.scala 22:26 93:34]
  wire  _GEN_2705 = ~quene ? valid_1_6 : _GEN_1168; // @[cache.scala 22:26 93:34]
  wire  _GEN_2706 = ~quene ? valid_1_7 : _GEN_1169; // @[cache.scala 22:26 93:34]
  wire  _GEN_2707 = ~quene ? valid_1_8 : _GEN_1170; // @[cache.scala 22:26 93:34]
  wire  _GEN_2708 = ~quene ? valid_1_9 : _GEN_1171; // @[cache.scala 22:26 93:34]
  wire  _GEN_2709 = ~quene ? valid_1_10 : _GEN_1172; // @[cache.scala 22:26 93:34]
  wire  _GEN_2710 = ~quene ? valid_1_11 : _GEN_1173; // @[cache.scala 22:26 93:34]
  wire  _GEN_2711 = ~quene ? valid_1_12 : _GEN_1174; // @[cache.scala 22:26 93:34]
  wire  _GEN_2712 = ~quene ? valid_1_13 : _GEN_1175; // @[cache.scala 22:26 93:34]
  wire  _GEN_2713 = ~quene ? valid_1_14 : _GEN_1176; // @[cache.scala 22:26 93:34]
  wire  _GEN_2714 = ~quene ? valid_1_15 : _GEN_1177; // @[cache.scala 22:26 93:34]
  wire  _GEN_2715 = ~quene ? valid_1_16 : _GEN_1178; // @[cache.scala 22:26 93:34]
  wire  _GEN_2716 = ~quene ? valid_1_17 : _GEN_1179; // @[cache.scala 22:26 93:34]
  wire  _GEN_2717 = ~quene ? valid_1_18 : _GEN_1180; // @[cache.scala 22:26 93:34]
  wire  _GEN_2718 = ~quene ? valid_1_19 : _GEN_1181; // @[cache.scala 22:26 93:34]
  wire  _GEN_2719 = ~quene ? valid_1_20 : _GEN_1182; // @[cache.scala 22:26 93:34]
  wire  _GEN_2720 = ~quene ? valid_1_21 : _GEN_1183; // @[cache.scala 22:26 93:34]
  wire  _GEN_2721 = ~quene ? valid_1_22 : _GEN_1184; // @[cache.scala 22:26 93:34]
  wire  _GEN_2722 = ~quene ? valid_1_23 : _GEN_1185; // @[cache.scala 22:26 93:34]
  wire  _GEN_2723 = ~quene ? valid_1_24 : _GEN_1186; // @[cache.scala 22:26 93:34]
  wire  _GEN_2724 = ~quene ? valid_1_25 : _GEN_1187; // @[cache.scala 22:26 93:34]
  wire  _GEN_2725 = ~quene ? valid_1_26 : _GEN_1188; // @[cache.scala 22:26 93:34]
  wire  _GEN_2726 = ~quene ? valid_1_27 : _GEN_1189; // @[cache.scala 22:26 93:34]
  wire  _GEN_2727 = ~quene ? valid_1_28 : _GEN_1190; // @[cache.scala 22:26 93:34]
  wire  _GEN_2728 = ~quene ? valid_1_29 : _GEN_1191; // @[cache.scala 22:26 93:34]
  wire  _GEN_2729 = ~quene ? valid_1_30 : _GEN_1192; // @[cache.scala 22:26 93:34]
  wire  _GEN_2730 = ~quene ? valid_1_31 : _GEN_1193; // @[cache.scala 22:26 93:34]
  wire  _GEN_2731 = ~quene ? valid_1_32 : _GEN_1194; // @[cache.scala 22:26 93:34]
  wire  _GEN_2732 = ~quene ? valid_1_33 : _GEN_1195; // @[cache.scala 22:26 93:34]
  wire  _GEN_2733 = ~quene ? valid_1_34 : _GEN_1196; // @[cache.scala 22:26 93:34]
  wire  _GEN_2734 = ~quene ? valid_1_35 : _GEN_1197; // @[cache.scala 22:26 93:34]
  wire  _GEN_2735 = ~quene ? valid_1_36 : _GEN_1198; // @[cache.scala 22:26 93:34]
  wire  _GEN_2736 = ~quene ? valid_1_37 : _GEN_1199; // @[cache.scala 22:26 93:34]
  wire  _GEN_2737 = ~quene ? valid_1_38 : _GEN_1200; // @[cache.scala 22:26 93:34]
  wire  _GEN_2738 = ~quene ? valid_1_39 : _GEN_1201; // @[cache.scala 22:26 93:34]
  wire  _GEN_2739 = ~quene ? valid_1_40 : _GEN_1202; // @[cache.scala 22:26 93:34]
  wire  _GEN_2740 = ~quene ? valid_1_41 : _GEN_1203; // @[cache.scala 22:26 93:34]
  wire  _GEN_2741 = ~quene ? valid_1_42 : _GEN_1204; // @[cache.scala 22:26 93:34]
  wire  _GEN_2742 = ~quene ? valid_1_43 : _GEN_1205; // @[cache.scala 22:26 93:34]
  wire  _GEN_2743 = ~quene ? valid_1_44 : _GEN_1206; // @[cache.scala 22:26 93:34]
  wire  _GEN_2744 = ~quene ? valid_1_45 : _GEN_1207; // @[cache.scala 22:26 93:34]
  wire  _GEN_2745 = ~quene ? valid_1_46 : _GEN_1208; // @[cache.scala 22:26 93:34]
  wire  _GEN_2746 = ~quene ? valid_1_47 : _GEN_1209; // @[cache.scala 22:26 93:34]
  wire  _GEN_2747 = ~quene ? valid_1_48 : _GEN_1210; // @[cache.scala 22:26 93:34]
  wire  _GEN_2748 = ~quene ? valid_1_49 : _GEN_1211; // @[cache.scala 22:26 93:34]
  wire  _GEN_2749 = ~quene ? valid_1_50 : _GEN_1212; // @[cache.scala 22:26 93:34]
  wire  _GEN_2750 = ~quene ? valid_1_51 : _GEN_1213; // @[cache.scala 22:26 93:34]
  wire  _GEN_2751 = ~quene ? valid_1_52 : _GEN_1214; // @[cache.scala 22:26 93:34]
  wire  _GEN_2752 = ~quene ? valid_1_53 : _GEN_1215; // @[cache.scala 22:26 93:34]
  wire  _GEN_2753 = ~quene ? valid_1_54 : _GEN_1216; // @[cache.scala 22:26 93:34]
  wire  _GEN_2754 = ~quene ? valid_1_55 : _GEN_1217; // @[cache.scala 22:26 93:34]
  wire  _GEN_2755 = ~quene ? valid_1_56 : _GEN_1218; // @[cache.scala 22:26 93:34]
  wire  _GEN_2756 = ~quene ? valid_1_57 : _GEN_1219; // @[cache.scala 22:26 93:34]
  wire  _GEN_2757 = ~quene ? valid_1_58 : _GEN_1220; // @[cache.scala 22:26 93:34]
  wire  _GEN_2758 = ~quene ? valid_1_59 : _GEN_1221; // @[cache.scala 22:26 93:34]
  wire  _GEN_2759 = ~quene ? valid_1_60 : _GEN_1222; // @[cache.scala 22:26 93:34]
  wire  _GEN_2760 = ~quene ? valid_1_61 : _GEN_1223; // @[cache.scala 22:26 93:34]
  wire  _GEN_2761 = ~quene ? valid_1_62 : _GEN_1224; // @[cache.scala 22:26 93:34]
  wire  _GEN_2762 = ~quene ? valid_1_63 : _GEN_1225; // @[cache.scala 22:26 93:34]
  wire  _GEN_2763 = ~quene ? valid_1_64 : _GEN_1226; // @[cache.scala 22:26 93:34]
  wire  _GEN_2764 = ~quene ? valid_1_65 : _GEN_1227; // @[cache.scala 22:26 93:34]
  wire  _GEN_2765 = ~quene ? valid_1_66 : _GEN_1228; // @[cache.scala 22:26 93:34]
  wire  _GEN_2766 = ~quene ? valid_1_67 : _GEN_1229; // @[cache.scala 22:26 93:34]
  wire  _GEN_2767 = ~quene ? valid_1_68 : _GEN_1230; // @[cache.scala 22:26 93:34]
  wire  _GEN_2768 = ~quene ? valid_1_69 : _GEN_1231; // @[cache.scala 22:26 93:34]
  wire  _GEN_2769 = ~quene ? valid_1_70 : _GEN_1232; // @[cache.scala 22:26 93:34]
  wire  _GEN_2770 = ~quene ? valid_1_71 : _GEN_1233; // @[cache.scala 22:26 93:34]
  wire  _GEN_2771 = ~quene ? valid_1_72 : _GEN_1234; // @[cache.scala 22:26 93:34]
  wire  _GEN_2772 = ~quene ? valid_1_73 : _GEN_1235; // @[cache.scala 22:26 93:34]
  wire  _GEN_2773 = ~quene ? valid_1_74 : _GEN_1236; // @[cache.scala 22:26 93:34]
  wire  _GEN_2774 = ~quene ? valid_1_75 : _GEN_1237; // @[cache.scala 22:26 93:34]
  wire  _GEN_2775 = ~quene ? valid_1_76 : _GEN_1238; // @[cache.scala 22:26 93:34]
  wire  _GEN_2776 = ~quene ? valid_1_77 : _GEN_1239; // @[cache.scala 22:26 93:34]
  wire  _GEN_2777 = ~quene ? valid_1_78 : _GEN_1240; // @[cache.scala 22:26 93:34]
  wire  _GEN_2778 = ~quene ? valid_1_79 : _GEN_1241; // @[cache.scala 22:26 93:34]
  wire  _GEN_2779 = ~quene ? valid_1_80 : _GEN_1242; // @[cache.scala 22:26 93:34]
  wire  _GEN_2780 = ~quene ? valid_1_81 : _GEN_1243; // @[cache.scala 22:26 93:34]
  wire  _GEN_2781 = ~quene ? valid_1_82 : _GEN_1244; // @[cache.scala 22:26 93:34]
  wire  _GEN_2782 = ~quene ? valid_1_83 : _GEN_1245; // @[cache.scala 22:26 93:34]
  wire  _GEN_2783 = ~quene ? valid_1_84 : _GEN_1246; // @[cache.scala 22:26 93:34]
  wire  _GEN_2784 = ~quene ? valid_1_85 : _GEN_1247; // @[cache.scala 22:26 93:34]
  wire  _GEN_2785 = ~quene ? valid_1_86 : _GEN_1248; // @[cache.scala 22:26 93:34]
  wire  _GEN_2786 = ~quene ? valid_1_87 : _GEN_1249; // @[cache.scala 22:26 93:34]
  wire  _GEN_2787 = ~quene ? valid_1_88 : _GEN_1250; // @[cache.scala 22:26 93:34]
  wire  _GEN_2788 = ~quene ? valid_1_89 : _GEN_1251; // @[cache.scala 22:26 93:34]
  wire  _GEN_2789 = ~quene ? valid_1_90 : _GEN_1252; // @[cache.scala 22:26 93:34]
  wire  _GEN_2790 = ~quene ? valid_1_91 : _GEN_1253; // @[cache.scala 22:26 93:34]
  wire  _GEN_2791 = ~quene ? valid_1_92 : _GEN_1254; // @[cache.scala 22:26 93:34]
  wire  _GEN_2792 = ~quene ? valid_1_93 : _GEN_1255; // @[cache.scala 22:26 93:34]
  wire  _GEN_2793 = ~quene ? valid_1_94 : _GEN_1256; // @[cache.scala 22:26 93:34]
  wire  _GEN_2794 = ~quene ? valid_1_95 : _GEN_1257; // @[cache.scala 22:26 93:34]
  wire  _GEN_2795 = ~quene ? valid_1_96 : _GEN_1258; // @[cache.scala 22:26 93:34]
  wire  _GEN_2796 = ~quene ? valid_1_97 : _GEN_1259; // @[cache.scala 22:26 93:34]
  wire  _GEN_2797 = ~quene ? valid_1_98 : _GEN_1260; // @[cache.scala 22:26 93:34]
  wire  _GEN_2798 = ~quene ? valid_1_99 : _GEN_1261; // @[cache.scala 22:26 93:34]
  wire  _GEN_2799 = ~quene ? valid_1_100 : _GEN_1262; // @[cache.scala 22:26 93:34]
  wire  _GEN_2800 = ~quene ? valid_1_101 : _GEN_1263; // @[cache.scala 22:26 93:34]
  wire  _GEN_2801 = ~quene ? valid_1_102 : _GEN_1264; // @[cache.scala 22:26 93:34]
  wire  _GEN_2802 = ~quene ? valid_1_103 : _GEN_1265; // @[cache.scala 22:26 93:34]
  wire  _GEN_2803 = ~quene ? valid_1_104 : _GEN_1266; // @[cache.scala 22:26 93:34]
  wire  _GEN_2804 = ~quene ? valid_1_105 : _GEN_1267; // @[cache.scala 22:26 93:34]
  wire  _GEN_2805 = ~quene ? valid_1_106 : _GEN_1268; // @[cache.scala 22:26 93:34]
  wire  _GEN_2806 = ~quene ? valid_1_107 : _GEN_1269; // @[cache.scala 22:26 93:34]
  wire  _GEN_2807 = ~quene ? valid_1_108 : _GEN_1270; // @[cache.scala 22:26 93:34]
  wire  _GEN_2808 = ~quene ? valid_1_109 : _GEN_1271; // @[cache.scala 22:26 93:34]
  wire  _GEN_2809 = ~quene ? valid_1_110 : _GEN_1272; // @[cache.scala 22:26 93:34]
  wire  _GEN_2810 = ~quene ? valid_1_111 : _GEN_1273; // @[cache.scala 22:26 93:34]
  wire  _GEN_2811 = ~quene ? valid_1_112 : _GEN_1274; // @[cache.scala 22:26 93:34]
  wire  _GEN_2812 = ~quene ? valid_1_113 : _GEN_1275; // @[cache.scala 22:26 93:34]
  wire  _GEN_2813 = ~quene ? valid_1_114 : _GEN_1276; // @[cache.scala 22:26 93:34]
  wire  _GEN_2814 = ~quene ? valid_1_115 : _GEN_1277; // @[cache.scala 22:26 93:34]
  wire  _GEN_2815 = ~quene ? valid_1_116 : _GEN_1278; // @[cache.scala 22:26 93:34]
  wire  _GEN_2816 = ~quene ? valid_1_117 : _GEN_1279; // @[cache.scala 22:26 93:34]
  wire  _GEN_2817 = ~quene ? valid_1_118 : _GEN_1280; // @[cache.scala 22:26 93:34]
  wire  _GEN_2818 = ~quene ? valid_1_119 : _GEN_1281; // @[cache.scala 22:26 93:34]
  wire  _GEN_2819 = ~quene ? valid_1_120 : _GEN_1282; // @[cache.scala 22:26 93:34]
  wire  _GEN_2820 = ~quene ? valid_1_121 : _GEN_1283; // @[cache.scala 22:26 93:34]
  wire  _GEN_2821 = ~quene ? valid_1_122 : _GEN_1284; // @[cache.scala 22:26 93:34]
  wire  _GEN_2822 = ~quene ? valid_1_123 : _GEN_1285; // @[cache.scala 22:26 93:34]
  wire  _GEN_2823 = ~quene ? valid_1_124 : _GEN_1286; // @[cache.scala 22:26 93:34]
  wire  _GEN_2824 = ~quene ? valid_1_125 : _GEN_1287; // @[cache.scala 22:26 93:34]
  wire  _GEN_2825 = ~quene ? valid_1_126 : _GEN_1288; // @[cache.scala 22:26 93:34]
  wire  _GEN_2826 = ~quene ? valid_1_127 : _GEN_1289; // @[cache.scala 22:26 93:34]
  wire [63:0] _GEN_2827 = unuse_way == 2'h2 ? _GEN_906 : _GEN_2443; // @[cache.scala 87:40]
  wire [63:0] _GEN_2828 = unuse_way == 2'h2 ? _GEN_907 : _GEN_2444; // @[cache.scala 87:40]
  wire [63:0] _GEN_2829 = unuse_way == 2'h2 ? _GEN_908 : _GEN_2445; // @[cache.scala 87:40]
  wire [63:0] _GEN_2830 = unuse_way == 2'h2 ? _GEN_909 : _GEN_2446; // @[cache.scala 87:40]
  wire [63:0] _GEN_2831 = unuse_way == 2'h2 ? _GEN_910 : _GEN_2447; // @[cache.scala 87:40]
  wire [63:0] _GEN_2832 = unuse_way == 2'h2 ? _GEN_911 : _GEN_2448; // @[cache.scala 87:40]
  wire [63:0] _GEN_2833 = unuse_way == 2'h2 ? _GEN_912 : _GEN_2449; // @[cache.scala 87:40]
  wire [63:0] _GEN_2834 = unuse_way == 2'h2 ? _GEN_913 : _GEN_2450; // @[cache.scala 87:40]
  wire [63:0] _GEN_2835 = unuse_way == 2'h2 ? _GEN_914 : _GEN_2451; // @[cache.scala 87:40]
  wire [63:0] _GEN_2836 = unuse_way == 2'h2 ? _GEN_915 : _GEN_2452; // @[cache.scala 87:40]
  wire [63:0] _GEN_2837 = unuse_way == 2'h2 ? _GEN_916 : _GEN_2453; // @[cache.scala 87:40]
  wire [63:0] _GEN_2838 = unuse_way == 2'h2 ? _GEN_917 : _GEN_2454; // @[cache.scala 87:40]
  wire [63:0] _GEN_2839 = unuse_way == 2'h2 ? _GEN_918 : _GEN_2455; // @[cache.scala 87:40]
  wire [63:0] _GEN_2840 = unuse_way == 2'h2 ? _GEN_919 : _GEN_2456; // @[cache.scala 87:40]
  wire [63:0] _GEN_2841 = unuse_way == 2'h2 ? _GEN_920 : _GEN_2457; // @[cache.scala 87:40]
  wire [63:0] _GEN_2842 = unuse_way == 2'h2 ? _GEN_921 : _GEN_2458; // @[cache.scala 87:40]
  wire [63:0] _GEN_2843 = unuse_way == 2'h2 ? _GEN_922 : _GEN_2459; // @[cache.scala 87:40]
  wire [63:0] _GEN_2844 = unuse_way == 2'h2 ? _GEN_923 : _GEN_2460; // @[cache.scala 87:40]
  wire [63:0] _GEN_2845 = unuse_way == 2'h2 ? _GEN_924 : _GEN_2461; // @[cache.scala 87:40]
  wire [63:0] _GEN_2846 = unuse_way == 2'h2 ? _GEN_925 : _GEN_2462; // @[cache.scala 87:40]
  wire [63:0] _GEN_2847 = unuse_way == 2'h2 ? _GEN_926 : _GEN_2463; // @[cache.scala 87:40]
  wire [63:0] _GEN_2848 = unuse_way == 2'h2 ? _GEN_927 : _GEN_2464; // @[cache.scala 87:40]
  wire [63:0] _GEN_2849 = unuse_way == 2'h2 ? _GEN_928 : _GEN_2465; // @[cache.scala 87:40]
  wire [63:0] _GEN_2850 = unuse_way == 2'h2 ? _GEN_929 : _GEN_2466; // @[cache.scala 87:40]
  wire [63:0] _GEN_2851 = unuse_way == 2'h2 ? _GEN_930 : _GEN_2467; // @[cache.scala 87:40]
  wire [63:0] _GEN_2852 = unuse_way == 2'h2 ? _GEN_931 : _GEN_2468; // @[cache.scala 87:40]
  wire [63:0] _GEN_2853 = unuse_way == 2'h2 ? _GEN_932 : _GEN_2469; // @[cache.scala 87:40]
  wire [63:0] _GEN_2854 = unuse_way == 2'h2 ? _GEN_933 : _GEN_2470; // @[cache.scala 87:40]
  wire [63:0] _GEN_2855 = unuse_way == 2'h2 ? _GEN_934 : _GEN_2471; // @[cache.scala 87:40]
  wire [63:0] _GEN_2856 = unuse_way == 2'h2 ? _GEN_935 : _GEN_2472; // @[cache.scala 87:40]
  wire [63:0] _GEN_2857 = unuse_way == 2'h2 ? _GEN_936 : _GEN_2473; // @[cache.scala 87:40]
  wire [63:0] _GEN_2858 = unuse_way == 2'h2 ? _GEN_937 : _GEN_2474; // @[cache.scala 87:40]
  wire [63:0] _GEN_2859 = unuse_way == 2'h2 ? _GEN_938 : _GEN_2475; // @[cache.scala 87:40]
  wire [63:0] _GEN_2860 = unuse_way == 2'h2 ? _GEN_939 : _GEN_2476; // @[cache.scala 87:40]
  wire [63:0] _GEN_2861 = unuse_way == 2'h2 ? _GEN_940 : _GEN_2477; // @[cache.scala 87:40]
  wire [63:0] _GEN_2862 = unuse_way == 2'h2 ? _GEN_941 : _GEN_2478; // @[cache.scala 87:40]
  wire [63:0] _GEN_2863 = unuse_way == 2'h2 ? _GEN_942 : _GEN_2479; // @[cache.scala 87:40]
  wire [63:0] _GEN_2864 = unuse_way == 2'h2 ? _GEN_943 : _GEN_2480; // @[cache.scala 87:40]
  wire [63:0] _GEN_2865 = unuse_way == 2'h2 ? _GEN_944 : _GEN_2481; // @[cache.scala 87:40]
  wire [63:0] _GEN_2866 = unuse_way == 2'h2 ? _GEN_945 : _GEN_2482; // @[cache.scala 87:40]
  wire [63:0] _GEN_2867 = unuse_way == 2'h2 ? _GEN_946 : _GEN_2483; // @[cache.scala 87:40]
  wire [63:0] _GEN_2868 = unuse_way == 2'h2 ? _GEN_947 : _GEN_2484; // @[cache.scala 87:40]
  wire [63:0] _GEN_2869 = unuse_way == 2'h2 ? _GEN_948 : _GEN_2485; // @[cache.scala 87:40]
  wire [63:0] _GEN_2870 = unuse_way == 2'h2 ? _GEN_949 : _GEN_2486; // @[cache.scala 87:40]
  wire [63:0] _GEN_2871 = unuse_way == 2'h2 ? _GEN_950 : _GEN_2487; // @[cache.scala 87:40]
  wire [63:0] _GEN_2872 = unuse_way == 2'h2 ? _GEN_951 : _GEN_2488; // @[cache.scala 87:40]
  wire [63:0] _GEN_2873 = unuse_way == 2'h2 ? _GEN_952 : _GEN_2489; // @[cache.scala 87:40]
  wire [63:0] _GEN_2874 = unuse_way == 2'h2 ? _GEN_953 : _GEN_2490; // @[cache.scala 87:40]
  wire [63:0] _GEN_2875 = unuse_way == 2'h2 ? _GEN_954 : _GEN_2491; // @[cache.scala 87:40]
  wire [63:0] _GEN_2876 = unuse_way == 2'h2 ? _GEN_955 : _GEN_2492; // @[cache.scala 87:40]
  wire [63:0] _GEN_2877 = unuse_way == 2'h2 ? _GEN_956 : _GEN_2493; // @[cache.scala 87:40]
  wire [63:0] _GEN_2878 = unuse_way == 2'h2 ? _GEN_957 : _GEN_2494; // @[cache.scala 87:40]
  wire [63:0] _GEN_2879 = unuse_way == 2'h2 ? _GEN_958 : _GEN_2495; // @[cache.scala 87:40]
  wire [63:0] _GEN_2880 = unuse_way == 2'h2 ? _GEN_959 : _GEN_2496; // @[cache.scala 87:40]
  wire [63:0] _GEN_2881 = unuse_way == 2'h2 ? _GEN_960 : _GEN_2497; // @[cache.scala 87:40]
  wire [63:0] _GEN_2882 = unuse_way == 2'h2 ? _GEN_961 : _GEN_2498; // @[cache.scala 87:40]
  wire [63:0] _GEN_2883 = unuse_way == 2'h2 ? _GEN_962 : _GEN_2499; // @[cache.scala 87:40]
  wire [63:0] _GEN_2884 = unuse_way == 2'h2 ? _GEN_963 : _GEN_2500; // @[cache.scala 87:40]
  wire [63:0] _GEN_2885 = unuse_way == 2'h2 ? _GEN_964 : _GEN_2501; // @[cache.scala 87:40]
  wire [63:0] _GEN_2886 = unuse_way == 2'h2 ? _GEN_965 : _GEN_2502; // @[cache.scala 87:40]
  wire [63:0] _GEN_2887 = unuse_way == 2'h2 ? _GEN_966 : _GEN_2503; // @[cache.scala 87:40]
  wire [63:0] _GEN_2888 = unuse_way == 2'h2 ? _GEN_967 : _GEN_2504; // @[cache.scala 87:40]
  wire [63:0] _GEN_2889 = unuse_way == 2'h2 ? _GEN_968 : _GEN_2505; // @[cache.scala 87:40]
  wire [63:0] _GEN_2890 = unuse_way == 2'h2 ? _GEN_969 : _GEN_2506; // @[cache.scala 87:40]
  wire [63:0] _GEN_2891 = unuse_way == 2'h2 ? _GEN_970 : _GEN_2507; // @[cache.scala 87:40]
  wire [63:0] _GEN_2892 = unuse_way == 2'h2 ? _GEN_971 : _GEN_2508; // @[cache.scala 87:40]
  wire [63:0] _GEN_2893 = unuse_way == 2'h2 ? _GEN_972 : _GEN_2509; // @[cache.scala 87:40]
  wire [63:0] _GEN_2894 = unuse_way == 2'h2 ? _GEN_973 : _GEN_2510; // @[cache.scala 87:40]
  wire [63:0] _GEN_2895 = unuse_way == 2'h2 ? _GEN_974 : _GEN_2511; // @[cache.scala 87:40]
  wire [63:0] _GEN_2896 = unuse_way == 2'h2 ? _GEN_975 : _GEN_2512; // @[cache.scala 87:40]
  wire [63:0] _GEN_2897 = unuse_way == 2'h2 ? _GEN_976 : _GEN_2513; // @[cache.scala 87:40]
  wire [63:0] _GEN_2898 = unuse_way == 2'h2 ? _GEN_977 : _GEN_2514; // @[cache.scala 87:40]
  wire [63:0] _GEN_2899 = unuse_way == 2'h2 ? _GEN_978 : _GEN_2515; // @[cache.scala 87:40]
  wire [63:0] _GEN_2900 = unuse_way == 2'h2 ? _GEN_979 : _GEN_2516; // @[cache.scala 87:40]
  wire [63:0] _GEN_2901 = unuse_way == 2'h2 ? _GEN_980 : _GEN_2517; // @[cache.scala 87:40]
  wire [63:0] _GEN_2902 = unuse_way == 2'h2 ? _GEN_981 : _GEN_2518; // @[cache.scala 87:40]
  wire [63:0] _GEN_2903 = unuse_way == 2'h2 ? _GEN_982 : _GEN_2519; // @[cache.scala 87:40]
  wire [63:0] _GEN_2904 = unuse_way == 2'h2 ? _GEN_983 : _GEN_2520; // @[cache.scala 87:40]
  wire [63:0] _GEN_2905 = unuse_way == 2'h2 ? _GEN_984 : _GEN_2521; // @[cache.scala 87:40]
  wire [63:0] _GEN_2906 = unuse_way == 2'h2 ? _GEN_985 : _GEN_2522; // @[cache.scala 87:40]
  wire [63:0] _GEN_2907 = unuse_way == 2'h2 ? _GEN_986 : _GEN_2523; // @[cache.scala 87:40]
  wire [63:0] _GEN_2908 = unuse_way == 2'h2 ? _GEN_987 : _GEN_2524; // @[cache.scala 87:40]
  wire [63:0] _GEN_2909 = unuse_way == 2'h2 ? _GEN_988 : _GEN_2525; // @[cache.scala 87:40]
  wire [63:0] _GEN_2910 = unuse_way == 2'h2 ? _GEN_989 : _GEN_2526; // @[cache.scala 87:40]
  wire [63:0] _GEN_2911 = unuse_way == 2'h2 ? _GEN_990 : _GEN_2527; // @[cache.scala 87:40]
  wire [63:0] _GEN_2912 = unuse_way == 2'h2 ? _GEN_991 : _GEN_2528; // @[cache.scala 87:40]
  wire [63:0] _GEN_2913 = unuse_way == 2'h2 ? _GEN_992 : _GEN_2529; // @[cache.scala 87:40]
  wire [63:0] _GEN_2914 = unuse_way == 2'h2 ? _GEN_993 : _GEN_2530; // @[cache.scala 87:40]
  wire [63:0] _GEN_2915 = unuse_way == 2'h2 ? _GEN_994 : _GEN_2531; // @[cache.scala 87:40]
  wire [63:0] _GEN_2916 = unuse_way == 2'h2 ? _GEN_995 : _GEN_2532; // @[cache.scala 87:40]
  wire [63:0] _GEN_2917 = unuse_way == 2'h2 ? _GEN_996 : _GEN_2533; // @[cache.scala 87:40]
  wire [63:0] _GEN_2918 = unuse_way == 2'h2 ? _GEN_997 : _GEN_2534; // @[cache.scala 87:40]
  wire [63:0] _GEN_2919 = unuse_way == 2'h2 ? _GEN_998 : _GEN_2535; // @[cache.scala 87:40]
  wire [63:0] _GEN_2920 = unuse_way == 2'h2 ? _GEN_999 : _GEN_2536; // @[cache.scala 87:40]
  wire [63:0] _GEN_2921 = unuse_way == 2'h2 ? _GEN_1000 : _GEN_2537; // @[cache.scala 87:40]
  wire [63:0] _GEN_2922 = unuse_way == 2'h2 ? _GEN_1001 : _GEN_2538; // @[cache.scala 87:40]
  wire [63:0] _GEN_2923 = unuse_way == 2'h2 ? _GEN_1002 : _GEN_2539; // @[cache.scala 87:40]
  wire [63:0] _GEN_2924 = unuse_way == 2'h2 ? _GEN_1003 : _GEN_2540; // @[cache.scala 87:40]
  wire [63:0] _GEN_2925 = unuse_way == 2'h2 ? _GEN_1004 : _GEN_2541; // @[cache.scala 87:40]
  wire [63:0] _GEN_2926 = unuse_way == 2'h2 ? _GEN_1005 : _GEN_2542; // @[cache.scala 87:40]
  wire [63:0] _GEN_2927 = unuse_way == 2'h2 ? _GEN_1006 : _GEN_2543; // @[cache.scala 87:40]
  wire [63:0] _GEN_2928 = unuse_way == 2'h2 ? _GEN_1007 : _GEN_2544; // @[cache.scala 87:40]
  wire [63:0] _GEN_2929 = unuse_way == 2'h2 ? _GEN_1008 : _GEN_2545; // @[cache.scala 87:40]
  wire [63:0] _GEN_2930 = unuse_way == 2'h2 ? _GEN_1009 : _GEN_2546; // @[cache.scala 87:40]
  wire [63:0] _GEN_2931 = unuse_way == 2'h2 ? _GEN_1010 : _GEN_2547; // @[cache.scala 87:40]
  wire [63:0] _GEN_2932 = unuse_way == 2'h2 ? _GEN_1011 : _GEN_2548; // @[cache.scala 87:40]
  wire [63:0] _GEN_2933 = unuse_way == 2'h2 ? _GEN_1012 : _GEN_2549; // @[cache.scala 87:40]
  wire [63:0] _GEN_2934 = unuse_way == 2'h2 ? _GEN_1013 : _GEN_2550; // @[cache.scala 87:40]
  wire [63:0] _GEN_2935 = unuse_way == 2'h2 ? _GEN_1014 : _GEN_2551; // @[cache.scala 87:40]
  wire [63:0] _GEN_2936 = unuse_way == 2'h2 ? _GEN_1015 : _GEN_2552; // @[cache.scala 87:40]
  wire [63:0] _GEN_2937 = unuse_way == 2'h2 ? _GEN_1016 : _GEN_2553; // @[cache.scala 87:40]
  wire [63:0] _GEN_2938 = unuse_way == 2'h2 ? _GEN_1017 : _GEN_2554; // @[cache.scala 87:40]
  wire [63:0] _GEN_2939 = unuse_way == 2'h2 ? _GEN_1018 : _GEN_2555; // @[cache.scala 87:40]
  wire [63:0] _GEN_2940 = unuse_way == 2'h2 ? _GEN_1019 : _GEN_2556; // @[cache.scala 87:40]
  wire [63:0] _GEN_2941 = unuse_way == 2'h2 ? _GEN_1020 : _GEN_2557; // @[cache.scala 87:40]
  wire [63:0] _GEN_2942 = unuse_way == 2'h2 ? _GEN_1021 : _GEN_2558; // @[cache.scala 87:40]
  wire [63:0] _GEN_2943 = unuse_way == 2'h2 ? _GEN_1022 : _GEN_2559; // @[cache.scala 87:40]
  wire [63:0] _GEN_2944 = unuse_way == 2'h2 ? _GEN_1023 : _GEN_2560; // @[cache.scala 87:40]
  wire [63:0] _GEN_2945 = unuse_way == 2'h2 ? _GEN_1024 : _GEN_2561; // @[cache.scala 87:40]
  wire [63:0] _GEN_2946 = unuse_way == 2'h2 ? _GEN_1025 : _GEN_2562; // @[cache.scala 87:40]
  wire [63:0] _GEN_2947 = unuse_way == 2'h2 ? _GEN_1026 : _GEN_2563; // @[cache.scala 87:40]
  wire [63:0] _GEN_2948 = unuse_way == 2'h2 ? _GEN_1027 : _GEN_2564; // @[cache.scala 87:40]
  wire [63:0] _GEN_2949 = unuse_way == 2'h2 ? _GEN_1028 : _GEN_2565; // @[cache.scala 87:40]
  wire [63:0] _GEN_2950 = unuse_way == 2'h2 ? _GEN_1029 : _GEN_2566; // @[cache.scala 87:40]
  wire [63:0] _GEN_2951 = unuse_way == 2'h2 ? _GEN_1030 : _GEN_2567; // @[cache.scala 87:40]
  wire [63:0] _GEN_2952 = unuse_way == 2'h2 ? _GEN_1031 : _GEN_2568; // @[cache.scala 87:40]
  wire [63:0] _GEN_2953 = unuse_way == 2'h2 ? _GEN_1032 : _GEN_2569; // @[cache.scala 87:40]
  wire [63:0] _GEN_2954 = unuse_way == 2'h2 ? _GEN_1033 : _GEN_2570; // @[cache.scala 87:40]
  wire [31:0] _GEN_2955 = unuse_way == 2'h2 ? _GEN_1034 : _GEN_2571; // @[cache.scala 87:40]
  wire [31:0] _GEN_2956 = unuse_way == 2'h2 ? _GEN_1035 : _GEN_2572; // @[cache.scala 87:40]
  wire [31:0] _GEN_2957 = unuse_way == 2'h2 ? _GEN_1036 : _GEN_2573; // @[cache.scala 87:40]
  wire [31:0] _GEN_2958 = unuse_way == 2'h2 ? _GEN_1037 : _GEN_2574; // @[cache.scala 87:40]
  wire [31:0] _GEN_2959 = unuse_way == 2'h2 ? _GEN_1038 : _GEN_2575; // @[cache.scala 87:40]
  wire [31:0] _GEN_2960 = unuse_way == 2'h2 ? _GEN_1039 : _GEN_2576; // @[cache.scala 87:40]
  wire [31:0] _GEN_2961 = unuse_way == 2'h2 ? _GEN_1040 : _GEN_2577; // @[cache.scala 87:40]
  wire [31:0] _GEN_2962 = unuse_way == 2'h2 ? _GEN_1041 : _GEN_2578; // @[cache.scala 87:40]
  wire [31:0] _GEN_2963 = unuse_way == 2'h2 ? _GEN_1042 : _GEN_2579; // @[cache.scala 87:40]
  wire [31:0] _GEN_2964 = unuse_way == 2'h2 ? _GEN_1043 : _GEN_2580; // @[cache.scala 87:40]
  wire [31:0] _GEN_2965 = unuse_way == 2'h2 ? _GEN_1044 : _GEN_2581; // @[cache.scala 87:40]
  wire [31:0] _GEN_2966 = unuse_way == 2'h2 ? _GEN_1045 : _GEN_2582; // @[cache.scala 87:40]
  wire [31:0] _GEN_2967 = unuse_way == 2'h2 ? _GEN_1046 : _GEN_2583; // @[cache.scala 87:40]
  wire [31:0] _GEN_2968 = unuse_way == 2'h2 ? _GEN_1047 : _GEN_2584; // @[cache.scala 87:40]
  wire [31:0] _GEN_2969 = unuse_way == 2'h2 ? _GEN_1048 : _GEN_2585; // @[cache.scala 87:40]
  wire [31:0] _GEN_2970 = unuse_way == 2'h2 ? _GEN_1049 : _GEN_2586; // @[cache.scala 87:40]
  wire [31:0] _GEN_2971 = unuse_way == 2'h2 ? _GEN_1050 : _GEN_2587; // @[cache.scala 87:40]
  wire [31:0] _GEN_2972 = unuse_way == 2'h2 ? _GEN_1051 : _GEN_2588; // @[cache.scala 87:40]
  wire [31:0] _GEN_2973 = unuse_way == 2'h2 ? _GEN_1052 : _GEN_2589; // @[cache.scala 87:40]
  wire [31:0] _GEN_2974 = unuse_way == 2'h2 ? _GEN_1053 : _GEN_2590; // @[cache.scala 87:40]
  wire [31:0] _GEN_2975 = unuse_way == 2'h2 ? _GEN_1054 : _GEN_2591; // @[cache.scala 87:40]
  wire [31:0] _GEN_2976 = unuse_way == 2'h2 ? _GEN_1055 : _GEN_2592; // @[cache.scala 87:40]
  wire [31:0] _GEN_2977 = unuse_way == 2'h2 ? _GEN_1056 : _GEN_2593; // @[cache.scala 87:40]
  wire [31:0] _GEN_2978 = unuse_way == 2'h2 ? _GEN_1057 : _GEN_2594; // @[cache.scala 87:40]
  wire [31:0] _GEN_2979 = unuse_way == 2'h2 ? _GEN_1058 : _GEN_2595; // @[cache.scala 87:40]
  wire [31:0] _GEN_2980 = unuse_way == 2'h2 ? _GEN_1059 : _GEN_2596; // @[cache.scala 87:40]
  wire [31:0] _GEN_2981 = unuse_way == 2'h2 ? _GEN_1060 : _GEN_2597; // @[cache.scala 87:40]
  wire [31:0] _GEN_2982 = unuse_way == 2'h2 ? _GEN_1061 : _GEN_2598; // @[cache.scala 87:40]
  wire [31:0] _GEN_2983 = unuse_way == 2'h2 ? _GEN_1062 : _GEN_2599; // @[cache.scala 87:40]
  wire [31:0] _GEN_2984 = unuse_way == 2'h2 ? _GEN_1063 : _GEN_2600; // @[cache.scala 87:40]
  wire [31:0] _GEN_2985 = unuse_way == 2'h2 ? _GEN_1064 : _GEN_2601; // @[cache.scala 87:40]
  wire [31:0] _GEN_2986 = unuse_way == 2'h2 ? _GEN_1065 : _GEN_2602; // @[cache.scala 87:40]
  wire [31:0] _GEN_2987 = unuse_way == 2'h2 ? _GEN_1066 : _GEN_2603; // @[cache.scala 87:40]
  wire [31:0] _GEN_2988 = unuse_way == 2'h2 ? _GEN_1067 : _GEN_2604; // @[cache.scala 87:40]
  wire [31:0] _GEN_2989 = unuse_way == 2'h2 ? _GEN_1068 : _GEN_2605; // @[cache.scala 87:40]
  wire [31:0] _GEN_2990 = unuse_way == 2'h2 ? _GEN_1069 : _GEN_2606; // @[cache.scala 87:40]
  wire [31:0] _GEN_2991 = unuse_way == 2'h2 ? _GEN_1070 : _GEN_2607; // @[cache.scala 87:40]
  wire [31:0] _GEN_2992 = unuse_way == 2'h2 ? _GEN_1071 : _GEN_2608; // @[cache.scala 87:40]
  wire [31:0] _GEN_2993 = unuse_way == 2'h2 ? _GEN_1072 : _GEN_2609; // @[cache.scala 87:40]
  wire [31:0] _GEN_2994 = unuse_way == 2'h2 ? _GEN_1073 : _GEN_2610; // @[cache.scala 87:40]
  wire [31:0] _GEN_2995 = unuse_way == 2'h2 ? _GEN_1074 : _GEN_2611; // @[cache.scala 87:40]
  wire [31:0] _GEN_2996 = unuse_way == 2'h2 ? _GEN_1075 : _GEN_2612; // @[cache.scala 87:40]
  wire [31:0] _GEN_2997 = unuse_way == 2'h2 ? _GEN_1076 : _GEN_2613; // @[cache.scala 87:40]
  wire [31:0] _GEN_2998 = unuse_way == 2'h2 ? _GEN_1077 : _GEN_2614; // @[cache.scala 87:40]
  wire [31:0] _GEN_2999 = unuse_way == 2'h2 ? _GEN_1078 : _GEN_2615; // @[cache.scala 87:40]
  wire [31:0] _GEN_3000 = unuse_way == 2'h2 ? _GEN_1079 : _GEN_2616; // @[cache.scala 87:40]
  wire [31:0] _GEN_3001 = unuse_way == 2'h2 ? _GEN_1080 : _GEN_2617; // @[cache.scala 87:40]
  wire [31:0] _GEN_3002 = unuse_way == 2'h2 ? _GEN_1081 : _GEN_2618; // @[cache.scala 87:40]
  wire [31:0] _GEN_3003 = unuse_way == 2'h2 ? _GEN_1082 : _GEN_2619; // @[cache.scala 87:40]
  wire [31:0] _GEN_3004 = unuse_way == 2'h2 ? _GEN_1083 : _GEN_2620; // @[cache.scala 87:40]
  wire [31:0] _GEN_3005 = unuse_way == 2'h2 ? _GEN_1084 : _GEN_2621; // @[cache.scala 87:40]
  wire [31:0] _GEN_3006 = unuse_way == 2'h2 ? _GEN_1085 : _GEN_2622; // @[cache.scala 87:40]
  wire [31:0] _GEN_3007 = unuse_way == 2'h2 ? _GEN_1086 : _GEN_2623; // @[cache.scala 87:40]
  wire [31:0] _GEN_3008 = unuse_way == 2'h2 ? _GEN_1087 : _GEN_2624; // @[cache.scala 87:40]
  wire [31:0] _GEN_3009 = unuse_way == 2'h2 ? _GEN_1088 : _GEN_2625; // @[cache.scala 87:40]
  wire [31:0] _GEN_3010 = unuse_way == 2'h2 ? _GEN_1089 : _GEN_2626; // @[cache.scala 87:40]
  wire [31:0] _GEN_3011 = unuse_way == 2'h2 ? _GEN_1090 : _GEN_2627; // @[cache.scala 87:40]
  wire [31:0] _GEN_3012 = unuse_way == 2'h2 ? _GEN_1091 : _GEN_2628; // @[cache.scala 87:40]
  wire [31:0] _GEN_3013 = unuse_way == 2'h2 ? _GEN_1092 : _GEN_2629; // @[cache.scala 87:40]
  wire [31:0] _GEN_3014 = unuse_way == 2'h2 ? _GEN_1093 : _GEN_2630; // @[cache.scala 87:40]
  wire [31:0] _GEN_3015 = unuse_way == 2'h2 ? _GEN_1094 : _GEN_2631; // @[cache.scala 87:40]
  wire [31:0] _GEN_3016 = unuse_way == 2'h2 ? _GEN_1095 : _GEN_2632; // @[cache.scala 87:40]
  wire [31:0] _GEN_3017 = unuse_way == 2'h2 ? _GEN_1096 : _GEN_2633; // @[cache.scala 87:40]
  wire [31:0] _GEN_3018 = unuse_way == 2'h2 ? _GEN_1097 : _GEN_2634; // @[cache.scala 87:40]
  wire [31:0] _GEN_3019 = unuse_way == 2'h2 ? _GEN_1098 : _GEN_2635; // @[cache.scala 87:40]
  wire [31:0] _GEN_3020 = unuse_way == 2'h2 ? _GEN_1099 : _GEN_2636; // @[cache.scala 87:40]
  wire [31:0] _GEN_3021 = unuse_way == 2'h2 ? _GEN_1100 : _GEN_2637; // @[cache.scala 87:40]
  wire [31:0] _GEN_3022 = unuse_way == 2'h2 ? _GEN_1101 : _GEN_2638; // @[cache.scala 87:40]
  wire [31:0] _GEN_3023 = unuse_way == 2'h2 ? _GEN_1102 : _GEN_2639; // @[cache.scala 87:40]
  wire [31:0] _GEN_3024 = unuse_way == 2'h2 ? _GEN_1103 : _GEN_2640; // @[cache.scala 87:40]
  wire [31:0] _GEN_3025 = unuse_way == 2'h2 ? _GEN_1104 : _GEN_2641; // @[cache.scala 87:40]
  wire [31:0] _GEN_3026 = unuse_way == 2'h2 ? _GEN_1105 : _GEN_2642; // @[cache.scala 87:40]
  wire [31:0] _GEN_3027 = unuse_way == 2'h2 ? _GEN_1106 : _GEN_2643; // @[cache.scala 87:40]
  wire [31:0] _GEN_3028 = unuse_way == 2'h2 ? _GEN_1107 : _GEN_2644; // @[cache.scala 87:40]
  wire [31:0] _GEN_3029 = unuse_way == 2'h2 ? _GEN_1108 : _GEN_2645; // @[cache.scala 87:40]
  wire [31:0] _GEN_3030 = unuse_way == 2'h2 ? _GEN_1109 : _GEN_2646; // @[cache.scala 87:40]
  wire [31:0] _GEN_3031 = unuse_way == 2'h2 ? _GEN_1110 : _GEN_2647; // @[cache.scala 87:40]
  wire [31:0] _GEN_3032 = unuse_way == 2'h2 ? _GEN_1111 : _GEN_2648; // @[cache.scala 87:40]
  wire [31:0] _GEN_3033 = unuse_way == 2'h2 ? _GEN_1112 : _GEN_2649; // @[cache.scala 87:40]
  wire [31:0] _GEN_3034 = unuse_way == 2'h2 ? _GEN_1113 : _GEN_2650; // @[cache.scala 87:40]
  wire [31:0] _GEN_3035 = unuse_way == 2'h2 ? _GEN_1114 : _GEN_2651; // @[cache.scala 87:40]
  wire [31:0] _GEN_3036 = unuse_way == 2'h2 ? _GEN_1115 : _GEN_2652; // @[cache.scala 87:40]
  wire [31:0] _GEN_3037 = unuse_way == 2'h2 ? _GEN_1116 : _GEN_2653; // @[cache.scala 87:40]
  wire [31:0] _GEN_3038 = unuse_way == 2'h2 ? _GEN_1117 : _GEN_2654; // @[cache.scala 87:40]
  wire [31:0] _GEN_3039 = unuse_way == 2'h2 ? _GEN_1118 : _GEN_2655; // @[cache.scala 87:40]
  wire [31:0] _GEN_3040 = unuse_way == 2'h2 ? _GEN_1119 : _GEN_2656; // @[cache.scala 87:40]
  wire [31:0] _GEN_3041 = unuse_way == 2'h2 ? _GEN_1120 : _GEN_2657; // @[cache.scala 87:40]
  wire [31:0] _GEN_3042 = unuse_way == 2'h2 ? _GEN_1121 : _GEN_2658; // @[cache.scala 87:40]
  wire [31:0] _GEN_3043 = unuse_way == 2'h2 ? _GEN_1122 : _GEN_2659; // @[cache.scala 87:40]
  wire [31:0] _GEN_3044 = unuse_way == 2'h2 ? _GEN_1123 : _GEN_2660; // @[cache.scala 87:40]
  wire [31:0] _GEN_3045 = unuse_way == 2'h2 ? _GEN_1124 : _GEN_2661; // @[cache.scala 87:40]
  wire [31:0] _GEN_3046 = unuse_way == 2'h2 ? _GEN_1125 : _GEN_2662; // @[cache.scala 87:40]
  wire [31:0] _GEN_3047 = unuse_way == 2'h2 ? _GEN_1126 : _GEN_2663; // @[cache.scala 87:40]
  wire [31:0] _GEN_3048 = unuse_way == 2'h2 ? _GEN_1127 : _GEN_2664; // @[cache.scala 87:40]
  wire [31:0] _GEN_3049 = unuse_way == 2'h2 ? _GEN_1128 : _GEN_2665; // @[cache.scala 87:40]
  wire [31:0] _GEN_3050 = unuse_way == 2'h2 ? _GEN_1129 : _GEN_2666; // @[cache.scala 87:40]
  wire [31:0] _GEN_3051 = unuse_way == 2'h2 ? _GEN_1130 : _GEN_2667; // @[cache.scala 87:40]
  wire [31:0] _GEN_3052 = unuse_way == 2'h2 ? _GEN_1131 : _GEN_2668; // @[cache.scala 87:40]
  wire [31:0] _GEN_3053 = unuse_way == 2'h2 ? _GEN_1132 : _GEN_2669; // @[cache.scala 87:40]
  wire [31:0] _GEN_3054 = unuse_way == 2'h2 ? _GEN_1133 : _GEN_2670; // @[cache.scala 87:40]
  wire [31:0] _GEN_3055 = unuse_way == 2'h2 ? _GEN_1134 : _GEN_2671; // @[cache.scala 87:40]
  wire [31:0] _GEN_3056 = unuse_way == 2'h2 ? _GEN_1135 : _GEN_2672; // @[cache.scala 87:40]
  wire [31:0] _GEN_3057 = unuse_way == 2'h2 ? _GEN_1136 : _GEN_2673; // @[cache.scala 87:40]
  wire [31:0] _GEN_3058 = unuse_way == 2'h2 ? _GEN_1137 : _GEN_2674; // @[cache.scala 87:40]
  wire [31:0] _GEN_3059 = unuse_way == 2'h2 ? _GEN_1138 : _GEN_2675; // @[cache.scala 87:40]
  wire [31:0] _GEN_3060 = unuse_way == 2'h2 ? _GEN_1139 : _GEN_2676; // @[cache.scala 87:40]
  wire [31:0] _GEN_3061 = unuse_way == 2'h2 ? _GEN_1140 : _GEN_2677; // @[cache.scala 87:40]
  wire [31:0] _GEN_3062 = unuse_way == 2'h2 ? _GEN_1141 : _GEN_2678; // @[cache.scala 87:40]
  wire [31:0] _GEN_3063 = unuse_way == 2'h2 ? _GEN_1142 : _GEN_2679; // @[cache.scala 87:40]
  wire [31:0] _GEN_3064 = unuse_way == 2'h2 ? _GEN_1143 : _GEN_2680; // @[cache.scala 87:40]
  wire [31:0] _GEN_3065 = unuse_way == 2'h2 ? _GEN_1144 : _GEN_2681; // @[cache.scala 87:40]
  wire [31:0] _GEN_3066 = unuse_way == 2'h2 ? _GEN_1145 : _GEN_2682; // @[cache.scala 87:40]
  wire [31:0] _GEN_3067 = unuse_way == 2'h2 ? _GEN_1146 : _GEN_2683; // @[cache.scala 87:40]
  wire [31:0] _GEN_3068 = unuse_way == 2'h2 ? _GEN_1147 : _GEN_2684; // @[cache.scala 87:40]
  wire [31:0] _GEN_3069 = unuse_way == 2'h2 ? _GEN_1148 : _GEN_2685; // @[cache.scala 87:40]
  wire [31:0] _GEN_3070 = unuse_way == 2'h2 ? _GEN_1149 : _GEN_2686; // @[cache.scala 87:40]
  wire [31:0] _GEN_3071 = unuse_way == 2'h2 ? _GEN_1150 : _GEN_2687; // @[cache.scala 87:40]
  wire [31:0] _GEN_3072 = unuse_way == 2'h2 ? _GEN_1151 : _GEN_2688; // @[cache.scala 87:40]
  wire [31:0] _GEN_3073 = unuse_way == 2'h2 ? _GEN_1152 : _GEN_2689; // @[cache.scala 87:40]
  wire [31:0] _GEN_3074 = unuse_way == 2'h2 ? _GEN_1153 : _GEN_2690; // @[cache.scala 87:40]
  wire [31:0] _GEN_3075 = unuse_way == 2'h2 ? _GEN_1154 : _GEN_2691; // @[cache.scala 87:40]
  wire [31:0] _GEN_3076 = unuse_way == 2'h2 ? _GEN_1155 : _GEN_2692; // @[cache.scala 87:40]
  wire [31:0] _GEN_3077 = unuse_way == 2'h2 ? _GEN_1156 : _GEN_2693; // @[cache.scala 87:40]
  wire [31:0] _GEN_3078 = unuse_way == 2'h2 ? _GEN_1157 : _GEN_2694; // @[cache.scala 87:40]
  wire [31:0] _GEN_3079 = unuse_way == 2'h2 ? _GEN_1158 : _GEN_2695; // @[cache.scala 87:40]
  wire [31:0] _GEN_3080 = unuse_way == 2'h2 ? _GEN_1159 : _GEN_2696; // @[cache.scala 87:40]
  wire [31:0] _GEN_3081 = unuse_way == 2'h2 ? _GEN_1160 : _GEN_2697; // @[cache.scala 87:40]
  wire [31:0] _GEN_3082 = unuse_way == 2'h2 ? _GEN_1161 : _GEN_2698; // @[cache.scala 87:40]
  wire  _GEN_3083 = unuse_way == 2'h2 ? _GEN_1162 : _GEN_2699; // @[cache.scala 87:40]
  wire  _GEN_3084 = unuse_way == 2'h2 ? _GEN_1163 : _GEN_2700; // @[cache.scala 87:40]
  wire  _GEN_3085 = unuse_way == 2'h2 ? _GEN_1164 : _GEN_2701; // @[cache.scala 87:40]
  wire  _GEN_3086 = unuse_way == 2'h2 ? _GEN_1165 : _GEN_2702; // @[cache.scala 87:40]
  wire  _GEN_3087 = unuse_way == 2'h2 ? _GEN_1166 : _GEN_2703; // @[cache.scala 87:40]
  wire  _GEN_3088 = unuse_way == 2'h2 ? _GEN_1167 : _GEN_2704; // @[cache.scala 87:40]
  wire  _GEN_3089 = unuse_way == 2'h2 ? _GEN_1168 : _GEN_2705; // @[cache.scala 87:40]
  wire  _GEN_3090 = unuse_way == 2'h2 ? _GEN_1169 : _GEN_2706; // @[cache.scala 87:40]
  wire  _GEN_3091 = unuse_way == 2'h2 ? _GEN_1170 : _GEN_2707; // @[cache.scala 87:40]
  wire  _GEN_3092 = unuse_way == 2'h2 ? _GEN_1171 : _GEN_2708; // @[cache.scala 87:40]
  wire  _GEN_3093 = unuse_way == 2'h2 ? _GEN_1172 : _GEN_2709; // @[cache.scala 87:40]
  wire  _GEN_3094 = unuse_way == 2'h2 ? _GEN_1173 : _GEN_2710; // @[cache.scala 87:40]
  wire  _GEN_3095 = unuse_way == 2'h2 ? _GEN_1174 : _GEN_2711; // @[cache.scala 87:40]
  wire  _GEN_3096 = unuse_way == 2'h2 ? _GEN_1175 : _GEN_2712; // @[cache.scala 87:40]
  wire  _GEN_3097 = unuse_way == 2'h2 ? _GEN_1176 : _GEN_2713; // @[cache.scala 87:40]
  wire  _GEN_3098 = unuse_way == 2'h2 ? _GEN_1177 : _GEN_2714; // @[cache.scala 87:40]
  wire  _GEN_3099 = unuse_way == 2'h2 ? _GEN_1178 : _GEN_2715; // @[cache.scala 87:40]
  wire  _GEN_3100 = unuse_way == 2'h2 ? _GEN_1179 : _GEN_2716; // @[cache.scala 87:40]
  wire  _GEN_3101 = unuse_way == 2'h2 ? _GEN_1180 : _GEN_2717; // @[cache.scala 87:40]
  wire  _GEN_3102 = unuse_way == 2'h2 ? _GEN_1181 : _GEN_2718; // @[cache.scala 87:40]
  wire  _GEN_3103 = unuse_way == 2'h2 ? _GEN_1182 : _GEN_2719; // @[cache.scala 87:40]
  wire  _GEN_3104 = unuse_way == 2'h2 ? _GEN_1183 : _GEN_2720; // @[cache.scala 87:40]
  wire  _GEN_3105 = unuse_way == 2'h2 ? _GEN_1184 : _GEN_2721; // @[cache.scala 87:40]
  wire  _GEN_3106 = unuse_way == 2'h2 ? _GEN_1185 : _GEN_2722; // @[cache.scala 87:40]
  wire  _GEN_3107 = unuse_way == 2'h2 ? _GEN_1186 : _GEN_2723; // @[cache.scala 87:40]
  wire  _GEN_3108 = unuse_way == 2'h2 ? _GEN_1187 : _GEN_2724; // @[cache.scala 87:40]
  wire  _GEN_3109 = unuse_way == 2'h2 ? _GEN_1188 : _GEN_2725; // @[cache.scala 87:40]
  wire  _GEN_3110 = unuse_way == 2'h2 ? _GEN_1189 : _GEN_2726; // @[cache.scala 87:40]
  wire  _GEN_3111 = unuse_way == 2'h2 ? _GEN_1190 : _GEN_2727; // @[cache.scala 87:40]
  wire  _GEN_3112 = unuse_way == 2'h2 ? _GEN_1191 : _GEN_2728; // @[cache.scala 87:40]
  wire  _GEN_3113 = unuse_way == 2'h2 ? _GEN_1192 : _GEN_2729; // @[cache.scala 87:40]
  wire  _GEN_3114 = unuse_way == 2'h2 ? _GEN_1193 : _GEN_2730; // @[cache.scala 87:40]
  wire  _GEN_3115 = unuse_way == 2'h2 ? _GEN_1194 : _GEN_2731; // @[cache.scala 87:40]
  wire  _GEN_3116 = unuse_way == 2'h2 ? _GEN_1195 : _GEN_2732; // @[cache.scala 87:40]
  wire  _GEN_3117 = unuse_way == 2'h2 ? _GEN_1196 : _GEN_2733; // @[cache.scala 87:40]
  wire  _GEN_3118 = unuse_way == 2'h2 ? _GEN_1197 : _GEN_2734; // @[cache.scala 87:40]
  wire  _GEN_3119 = unuse_way == 2'h2 ? _GEN_1198 : _GEN_2735; // @[cache.scala 87:40]
  wire  _GEN_3120 = unuse_way == 2'h2 ? _GEN_1199 : _GEN_2736; // @[cache.scala 87:40]
  wire  _GEN_3121 = unuse_way == 2'h2 ? _GEN_1200 : _GEN_2737; // @[cache.scala 87:40]
  wire  _GEN_3122 = unuse_way == 2'h2 ? _GEN_1201 : _GEN_2738; // @[cache.scala 87:40]
  wire  _GEN_3123 = unuse_way == 2'h2 ? _GEN_1202 : _GEN_2739; // @[cache.scala 87:40]
  wire  _GEN_3124 = unuse_way == 2'h2 ? _GEN_1203 : _GEN_2740; // @[cache.scala 87:40]
  wire  _GEN_3125 = unuse_way == 2'h2 ? _GEN_1204 : _GEN_2741; // @[cache.scala 87:40]
  wire  _GEN_3126 = unuse_way == 2'h2 ? _GEN_1205 : _GEN_2742; // @[cache.scala 87:40]
  wire  _GEN_3127 = unuse_way == 2'h2 ? _GEN_1206 : _GEN_2743; // @[cache.scala 87:40]
  wire  _GEN_3128 = unuse_way == 2'h2 ? _GEN_1207 : _GEN_2744; // @[cache.scala 87:40]
  wire  _GEN_3129 = unuse_way == 2'h2 ? _GEN_1208 : _GEN_2745; // @[cache.scala 87:40]
  wire  _GEN_3130 = unuse_way == 2'h2 ? _GEN_1209 : _GEN_2746; // @[cache.scala 87:40]
  wire  _GEN_3131 = unuse_way == 2'h2 ? _GEN_1210 : _GEN_2747; // @[cache.scala 87:40]
  wire  _GEN_3132 = unuse_way == 2'h2 ? _GEN_1211 : _GEN_2748; // @[cache.scala 87:40]
  wire  _GEN_3133 = unuse_way == 2'h2 ? _GEN_1212 : _GEN_2749; // @[cache.scala 87:40]
  wire  _GEN_3134 = unuse_way == 2'h2 ? _GEN_1213 : _GEN_2750; // @[cache.scala 87:40]
  wire  _GEN_3135 = unuse_way == 2'h2 ? _GEN_1214 : _GEN_2751; // @[cache.scala 87:40]
  wire  _GEN_3136 = unuse_way == 2'h2 ? _GEN_1215 : _GEN_2752; // @[cache.scala 87:40]
  wire  _GEN_3137 = unuse_way == 2'h2 ? _GEN_1216 : _GEN_2753; // @[cache.scala 87:40]
  wire  _GEN_3138 = unuse_way == 2'h2 ? _GEN_1217 : _GEN_2754; // @[cache.scala 87:40]
  wire  _GEN_3139 = unuse_way == 2'h2 ? _GEN_1218 : _GEN_2755; // @[cache.scala 87:40]
  wire  _GEN_3140 = unuse_way == 2'h2 ? _GEN_1219 : _GEN_2756; // @[cache.scala 87:40]
  wire  _GEN_3141 = unuse_way == 2'h2 ? _GEN_1220 : _GEN_2757; // @[cache.scala 87:40]
  wire  _GEN_3142 = unuse_way == 2'h2 ? _GEN_1221 : _GEN_2758; // @[cache.scala 87:40]
  wire  _GEN_3143 = unuse_way == 2'h2 ? _GEN_1222 : _GEN_2759; // @[cache.scala 87:40]
  wire  _GEN_3144 = unuse_way == 2'h2 ? _GEN_1223 : _GEN_2760; // @[cache.scala 87:40]
  wire  _GEN_3145 = unuse_way == 2'h2 ? _GEN_1224 : _GEN_2761; // @[cache.scala 87:40]
  wire  _GEN_3146 = unuse_way == 2'h2 ? _GEN_1225 : _GEN_2762; // @[cache.scala 87:40]
  wire  _GEN_3147 = unuse_way == 2'h2 ? _GEN_1226 : _GEN_2763; // @[cache.scala 87:40]
  wire  _GEN_3148 = unuse_way == 2'h2 ? _GEN_1227 : _GEN_2764; // @[cache.scala 87:40]
  wire  _GEN_3149 = unuse_way == 2'h2 ? _GEN_1228 : _GEN_2765; // @[cache.scala 87:40]
  wire  _GEN_3150 = unuse_way == 2'h2 ? _GEN_1229 : _GEN_2766; // @[cache.scala 87:40]
  wire  _GEN_3151 = unuse_way == 2'h2 ? _GEN_1230 : _GEN_2767; // @[cache.scala 87:40]
  wire  _GEN_3152 = unuse_way == 2'h2 ? _GEN_1231 : _GEN_2768; // @[cache.scala 87:40]
  wire  _GEN_3153 = unuse_way == 2'h2 ? _GEN_1232 : _GEN_2769; // @[cache.scala 87:40]
  wire  _GEN_3154 = unuse_way == 2'h2 ? _GEN_1233 : _GEN_2770; // @[cache.scala 87:40]
  wire  _GEN_3155 = unuse_way == 2'h2 ? _GEN_1234 : _GEN_2771; // @[cache.scala 87:40]
  wire  _GEN_3156 = unuse_way == 2'h2 ? _GEN_1235 : _GEN_2772; // @[cache.scala 87:40]
  wire  _GEN_3157 = unuse_way == 2'h2 ? _GEN_1236 : _GEN_2773; // @[cache.scala 87:40]
  wire  _GEN_3158 = unuse_way == 2'h2 ? _GEN_1237 : _GEN_2774; // @[cache.scala 87:40]
  wire  _GEN_3159 = unuse_way == 2'h2 ? _GEN_1238 : _GEN_2775; // @[cache.scala 87:40]
  wire  _GEN_3160 = unuse_way == 2'h2 ? _GEN_1239 : _GEN_2776; // @[cache.scala 87:40]
  wire  _GEN_3161 = unuse_way == 2'h2 ? _GEN_1240 : _GEN_2777; // @[cache.scala 87:40]
  wire  _GEN_3162 = unuse_way == 2'h2 ? _GEN_1241 : _GEN_2778; // @[cache.scala 87:40]
  wire  _GEN_3163 = unuse_way == 2'h2 ? _GEN_1242 : _GEN_2779; // @[cache.scala 87:40]
  wire  _GEN_3164 = unuse_way == 2'h2 ? _GEN_1243 : _GEN_2780; // @[cache.scala 87:40]
  wire  _GEN_3165 = unuse_way == 2'h2 ? _GEN_1244 : _GEN_2781; // @[cache.scala 87:40]
  wire  _GEN_3166 = unuse_way == 2'h2 ? _GEN_1245 : _GEN_2782; // @[cache.scala 87:40]
  wire  _GEN_3167 = unuse_way == 2'h2 ? _GEN_1246 : _GEN_2783; // @[cache.scala 87:40]
  wire  _GEN_3168 = unuse_way == 2'h2 ? _GEN_1247 : _GEN_2784; // @[cache.scala 87:40]
  wire  _GEN_3169 = unuse_way == 2'h2 ? _GEN_1248 : _GEN_2785; // @[cache.scala 87:40]
  wire  _GEN_3170 = unuse_way == 2'h2 ? _GEN_1249 : _GEN_2786; // @[cache.scala 87:40]
  wire  _GEN_3171 = unuse_way == 2'h2 ? _GEN_1250 : _GEN_2787; // @[cache.scala 87:40]
  wire  _GEN_3172 = unuse_way == 2'h2 ? _GEN_1251 : _GEN_2788; // @[cache.scala 87:40]
  wire  _GEN_3173 = unuse_way == 2'h2 ? _GEN_1252 : _GEN_2789; // @[cache.scala 87:40]
  wire  _GEN_3174 = unuse_way == 2'h2 ? _GEN_1253 : _GEN_2790; // @[cache.scala 87:40]
  wire  _GEN_3175 = unuse_way == 2'h2 ? _GEN_1254 : _GEN_2791; // @[cache.scala 87:40]
  wire  _GEN_3176 = unuse_way == 2'h2 ? _GEN_1255 : _GEN_2792; // @[cache.scala 87:40]
  wire  _GEN_3177 = unuse_way == 2'h2 ? _GEN_1256 : _GEN_2793; // @[cache.scala 87:40]
  wire  _GEN_3178 = unuse_way == 2'h2 ? _GEN_1257 : _GEN_2794; // @[cache.scala 87:40]
  wire  _GEN_3179 = unuse_way == 2'h2 ? _GEN_1258 : _GEN_2795; // @[cache.scala 87:40]
  wire  _GEN_3180 = unuse_way == 2'h2 ? _GEN_1259 : _GEN_2796; // @[cache.scala 87:40]
  wire  _GEN_3181 = unuse_way == 2'h2 ? _GEN_1260 : _GEN_2797; // @[cache.scala 87:40]
  wire  _GEN_3182 = unuse_way == 2'h2 ? _GEN_1261 : _GEN_2798; // @[cache.scala 87:40]
  wire  _GEN_3183 = unuse_way == 2'h2 ? _GEN_1262 : _GEN_2799; // @[cache.scala 87:40]
  wire  _GEN_3184 = unuse_way == 2'h2 ? _GEN_1263 : _GEN_2800; // @[cache.scala 87:40]
  wire  _GEN_3185 = unuse_way == 2'h2 ? _GEN_1264 : _GEN_2801; // @[cache.scala 87:40]
  wire  _GEN_3186 = unuse_way == 2'h2 ? _GEN_1265 : _GEN_2802; // @[cache.scala 87:40]
  wire  _GEN_3187 = unuse_way == 2'h2 ? _GEN_1266 : _GEN_2803; // @[cache.scala 87:40]
  wire  _GEN_3188 = unuse_way == 2'h2 ? _GEN_1267 : _GEN_2804; // @[cache.scala 87:40]
  wire  _GEN_3189 = unuse_way == 2'h2 ? _GEN_1268 : _GEN_2805; // @[cache.scala 87:40]
  wire  _GEN_3190 = unuse_way == 2'h2 ? _GEN_1269 : _GEN_2806; // @[cache.scala 87:40]
  wire  _GEN_3191 = unuse_way == 2'h2 ? _GEN_1270 : _GEN_2807; // @[cache.scala 87:40]
  wire  _GEN_3192 = unuse_way == 2'h2 ? _GEN_1271 : _GEN_2808; // @[cache.scala 87:40]
  wire  _GEN_3193 = unuse_way == 2'h2 ? _GEN_1272 : _GEN_2809; // @[cache.scala 87:40]
  wire  _GEN_3194 = unuse_way == 2'h2 ? _GEN_1273 : _GEN_2810; // @[cache.scala 87:40]
  wire  _GEN_3195 = unuse_way == 2'h2 ? _GEN_1274 : _GEN_2811; // @[cache.scala 87:40]
  wire  _GEN_3196 = unuse_way == 2'h2 ? _GEN_1275 : _GEN_2812; // @[cache.scala 87:40]
  wire  _GEN_3197 = unuse_way == 2'h2 ? _GEN_1276 : _GEN_2813; // @[cache.scala 87:40]
  wire  _GEN_3198 = unuse_way == 2'h2 ? _GEN_1277 : _GEN_2814; // @[cache.scala 87:40]
  wire  _GEN_3199 = unuse_way == 2'h2 ? _GEN_1278 : _GEN_2815; // @[cache.scala 87:40]
  wire  _GEN_3200 = unuse_way == 2'h2 ? _GEN_1279 : _GEN_2816; // @[cache.scala 87:40]
  wire  _GEN_3201 = unuse_way == 2'h2 ? _GEN_1280 : _GEN_2817; // @[cache.scala 87:40]
  wire  _GEN_3202 = unuse_way == 2'h2 ? _GEN_1281 : _GEN_2818; // @[cache.scala 87:40]
  wire  _GEN_3203 = unuse_way == 2'h2 ? _GEN_1282 : _GEN_2819; // @[cache.scala 87:40]
  wire  _GEN_3204 = unuse_way == 2'h2 ? _GEN_1283 : _GEN_2820; // @[cache.scala 87:40]
  wire  _GEN_3205 = unuse_way == 2'h2 ? _GEN_1284 : _GEN_2821; // @[cache.scala 87:40]
  wire  _GEN_3206 = unuse_way == 2'h2 ? _GEN_1285 : _GEN_2822; // @[cache.scala 87:40]
  wire  _GEN_3207 = unuse_way == 2'h2 ? _GEN_1286 : _GEN_2823; // @[cache.scala 87:40]
  wire  _GEN_3208 = unuse_way == 2'h2 ? _GEN_1287 : _GEN_2824; // @[cache.scala 87:40]
  wire  _GEN_3209 = unuse_way == 2'h2 ? _GEN_1288 : _GEN_2825; // @[cache.scala 87:40]
  wire  _GEN_3210 = unuse_way == 2'h2 ? _GEN_1289 : _GEN_2826; // @[cache.scala 87:40]
  wire  _GEN_3211 = unuse_way == 2'h2 ? 1'h0 : _T_18; // @[cache.scala 87:40 91:23]
  wire [63:0] _GEN_3212 = unuse_way == 2'h2 ? ram_0_0 : _GEN_2058; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3213 = unuse_way == 2'h2 ? ram_0_1 : _GEN_2059; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3214 = unuse_way == 2'h2 ? ram_0_2 : _GEN_2060; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3215 = unuse_way == 2'h2 ? ram_0_3 : _GEN_2061; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3216 = unuse_way == 2'h2 ? ram_0_4 : _GEN_2062; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3217 = unuse_way == 2'h2 ? ram_0_5 : _GEN_2063; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3218 = unuse_way == 2'h2 ? ram_0_6 : _GEN_2064; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3219 = unuse_way == 2'h2 ? ram_0_7 : _GEN_2065; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3220 = unuse_way == 2'h2 ? ram_0_8 : _GEN_2066; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3221 = unuse_way == 2'h2 ? ram_0_9 : _GEN_2067; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3222 = unuse_way == 2'h2 ? ram_0_10 : _GEN_2068; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3223 = unuse_way == 2'h2 ? ram_0_11 : _GEN_2069; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3224 = unuse_way == 2'h2 ? ram_0_12 : _GEN_2070; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3225 = unuse_way == 2'h2 ? ram_0_13 : _GEN_2071; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3226 = unuse_way == 2'h2 ? ram_0_14 : _GEN_2072; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3227 = unuse_way == 2'h2 ? ram_0_15 : _GEN_2073; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3228 = unuse_way == 2'h2 ? ram_0_16 : _GEN_2074; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3229 = unuse_way == 2'h2 ? ram_0_17 : _GEN_2075; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3230 = unuse_way == 2'h2 ? ram_0_18 : _GEN_2076; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3231 = unuse_way == 2'h2 ? ram_0_19 : _GEN_2077; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3232 = unuse_way == 2'h2 ? ram_0_20 : _GEN_2078; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3233 = unuse_way == 2'h2 ? ram_0_21 : _GEN_2079; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3234 = unuse_way == 2'h2 ? ram_0_22 : _GEN_2080; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3235 = unuse_way == 2'h2 ? ram_0_23 : _GEN_2081; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3236 = unuse_way == 2'h2 ? ram_0_24 : _GEN_2082; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3237 = unuse_way == 2'h2 ? ram_0_25 : _GEN_2083; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3238 = unuse_way == 2'h2 ? ram_0_26 : _GEN_2084; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3239 = unuse_way == 2'h2 ? ram_0_27 : _GEN_2085; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3240 = unuse_way == 2'h2 ? ram_0_28 : _GEN_2086; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3241 = unuse_way == 2'h2 ? ram_0_29 : _GEN_2087; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3242 = unuse_way == 2'h2 ? ram_0_30 : _GEN_2088; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3243 = unuse_way == 2'h2 ? ram_0_31 : _GEN_2089; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3244 = unuse_way == 2'h2 ? ram_0_32 : _GEN_2090; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3245 = unuse_way == 2'h2 ? ram_0_33 : _GEN_2091; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3246 = unuse_way == 2'h2 ? ram_0_34 : _GEN_2092; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3247 = unuse_way == 2'h2 ? ram_0_35 : _GEN_2093; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3248 = unuse_way == 2'h2 ? ram_0_36 : _GEN_2094; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3249 = unuse_way == 2'h2 ? ram_0_37 : _GEN_2095; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3250 = unuse_way == 2'h2 ? ram_0_38 : _GEN_2096; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3251 = unuse_way == 2'h2 ? ram_0_39 : _GEN_2097; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3252 = unuse_way == 2'h2 ? ram_0_40 : _GEN_2098; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3253 = unuse_way == 2'h2 ? ram_0_41 : _GEN_2099; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3254 = unuse_way == 2'h2 ? ram_0_42 : _GEN_2100; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3255 = unuse_way == 2'h2 ? ram_0_43 : _GEN_2101; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3256 = unuse_way == 2'h2 ? ram_0_44 : _GEN_2102; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3257 = unuse_way == 2'h2 ? ram_0_45 : _GEN_2103; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3258 = unuse_way == 2'h2 ? ram_0_46 : _GEN_2104; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3259 = unuse_way == 2'h2 ? ram_0_47 : _GEN_2105; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3260 = unuse_way == 2'h2 ? ram_0_48 : _GEN_2106; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3261 = unuse_way == 2'h2 ? ram_0_49 : _GEN_2107; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3262 = unuse_way == 2'h2 ? ram_0_50 : _GEN_2108; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3263 = unuse_way == 2'h2 ? ram_0_51 : _GEN_2109; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3264 = unuse_way == 2'h2 ? ram_0_52 : _GEN_2110; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3265 = unuse_way == 2'h2 ? ram_0_53 : _GEN_2111; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3266 = unuse_way == 2'h2 ? ram_0_54 : _GEN_2112; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3267 = unuse_way == 2'h2 ? ram_0_55 : _GEN_2113; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3268 = unuse_way == 2'h2 ? ram_0_56 : _GEN_2114; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3269 = unuse_way == 2'h2 ? ram_0_57 : _GEN_2115; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3270 = unuse_way == 2'h2 ? ram_0_58 : _GEN_2116; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3271 = unuse_way == 2'h2 ? ram_0_59 : _GEN_2117; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3272 = unuse_way == 2'h2 ? ram_0_60 : _GEN_2118; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3273 = unuse_way == 2'h2 ? ram_0_61 : _GEN_2119; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3274 = unuse_way == 2'h2 ? ram_0_62 : _GEN_2120; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3275 = unuse_way == 2'h2 ? ram_0_63 : _GEN_2121; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3276 = unuse_way == 2'h2 ? ram_0_64 : _GEN_2122; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3277 = unuse_way == 2'h2 ? ram_0_65 : _GEN_2123; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3278 = unuse_way == 2'h2 ? ram_0_66 : _GEN_2124; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3279 = unuse_way == 2'h2 ? ram_0_67 : _GEN_2125; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3280 = unuse_way == 2'h2 ? ram_0_68 : _GEN_2126; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3281 = unuse_way == 2'h2 ? ram_0_69 : _GEN_2127; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3282 = unuse_way == 2'h2 ? ram_0_70 : _GEN_2128; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3283 = unuse_way == 2'h2 ? ram_0_71 : _GEN_2129; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3284 = unuse_way == 2'h2 ? ram_0_72 : _GEN_2130; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3285 = unuse_way == 2'h2 ? ram_0_73 : _GEN_2131; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3286 = unuse_way == 2'h2 ? ram_0_74 : _GEN_2132; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3287 = unuse_way == 2'h2 ? ram_0_75 : _GEN_2133; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3288 = unuse_way == 2'h2 ? ram_0_76 : _GEN_2134; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3289 = unuse_way == 2'h2 ? ram_0_77 : _GEN_2135; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3290 = unuse_way == 2'h2 ? ram_0_78 : _GEN_2136; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3291 = unuse_way == 2'h2 ? ram_0_79 : _GEN_2137; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3292 = unuse_way == 2'h2 ? ram_0_80 : _GEN_2138; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3293 = unuse_way == 2'h2 ? ram_0_81 : _GEN_2139; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3294 = unuse_way == 2'h2 ? ram_0_82 : _GEN_2140; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3295 = unuse_way == 2'h2 ? ram_0_83 : _GEN_2141; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3296 = unuse_way == 2'h2 ? ram_0_84 : _GEN_2142; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3297 = unuse_way == 2'h2 ? ram_0_85 : _GEN_2143; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3298 = unuse_way == 2'h2 ? ram_0_86 : _GEN_2144; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3299 = unuse_way == 2'h2 ? ram_0_87 : _GEN_2145; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3300 = unuse_way == 2'h2 ? ram_0_88 : _GEN_2146; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3301 = unuse_way == 2'h2 ? ram_0_89 : _GEN_2147; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3302 = unuse_way == 2'h2 ? ram_0_90 : _GEN_2148; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3303 = unuse_way == 2'h2 ? ram_0_91 : _GEN_2149; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3304 = unuse_way == 2'h2 ? ram_0_92 : _GEN_2150; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3305 = unuse_way == 2'h2 ? ram_0_93 : _GEN_2151; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3306 = unuse_way == 2'h2 ? ram_0_94 : _GEN_2152; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3307 = unuse_way == 2'h2 ? ram_0_95 : _GEN_2153; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3308 = unuse_way == 2'h2 ? ram_0_96 : _GEN_2154; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3309 = unuse_way == 2'h2 ? ram_0_97 : _GEN_2155; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3310 = unuse_way == 2'h2 ? ram_0_98 : _GEN_2156; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3311 = unuse_way == 2'h2 ? ram_0_99 : _GEN_2157; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3312 = unuse_way == 2'h2 ? ram_0_100 : _GEN_2158; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3313 = unuse_way == 2'h2 ? ram_0_101 : _GEN_2159; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3314 = unuse_way == 2'h2 ? ram_0_102 : _GEN_2160; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3315 = unuse_way == 2'h2 ? ram_0_103 : _GEN_2161; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3316 = unuse_way == 2'h2 ? ram_0_104 : _GEN_2162; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3317 = unuse_way == 2'h2 ? ram_0_105 : _GEN_2163; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3318 = unuse_way == 2'h2 ? ram_0_106 : _GEN_2164; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3319 = unuse_way == 2'h2 ? ram_0_107 : _GEN_2165; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3320 = unuse_way == 2'h2 ? ram_0_108 : _GEN_2166; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3321 = unuse_way == 2'h2 ? ram_0_109 : _GEN_2167; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3322 = unuse_way == 2'h2 ? ram_0_110 : _GEN_2168; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3323 = unuse_way == 2'h2 ? ram_0_111 : _GEN_2169; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3324 = unuse_way == 2'h2 ? ram_0_112 : _GEN_2170; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3325 = unuse_way == 2'h2 ? ram_0_113 : _GEN_2171; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3326 = unuse_way == 2'h2 ? ram_0_114 : _GEN_2172; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3327 = unuse_way == 2'h2 ? ram_0_115 : _GEN_2173; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3328 = unuse_way == 2'h2 ? ram_0_116 : _GEN_2174; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3329 = unuse_way == 2'h2 ? ram_0_117 : _GEN_2175; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3330 = unuse_way == 2'h2 ? ram_0_118 : _GEN_2176; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3331 = unuse_way == 2'h2 ? ram_0_119 : _GEN_2177; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3332 = unuse_way == 2'h2 ? ram_0_120 : _GEN_2178; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3333 = unuse_way == 2'h2 ? ram_0_121 : _GEN_2179; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3334 = unuse_way == 2'h2 ? ram_0_122 : _GEN_2180; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3335 = unuse_way == 2'h2 ? ram_0_123 : _GEN_2181; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3336 = unuse_way == 2'h2 ? ram_0_124 : _GEN_2182; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3337 = unuse_way == 2'h2 ? ram_0_125 : _GEN_2183; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3338 = unuse_way == 2'h2 ? ram_0_126 : _GEN_2184; // @[cache.scala 17:24 87:40]
  wire [63:0] _GEN_3339 = unuse_way == 2'h2 ? ram_0_127 : _GEN_2185; // @[cache.scala 17:24 87:40]
  wire [31:0] _GEN_3340 = unuse_way == 2'h2 ? tag_0_0 : _GEN_2186; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3341 = unuse_way == 2'h2 ? tag_0_1 : _GEN_2187; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3342 = unuse_way == 2'h2 ? tag_0_2 : _GEN_2188; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3343 = unuse_way == 2'h2 ? tag_0_3 : _GEN_2189; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3344 = unuse_way == 2'h2 ? tag_0_4 : _GEN_2190; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3345 = unuse_way == 2'h2 ? tag_0_5 : _GEN_2191; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3346 = unuse_way == 2'h2 ? tag_0_6 : _GEN_2192; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3347 = unuse_way == 2'h2 ? tag_0_7 : _GEN_2193; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3348 = unuse_way == 2'h2 ? tag_0_8 : _GEN_2194; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3349 = unuse_way == 2'h2 ? tag_0_9 : _GEN_2195; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3350 = unuse_way == 2'h2 ? tag_0_10 : _GEN_2196; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3351 = unuse_way == 2'h2 ? tag_0_11 : _GEN_2197; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3352 = unuse_way == 2'h2 ? tag_0_12 : _GEN_2198; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3353 = unuse_way == 2'h2 ? tag_0_13 : _GEN_2199; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3354 = unuse_way == 2'h2 ? tag_0_14 : _GEN_2200; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3355 = unuse_way == 2'h2 ? tag_0_15 : _GEN_2201; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3356 = unuse_way == 2'h2 ? tag_0_16 : _GEN_2202; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3357 = unuse_way == 2'h2 ? tag_0_17 : _GEN_2203; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3358 = unuse_way == 2'h2 ? tag_0_18 : _GEN_2204; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3359 = unuse_way == 2'h2 ? tag_0_19 : _GEN_2205; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3360 = unuse_way == 2'h2 ? tag_0_20 : _GEN_2206; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3361 = unuse_way == 2'h2 ? tag_0_21 : _GEN_2207; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3362 = unuse_way == 2'h2 ? tag_0_22 : _GEN_2208; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3363 = unuse_way == 2'h2 ? tag_0_23 : _GEN_2209; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3364 = unuse_way == 2'h2 ? tag_0_24 : _GEN_2210; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3365 = unuse_way == 2'h2 ? tag_0_25 : _GEN_2211; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3366 = unuse_way == 2'h2 ? tag_0_26 : _GEN_2212; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3367 = unuse_way == 2'h2 ? tag_0_27 : _GEN_2213; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3368 = unuse_way == 2'h2 ? tag_0_28 : _GEN_2214; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3369 = unuse_way == 2'h2 ? tag_0_29 : _GEN_2215; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3370 = unuse_way == 2'h2 ? tag_0_30 : _GEN_2216; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3371 = unuse_way == 2'h2 ? tag_0_31 : _GEN_2217; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3372 = unuse_way == 2'h2 ? tag_0_32 : _GEN_2218; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3373 = unuse_way == 2'h2 ? tag_0_33 : _GEN_2219; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3374 = unuse_way == 2'h2 ? tag_0_34 : _GEN_2220; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3375 = unuse_way == 2'h2 ? tag_0_35 : _GEN_2221; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3376 = unuse_way == 2'h2 ? tag_0_36 : _GEN_2222; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3377 = unuse_way == 2'h2 ? tag_0_37 : _GEN_2223; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3378 = unuse_way == 2'h2 ? tag_0_38 : _GEN_2224; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3379 = unuse_way == 2'h2 ? tag_0_39 : _GEN_2225; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3380 = unuse_way == 2'h2 ? tag_0_40 : _GEN_2226; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3381 = unuse_way == 2'h2 ? tag_0_41 : _GEN_2227; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3382 = unuse_way == 2'h2 ? tag_0_42 : _GEN_2228; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3383 = unuse_way == 2'h2 ? tag_0_43 : _GEN_2229; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3384 = unuse_way == 2'h2 ? tag_0_44 : _GEN_2230; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3385 = unuse_way == 2'h2 ? tag_0_45 : _GEN_2231; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3386 = unuse_way == 2'h2 ? tag_0_46 : _GEN_2232; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3387 = unuse_way == 2'h2 ? tag_0_47 : _GEN_2233; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3388 = unuse_way == 2'h2 ? tag_0_48 : _GEN_2234; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3389 = unuse_way == 2'h2 ? tag_0_49 : _GEN_2235; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3390 = unuse_way == 2'h2 ? tag_0_50 : _GEN_2236; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3391 = unuse_way == 2'h2 ? tag_0_51 : _GEN_2237; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3392 = unuse_way == 2'h2 ? tag_0_52 : _GEN_2238; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3393 = unuse_way == 2'h2 ? tag_0_53 : _GEN_2239; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3394 = unuse_way == 2'h2 ? tag_0_54 : _GEN_2240; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3395 = unuse_way == 2'h2 ? tag_0_55 : _GEN_2241; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3396 = unuse_way == 2'h2 ? tag_0_56 : _GEN_2242; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3397 = unuse_way == 2'h2 ? tag_0_57 : _GEN_2243; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3398 = unuse_way == 2'h2 ? tag_0_58 : _GEN_2244; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3399 = unuse_way == 2'h2 ? tag_0_59 : _GEN_2245; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3400 = unuse_way == 2'h2 ? tag_0_60 : _GEN_2246; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3401 = unuse_way == 2'h2 ? tag_0_61 : _GEN_2247; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3402 = unuse_way == 2'h2 ? tag_0_62 : _GEN_2248; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3403 = unuse_way == 2'h2 ? tag_0_63 : _GEN_2249; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3404 = unuse_way == 2'h2 ? tag_0_64 : _GEN_2250; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3405 = unuse_way == 2'h2 ? tag_0_65 : _GEN_2251; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3406 = unuse_way == 2'h2 ? tag_0_66 : _GEN_2252; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3407 = unuse_way == 2'h2 ? tag_0_67 : _GEN_2253; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3408 = unuse_way == 2'h2 ? tag_0_68 : _GEN_2254; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3409 = unuse_way == 2'h2 ? tag_0_69 : _GEN_2255; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3410 = unuse_way == 2'h2 ? tag_0_70 : _GEN_2256; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3411 = unuse_way == 2'h2 ? tag_0_71 : _GEN_2257; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3412 = unuse_way == 2'h2 ? tag_0_72 : _GEN_2258; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3413 = unuse_way == 2'h2 ? tag_0_73 : _GEN_2259; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3414 = unuse_way == 2'h2 ? tag_0_74 : _GEN_2260; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3415 = unuse_way == 2'h2 ? tag_0_75 : _GEN_2261; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3416 = unuse_way == 2'h2 ? tag_0_76 : _GEN_2262; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3417 = unuse_way == 2'h2 ? tag_0_77 : _GEN_2263; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3418 = unuse_way == 2'h2 ? tag_0_78 : _GEN_2264; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3419 = unuse_way == 2'h2 ? tag_0_79 : _GEN_2265; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3420 = unuse_way == 2'h2 ? tag_0_80 : _GEN_2266; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3421 = unuse_way == 2'h2 ? tag_0_81 : _GEN_2267; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3422 = unuse_way == 2'h2 ? tag_0_82 : _GEN_2268; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3423 = unuse_way == 2'h2 ? tag_0_83 : _GEN_2269; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3424 = unuse_way == 2'h2 ? tag_0_84 : _GEN_2270; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3425 = unuse_way == 2'h2 ? tag_0_85 : _GEN_2271; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3426 = unuse_way == 2'h2 ? tag_0_86 : _GEN_2272; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3427 = unuse_way == 2'h2 ? tag_0_87 : _GEN_2273; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3428 = unuse_way == 2'h2 ? tag_0_88 : _GEN_2274; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3429 = unuse_way == 2'h2 ? tag_0_89 : _GEN_2275; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3430 = unuse_way == 2'h2 ? tag_0_90 : _GEN_2276; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3431 = unuse_way == 2'h2 ? tag_0_91 : _GEN_2277; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3432 = unuse_way == 2'h2 ? tag_0_92 : _GEN_2278; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3433 = unuse_way == 2'h2 ? tag_0_93 : _GEN_2279; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3434 = unuse_way == 2'h2 ? tag_0_94 : _GEN_2280; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3435 = unuse_way == 2'h2 ? tag_0_95 : _GEN_2281; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3436 = unuse_way == 2'h2 ? tag_0_96 : _GEN_2282; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3437 = unuse_way == 2'h2 ? tag_0_97 : _GEN_2283; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3438 = unuse_way == 2'h2 ? tag_0_98 : _GEN_2284; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3439 = unuse_way == 2'h2 ? tag_0_99 : _GEN_2285; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3440 = unuse_way == 2'h2 ? tag_0_100 : _GEN_2286; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3441 = unuse_way == 2'h2 ? tag_0_101 : _GEN_2287; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3442 = unuse_way == 2'h2 ? tag_0_102 : _GEN_2288; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3443 = unuse_way == 2'h2 ? tag_0_103 : _GEN_2289; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3444 = unuse_way == 2'h2 ? tag_0_104 : _GEN_2290; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3445 = unuse_way == 2'h2 ? tag_0_105 : _GEN_2291; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3446 = unuse_way == 2'h2 ? tag_0_106 : _GEN_2292; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3447 = unuse_way == 2'h2 ? tag_0_107 : _GEN_2293; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3448 = unuse_way == 2'h2 ? tag_0_108 : _GEN_2294; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3449 = unuse_way == 2'h2 ? tag_0_109 : _GEN_2295; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3450 = unuse_way == 2'h2 ? tag_0_110 : _GEN_2296; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3451 = unuse_way == 2'h2 ? tag_0_111 : _GEN_2297; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3452 = unuse_way == 2'h2 ? tag_0_112 : _GEN_2298; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3453 = unuse_way == 2'h2 ? tag_0_113 : _GEN_2299; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3454 = unuse_way == 2'h2 ? tag_0_114 : _GEN_2300; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3455 = unuse_way == 2'h2 ? tag_0_115 : _GEN_2301; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3456 = unuse_way == 2'h2 ? tag_0_116 : _GEN_2302; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3457 = unuse_way == 2'h2 ? tag_0_117 : _GEN_2303; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3458 = unuse_way == 2'h2 ? tag_0_118 : _GEN_2304; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3459 = unuse_way == 2'h2 ? tag_0_119 : _GEN_2305; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3460 = unuse_way == 2'h2 ? tag_0_120 : _GEN_2306; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3461 = unuse_way == 2'h2 ? tag_0_121 : _GEN_2307; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3462 = unuse_way == 2'h2 ? tag_0_122 : _GEN_2308; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3463 = unuse_way == 2'h2 ? tag_0_123 : _GEN_2309; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3464 = unuse_way == 2'h2 ? tag_0_124 : _GEN_2310; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3465 = unuse_way == 2'h2 ? tag_0_125 : _GEN_2311; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3466 = unuse_way == 2'h2 ? tag_0_126 : _GEN_2312; // @[cache.scala 19:24 87:40]
  wire [31:0] _GEN_3467 = unuse_way == 2'h2 ? tag_0_127 : _GEN_2313; // @[cache.scala 19:24 87:40]
  wire  _GEN_3468 = unuse_way == 2'h2 ? valid_0_0 : _GEN_2314; // @[cache.scala 21:26 87:40]
  wire  _GEN_3469 = unuse_way == 2'h2 ? valid_0_1 : _GEN_2315; // @[cache.scala 21:26 87:40]
  wire  _GEN_3470 = unuse_way == 2'h2 ? valid_0_2 : _GEN_2316; // @[cache.scala 21:26 87:40]
  wire  _GEN_3471 = unuse_way == 2'h2 ? valid_0_3 : _GEN_2317; // @[cache.scala 21:26 87:40]
  wire  _GEN_3472 = unuse_way == 2'h2 ? valid_0_4 : _GEN_2318; // @[cache.scala 21:26 87:40]
  wire  _GEN_3473 = unuse_way == 2'h2 ? valid_0_5 : _GEN_2319; // @[cache.scala 21:26 87:40]
  wire  _GEN_3474 = unuse_way == 2'h2 ? valid_0_6 : _GEN_2320; // @[cache.scala 21:26 87:40]
  wire  _GEN_3475 = unuse_way == 2'h2 ? valid_0_7 : _GEN_2321; // @[cache.scala 21:26 87:40]
  wire  _GEN_3476 = unuse_way == 2'h2 ? valid_0_8 : _GEN_2322; // @[cache.scala 21:26 87:40]
  wire  _GEN_3477 = unuse_way == 2'h2 ? valid_0_9 : _GEN_2323; // @[cache.scala 21:26 87:40]
  wire  _GEN_3478 = unuse_way == 2'h2 ? valid_0_10 : _GEN_2324; // @[cache.scala 21:26 87:40]
  wire  _GEN_3479 = unuse_way == 2'h2 ? valid_0_11 : _GEN_2325; // @[cache.scala 21:26 87:40]
  wire  _GEN_3480 = unuse_way == 2'h2 ? valid_0_12 : _GEN_2326; // @[cache.scala 21:26 87:40]
  wire  _GEN_3481 = unuse_way == 2'h2 ? valid_0_13 : _GEN_2327; // @[cache.scala 21:26 87:40]
  wire  _GEN_3482 = unuse_way == 2'h2 ? valid_0_14 : _GEN_2328; // @[cache.scala 21:26 87:40]
  wire  _GEN_3483 = unuse_way == 2'h2 ? valid_0_15 : _GEN_2329; // @[cache.scala 21:26 87:40]
  wire  _GEN_3484 = unuse_way == 2'h2 ? valid_0_16 : _GEN_2330; // @[cache.scala 21:26 87:40]
  wire  _GEN_3485 = unuse_way == 2'h2 ? valid_0_17 : _GEN_2331; // @[cache.scala 21:26 87:40]
  wire  _GEN_3486 = unuse_way == 2'h2 ? valid_0_18 : _GEN_2332; // @[cache.scala 21:26 87:40]
  wire  _GEN_3487 = unuse_way == 2'h2 ? valid_0_19 : _GEN_2333; // @[cache.scala 21:26 87:40]
  wire  _GEN_3488 = unuse_way == 2'h2 ? valid_0_20 : _GEN_2334; // @[cache.scala 21:26 87:40]
  wire  _GEN_3489 = unuse_way == 2'h2 ? valid_0_21 : _GEN_2335; // @[cache.scala 21:26 87:40]
  wire  _GEN_3490 = unuse_way == 2'h2 ? valid_0_22 : _GEN_2336; // @[cache.scala 21:26 87:40]
  wire  _GEN_3491 = unuse_way == 2'h2 ? valid_0_23 : _GEN_2337; // @[cache.scala 21:26 87:40]
  wire  _GEN_3492 = unuse_way == 2'h2 ? valid_0_24 : _GEN_2338; // @[cache.scala 21:26 87:40]
  wire  _GEN_3493 = unuse_way == 2'h2 ? valid_0_25 : _GEN_2339; // @[cache.scala 21:26 87:40]
  wire  _GEN_3494 = unuse_way == 2'h2 ? valid_0_26 : _GEN_2340; // @[cache.scala 21:26 87:40]
  wire  _GEN_3495 = unuse_way == 2'h2 ? valid_0_27 : _GEN_2341; // @[cache.scala 21:26 87:40]
  wire  _GEN_3496 = unuse_way == 2'h2 ? valid_0_28 : _GEN_2342; // @[cache.scala 21:26 87:40]
  wire  _GEN_3497 = unuse_way == 2'h2 ? valid_0_29 : _GEN_2343; // @[cache.scala 21:26 87:40]
  wire  _GEN_3498 = unuse_way == 2'h2 ? valid_0_30 : _GEN_2344; // @[cache.scala 21:26 87:40]
  wire  _GEN_3499 = unuse_way == 2'h2 ? valid_0_31 : _GEN_2345; // @[cache.scala 21:26 87:40]
  wire  _GEN_3500 = unuse_way == 2'h2 ? valid_0_32 : _GEN_2346; // @[cache.scala 21:26 87:40]
  wire  _GEN_3501 = unuse_way == 2'h2 ? valid_0_33 : _GEN_2347; // @[cache.scala 21:26 87:40]
  wire  _GEN_3502 = unuse_way == 2'h2 ? valid_0_34 : _GEN_2348; // @[cache.scala 21:26 87:40]
  wire  _GEN_3503 = unuse_way == 2'h2 ? valid_0_35 : _GEN_2349; // @[cache.scala 21:26 87:40]
  wire  _GEN_3504 = unuse_way == 2'h2 ? valid_0_36 : _GEN_2350; // @[cache.scala 21:26 87:40]
  wire  _GEN_3505 = unuse_way == 2'h2 ? valid_0_37 : _GEN_2351; // @[cache.scala 21:26 87:40]
  wire  _GEN_3506 = unuse_way == 2'h2 ? valid_0_38 : _GEN_2352; // @[cache.scala 21:26 87:40]
  wire  _GEN_3507 = unuse_way == 2'h2 ? valid_0_39 : _GEN_2353; // @[cache.scala 21:26 87:40]
  wire  _GEN_3508 = unuse_way == 2'h2 ? valid_0_40 : _GEN_2354; // @[cache.scala 21:26 87:40]
  wire  _GEN_3509 = unuse_way == 2'h2 ? valid_0_41 : _GEN_2355; // @[cache.scala 21:26 87:40]
  wire  _GEN_3510 = unuse_way == 2'h2 ? valid_0_42 : _GEN_2356; // @[cache.scala 21:26 87:40]
  wire  _GEN_3511 = unuse_way == 2'h2 ? valid_0_43 : _GEN_2357; // @[cache.scala 21:26 87:40]
  wire  _GEN_3512 = unuse_way == 2'h2 ? valid_0_44 : _GEN_2358; // @[cache.scala 21:26 87:40]
  wire  _GEN_3513 = unuse_way == 2'h2 ? valid_0_45 : _GEN_2359; // @[cache.scala 21:26 87:40]
  wire  _GEN_3514 = unuse_way == 2'h2 ? valid_0_46 : _GEN_2360; // @[cache.scala 21:26 87:40]
  wire  _GEN_3515 = unuse_way == 2'h2 ? valid_0_47 : _GEN_2361; // @[cache.scala 21:26 87:40]
  wire  _GEN_3516 = unuse_way == 2'h2 ? valid_0_48 : _GEN_2362; // @[cache.scala 21:26 87:40]
  wire  _GEN_3517 = unuse_way == 2'h2 ? valid_0_49 : _GEN_2363; // @[cache.scala 21:26 87:40]
  wire  _GEN_3518 = unuse_way == 2'h2 ? valid_0_50 : _GEN_2364; // @[cache.scala 21:26 87:40]
  wire  _GEN_3519 = unuse_way == 2'h2 ? valid_0_51 : _GEN_2365; // @[cache.scala 21:26 87:40]
  wire  _GEN_3520 = unuse_way == 2'h2 ? valid_0_52 : _GEN_2366; // @[cache.scala 21:26 87:40]
  wire  _GEN_3521 = unuse_way == 2'h2 ? valid_0_53 : _GEN_2367; // @[cache.scala 21:26 87:40]
  wire  _GEN_3522 = unuse_way == 2'h2 ? valid_0_54 : _GEN_2368; // @[cache.scala 21:26 87:40]
  wire  _GEN_3523 = unuse_way == 2'h2 ? valid_0_55 : _GEN_2369; // @[cache.scala 21:26 87:40]
  wire  _GEN_3524 = unuse_way == 2'h2 ? valid_0_56 : _GEN_2370; // @[cache.scala 21:26 87:40]
  wire  _GEN_3525 = unuse_way == 2'h2 ? valid_0_57 : _GEN_2371; // @[cache.scala 21:26 87:40]
  wire  _GEN_3526 = unuse_way == 2'h2 ? valid_0_58 : _GEN_2372; // @[cache.scala 21:26 87:40]
  wire  _GEN_3527 = unuse_way == 2'h2 ? valid_0_59 : _GEN_2373; // @[cache.scala 21:26 87:40]
  wire  _GEN_3528 = unuse_way == 2'h2 ? valid_0_60 : _GEN_2374; // @[cache.scala 21:26 87:40]
  wire  _GEN_3529 = unuse_way == 2'h2 ? valid_0_61 : _GEN_2375; // @[cache.scala 21:26 87:40]
  wire  _GEN_3530 = unuse_way == 2'h2 ? valid_0_62 : _GEN_2376; // @[cache.scala 21:26 87:40]
  wire  _GEN_3531 = unuse_way == 2'h2 ? valid_0_63 : _GEN_2377; // @[cache.scala 21:26 87:40]
  wire  _GEN_3532 = unuse_way == 2'h2 ? valid_0_64 : _GEN_2378; // @[cache.scala 21:26 87:40]
  wire  _GEN_3533 = unuse_way == 2'h2 ? valid_0_65 : _GEN_2379; // @[cache.scala 21:26 87:40]
  wire  _GEN_3534 = unuse_way == 2'h2 ? valid_0_66 : _GEN_2380; // @[cache.scala 21:26 87:40]
  wire  _GEN_3535 = unuse_way == 2'h2 ? valid_0_67 : _GEN_2381; // @[cache.scala 21:26 87:40]
  wire  _GEN_3536 = unuse_way == 2'h2 ? valid_0_68 : _GEN_2382; // @[cache.scala 21:26 87:40]
  wire  _GEN_3537 = unuse_way == 2'h2 ? valid_0_69 : _GEN_2383; // @[cache.scala 21:26 87:40]
  wire  _GEN_3538 = unuse_way == 2'h2 ? valid_0_70 : _GEN_2384; // @[cache.scala 21:26 87:40]
  wire  _GEN_3539 = unuse_way == 2'h2 ? valid_0_71 : _GEN_2385; // @[cache.scala 21:26 87:40]
  wire  _GEN_3540 = unuse_way == 2'h2 ? valid_0_72 : _GEN_2386; // @[cache.scala 21:26 87:40]
  wire  _GEN_3541 = unuse_way == 2'h2 ? valid_0_73 : _GEN_2387; // @[cache.scala 21:26 87:40]
  wire  _GEN_3542 = unuse_way == 2'h2 ? valid_0_74 : _GEN_2388; // @[cache.scala 21:26 87:40]
  wire  _GEN_3543 = unuse_way == 2'h2 ? valid_0_75 : _GEN_2389; // @[cache.scala 21:26 87:40]
  wire  _GEN_3544 = unuse_way == 2'h2 ? valid_0_76 : _GEN_2390; // @[cache.scala 21:26 87:40]
  wire  _GEN_3545 = unuse_way == 2'h2 ? valid_0_77 : _GEN_2391; // @[cache.scala 21:26 87:40]
  wire  _GEN_3546 = unuse_way == 2'h2 ? valid_0_78 : _GEN_2392; // @[cache.scala 21:26 87:40]
  wire  _GEN_3547 = unuse_way == 2'h2 ? valid_0_79 : _GEN_2393; // @[cache.scala 21:26 87:40]
  wire  _GEN_3548 = unuse_way == 2'h2 ? valid_0_80 : _GEN_2394; // @[cache.scala 21:26 87:40]
  wire  _GEN_3549 = unuse_way == 2'h2 ? valid_0_81 : _GEN_2395; // @[cache.scala 21:26 87:40]
  wire  _GEN_3550 = unuse_way == 2'h2 ? valid_0_82 : _GEN_2396; // @[cache.scala 21:26 87:40]
  wire  _GEN_3551 = unuse_way == 2'h2 ? valid_0_83 : _GEN_2397; // @[cache.scala 21:26 87:40]
  wire  _GEN_3552 = unuse_way == 2'h2 ? valid_0_84 : _GEN_2398; // @[cache.scala 21:26 87:40]
  wire  _GEN_3553 = unuse_way == 2'h2 ? valid_0_85 : _GEN_2399; // @[cache.scala 21:26 87:40]
  wire  _GEN_3554 = unuse_way == 2'h2 ? valid_0_86 : _GEN_2400; // @[cache.scala 21:26 87:40]
  wire  _GEN_3555 = unuse_way == 2'h2 ? valid_0_87 : _GEN_2401; // @[cache.scala 21:26 87:40]
  wire  _GEN_3556 = unuse_way == 2'h2 ? valid_0_88 : _GEN_2402; // @[cache.scala 21:26 87:40]
  wire  _GEN_3557 = unuse_way == 2'h2 ? valid_0_89 : _GEN_2403; // @[cache.scala 21:26 87:40]
  wire  _GEN_3558 = unuse_way == 2'h2 ? valid_0_90 : _GEN_2404; // @[cache.scala 21:26 87:40]
  wire  _GEN_3559 = unuse_way == 2'h2 ? valid_0_91 : _GEN_2405; // @[cache.scala 21:26 87:40]
  wire  _GEN_3560 = unuse_way == 2'h2 ? valid_0_92 : _GEN_2406; // @[cache.scala 21:26 87:40]
  wire  _GEN_3561 = unuse_way == 2'h2 ? valid_0_93 : _GEN_2407; // @[cache.scala 21:26 87:40]
  wire  _GEN_3562 = unuse_way == 2'h2 ? valid_0_94 : _GEN_2408; // @[cache.scala 21:26 87:40]
  wire  _GEN_3563 = unuse_way == 2'h2 ? valid_0_95 : _GEN_2409; // @[cache.scala 21:26 87:40]
  wire  _GEN_3564 = unuse_way == 2'h2 ? valid_0_96 : _GEN_2410; // @[cache.scala 21:26 87:40]
  wire  _GEN_3565 = unuse_way == 2'h2 ? valid_0_97 : _GEN_2411; // @[cache.scala 21:26 87:40]
  wire  _GEN_3566 = unuse_way == 2'h2 ? valid_0_98 : _GEN_2412; // @[cache.scala 21:26 87:40]
  wire  _GEN_3567 = unuse_way == 2'h2 ? valid_0_99 : _GEN_2413; // @[cache.scala 21:26 87:40]
  wire  _GEN_3568 = unuse_way == 2'h2 ? valid_0_100 : _GEN_2414; // @[cache.scala 21:26 87:40]
  wire  _GEN_3569 = unuse_way == 2'h2 ? valid_0_101 : _GEN_2415; // @[cache.scala 21:26 87:40]
  wire  _GEN_3570 = unuse_way == 2'h2 ? valid_0_102 : _GEN_2416; // @[cache.scala 21:26 87:40]
  wire  _GEN_3571 = unuse_way == 2'h2 ? valid_0_103 : _GEN_2417; // @[cache.scala 21:26 87:40]
  wire  _GEN_3572 = unuse_way == 2'h2 ? valid_0_104 : _GEN_2418; // @[cache.scala 21:26 87:40]
  wire  _GEN_3573 = unuse_way == 2'h2 ? valid_0_105 : _GEN_2419; // @[cache.scala 21:26 87:40]
  wire  _GEN_3574 = unuse_way == 2'h2 ? valid_0_106 : _GEN_2420; // @[cache.scala 21:26 87:40]
  wire  _GEN_3575 = unuse_way == 2'h2 ? valid_0_107 : _GEN_2421; // @[cache.scala 21:26 87:40]
  wire  _GEN_3576 = unuse_way == 2'h2 ? valid_0_108 : _GEN_2422; // @[cache.scala 21:26 87:40]
  wire  _GEN_3577 = unuse_way == 2'h2 ? valid_0_109 : _GEN_2423; // @[cache.scala 21:26 87:40]
  wire  _GEN_3578 = unuse_way == 2'h2 ? valid_0_110 : _GEN_2424; // @[cache.scala 21:26 87:40]
  wire  _GEN_3579 = unuse_way == 2'h2 ? valid_0_111 : _GEN_2425; // @[cache.scala 21:26 87:40]
  wire  _GEN_3580 = unuse_way == 2'h2 ? valid_0_112 : _GEN_2426; // @[cache.scala 21:26 87:40]
  wire  _GEN_3581 = unuse_way == 2'h2 ? valid_0_113 : _GEN_2427; // @[cache.scala 21:26 87:40]
  wire  _GEN_3582 = unuse_way == 2'h2 ? valid_0_114 : _GEN_2428; // @[cache.scala 21:26 87:40]
  wire  _GEN_3583 = unuse_way == 2'h2 ? valid_0_115 : _GEN_2429; // @[cache.scala 21:26 87:40]
  wire  _GEN_3584 = unuse_way == 2'h2 ? valid_0_116 : _GEN_2430; // @[cache.scala 21:26 87:40]
  wire  _GEN_3585 = unuse_way == 2'h2 ? valid_0_117 : _GEN_2431; // @[cache.scala 21:26 87:40]
  wire  _GEN_3586 = unuse_way == 2'h2 ? valid_0_118 : _GEN_2432; // @[cache.scala 21:26 87:40]
  wire  _GEN_3587 = unuse_way == 2'h2 ? valid_0_119 : _GEN_2433; // @[cache.scala 21:26 87:40]
  wire  _GEN_3588 = unuse_way == 2'h2 ? valid_0_120 : _GEN_2434; // @[cache.scala 21:26 87:40]
  wire  _GEN_3589 = unuse_way == 2'h2 ? valid_0_121 : _GEN_2435; // @[cache.scala 21:26 87:40]
  wire  _GEN_3590 = unuse_way == 2'h2 ? valid_0_122 : _GEN_2436; // @[cache.scala 21:26 87:40]
  wire  _GEN_3591 = unuse_way == 2'h2 ? valid_0_123 : _GEN_2437; // @[cache.scala 21:26 87:40]
  wire  _GEN_3592 = unuse_way == 2'h2 ? valid_0_124 : _GEN_2438; // @[cache.scala 21:26 87:40]
  wire  _GEN_3593 = unuse_way == 2'h2 ? valid_0_125 : _GEN_2439; // @[cache.scala 21:26 87:40]
  wire  _GEN_3594 = unuse_way == 2'h2 ? valid_0_126 : _GEN_2440; // @[cache.scala 21:26 87:40]
  wire  _GEN_3595 = unuse_way == 2'h2 ? valid_0_127 : _GEN_2441; // @[cache.scala 21:26 87:40]
  wire [63:0] _GEN_3596 = unuse_way == 2'h1 ? _GEN_522 : _GEN_3212; // @[cache.scala 82:34]
  wire [63:0] _GEN_3597 = unuse_way == 2'h1 ? _GEN_523 : _GEN_3213; // @[cache.scala 82:34]
  wire [63:0] _GEN_3598 = unuse_way == 2'h1 ? _GEN_524 : _GEN_3214; // @[cache.scala 82:34]
  wire [63:0] _GEN_3599 = unuse_way == 2'h1 ? _GEN_525 : _GEN_3215; // @[cache.scala 82:34]
  wire [63:0] _GEN_3600 = unuse_way == 2'h1 ? _GEN_526 : _GEN_3216; // @[cache.scala 82:34]
  wire [63:0] _GEN_3601 = unuse_way == 2'h1 ? _GEN_527 : _GEN_3217; // @[cache.scala 82:34]
  wire [63:0] _GEN_3602 = unuse_way == 2'h1 ? _GEN_528 : _GEN_3218; // @[cache.scala 82:34]
  wire [63:0] _GEN_3603 = unuse_way == 2'h1 ? _GEN_529 : _GEN_3219; // @[cache.scala 82:34]
  wire [63:0] _GEN_3604 = unuse_way == 2'h1 ? _GEN_530 : _GEN_3220; // @[cache.scala 82:34]
  wire [63:0] _GEN_3605 = unuse_way == 2'h1 ? _GEN_531 : _GEN_3221; // @[cache.scala 82:34]
  wire [63:0] _GEN_3606 = unuse_way == 2'h1 ? _GEN_532 : _GEN_3222; // @[cache.scala 82:34]
  wire [63:0] _GEN_3607 = unuse_way == 2'h1 ? _GEN_533 : _GEN_3223; // @[cache.scala 82:34]
  wire [63:0] _GEN_3608 = unuse_way == 2'h1 ? _GEN_534 : _GEN_3224; // @[cache.scala 82:34]
  wire [63:0] _GEN_3609 = unuse_way == 2'h1 ? _GEN_535 : _GEN_3225; // @[cache.scala 82:34]
  wire [63:0] _GEN_3610 = unuse_way == 2'h1 ? _GEN_536 : _GEN_3226; // @[cache.scala 82:34]
  wire [63:0] _GEN_3611 = unuse_way == 2'h1 ? _GEN_537 : _GEN_3227; // @[cache.scala 82:34]
  wire [63:0] _GEN_3612 = unuse_way == 2'h1 ? _GEN_538 : _GEN_3228; // @[cache.scala 82:34]
  wire [63:0] _GEN_3613 = unuse_way == 2'h1 ? _GEN_539 : _GEN_3229; // @[cache.scala 82:34]
  wire [63:0] _GEN_3614 = unuse_way == 2'h1 ? _GEN_540 : _GEN_3230; // @[cache.scala 82:34]
  wire [63:0] _GEN_3615 = unuse_way == 2'h1 ? _GEN_541 : _GEN_3231; // @[cache.scala 82:34]
  wire [63:0] _GEN_3616 = unuse_way == 2'h1 ? _GEN_542 : _GEN_3232; // @[cache.scala 82:34]
  wire [63:0] _GEN_3617 = unuse_way == 2'h1 ? _GEN_543 : _GEN_3233; // @[cache.scala 82:34]
  wire [63:0] _GEN_3618 = unuse_way == 2'h1 ? _GEN_544 : _GEN_3234; // @[cache.scala 82:34]
  wire [63:0] _GEN_3619 = unuse_way == 2'h1 ? _GEN_545 : _GEN_3235; // @[cache.scala 82:34]
  wire [63:0] _GEN_3620 = unuse_way == 2'h1 ? _GEN_546 : _GEN_3236; // @[cache.scala 82:34]
  wire [63:0] _GEN_3621 = unuse_way == 2'h1 ? _GEN_547 : _GEN_3237; // @[cache.scala 82:34]
  wire [63:0] _GEN_3622 = unuse_way == 2'h1 ? _GEN_548 : _GEN_3238; // @[cache.scala 82:34]
  wire [63:0] _GEN_3623 = unuse_way == 2'h1 ? _GEN_549 : _GEN_3239; // @[cache.scala 82:34]
  wire [63:0] _GEN_3624 = unuse_way == 2'h1 ? _GEN_550 : _GEN_3240; // @[cache.scala 82:34]
  wire [63:0] _GEN_3625 = unuse_way == 2'h1 ? _GEN_551 : _GEN_3241; // @[cache.scala 82:34]
  wire [63:0] _GEN_3626 = unuse_way == 2'h1 ? _GEN_552 : _GEN_3242; // @[cache.scala 82:34]
  wire [63:0] _GEN_3627 = unuse_way == 2'h1 ? _GEN_553 : _GEN_3243; // @[cache.scala 82:34]
  wire [63:0] _GEN_3628 = unuse_way == 2'h1 ? _GEN_554 : _GEN_3244; // @[cache.scala 82:34]
  wire [63:0] _GEN_3629 = unuse_way == 2'h1 ? _GEN_555 : _GEN_3245; // @[cache.scala 82:34]
  wire [63:0] _GEN_3630 = unuse_way == 2'h1 ? _GEN_556 : _GEN_3246; // @[cache.scala 82:34]
  wire [63:0] _GEN_3631 = unuse_way == 2'h1 ? _GEN_557 : _GEN_3247; // @[cache.scala 82:34]
  wire [63:0] _GEN_3632 = unuse_way == 2'h1 ? _GEN_558 : _GEN_3248; // @[cache.scala 82:34]
  wire [63:0] _GEN_3633 = unuse_way == 2'h1 ? _GEN_559 : _GEN_3249; // @[cache.scala 82:34]
  wire [63:0] _GEN_3634 = unuse_way == 2'h1 ? _GEN_560 : _GEN_3250; // @[cache.scala 82:34]
  wire [63:0] _GEN_3635 = unuse_way == 2'h1 ? _GEN_561 : _GEN_3251; // @[cache.scala 82:34]
  wire [63:0] _GEN_3636 = unuse_way == 2'h1 ? _GEN_562 : _GEN_3252; // @[cache.scala 82:34]
  wire [63:0] _GEN_3637 = unuse_way == 2'h1 ? _GEN_563 : _GEN_3253; // @[cache.scala 82:34]
  wire [63:0] _GEN_3638 = unuse_way == 2'h1 ? _GEN_564 : _GEN_3254; // @[cache.scala 82:34]
  wire [63:0] _GEN_3639 = unuse_way == 2'h1 ? _GEN_565 : _GEN_3255; // @[cache.scala 82:34]
  wire [63:0] _GEN_3640 = unuse_way == 2'h1 ? _GEN_566 : _GEN_3256; // @[cache.scala 82:34]
  wire [63:0] _GEN_3641 = unuse_way == 2'h1 ? _GEN_567 : _GEN_3257; // @[cache.scala 82:34]
  wire [63:0] _GEN_3642 = unuse_way == 2'h1 ? _GEN_568 : _GEN_3258; // @[cache.scala 82:34]
  wire [63:0] _GEN_3643 = unuse_way == 2'h1 ? _GEN_569 : _GEN_3259; // @[cache.scala 82:34]
  wire [63:0] _GEN_3644 = unuse_way == 2'h1 ? _GEN_570 : _GEN_3260; // @[cache.scala 82:34]
  wire [63:0] _GEN_3645 = unuse_way == 2'h1 ? _GEN_571 : _GEN_3261; // @[cache.scala 82:34]
  wire [63:0] _GEN_3646 = unuse_way == 2'h1 ? _GEN_572 : _GEN_3262; // @[cache.scala 82:34]
  wire [63:0] _GEN_3647 = unuse_way == 2'h1 ? _GEN_573 : _GEN_3263; // @[cache.scala 82:34]
  wire [63:0] _GEN_3648 = unuse_way == 2'h1 ? _GEN_574 : _GEN_3264; // @[cache.scala 82:34]
  wire [63:0] _GEN_3649 = unuse_way == 2'h1 ? _GEN_575 : _GEN_3265; // @[cache.scala 82:34]
  wire [63:0] _GEN_3650 = unuse_way == 2'h1 ? _GEN_576 : _GEN_3266; // @[cache.scala 82:34]
  wire [63:0] _GEN_3651 = unuse_way == 2'h1 ? _GEN_577 : _GEN_3267; // @[cache.scala 82:34]
  wire [63:0] _GEN_3652 = unuse_way == 2'h1 ? _GEN_578 : _GEN_3268; // @[cache.scala 82:34]
  wire [63:0] _GEN_3653 = unuse_way == 2'h1 ? _GEN_579 : _GEN_3269; // @[cache.scala 82:34]
  wire [63:0] _GEN_3654 = unuse_way == 2'h1 ? _GEN_580 : _GEN_3270; // @[cache.scala 82:34]
  wire [63:0] _GEN_3655 = unuse_way == 2'h1 ? _GEN_581 : _GEN_3271; // @[cache.scala 82:34]
  wire [63:0] _GEN_3656 = unuse_way == 2'h1 ? _GEN_582 : _GEN_3272; // @[cache.scala 82:34]
  wire [63:0] _GEN_3657 = unuse_way == 2'h1 ? _GEN_583 : _GEN_3273; // @[cache.scala 82:34]
  wire [63:0] _GEN_3658 = unuse_way == 2'h1 ? _GEN_584 : _GEN_3274; // @[cache.scala 82:34]
  wire [63:0] _GEN_3659 = unuse_way == 2'h1 ? _GEN_585 : _GEN_3275; // @[cache.scala 82:34]
  wire [63:0] _GEN_3660 = unuse_way == 2'h1 ? _GEN_586 : _GEN_3276; // @[cache.scala 82:34]
  wire [63:0] _GEN_3661 = unuse_way == 2'h1 ? _GEN_587 : _GEN_3277; // @[cache.scala 82:34]
  wire [63:0] _GEN_3662 = unuse_way == 2'h1 ? _GEN_588 : _GEN_3278; // @[cache.scala 82:34]
  wire [63:0] _GEN_3663 = unuse_way == 2'h1 ? _GEN_589 : _GEN_3279; // @[cache.scala 82:34]
  wire [63:0] _GEN_3664 = unuse_way == 2'h1 ? _GEN_590 : _GEN_3280; // @[cache.scala 82:34]
  wire [63:0] _GEN_3665 = unuse_way == 2'h1 ? _GEN_591 : _GEN_3281; // @[cache.scala 82:34]
  wire [63:0] _GEN_3666 = unuse_way == 2'h1 ? _GEN_592 : _GEN_3282; // @[cache.scala 82:34]
  wire [63:0] _GEN_3667 = unuse_way == 2'h1 ? _GEN_593 : _GEN_3283; // @[cache.scala 82:34]
  wire [63:0] _GEN_3668 = unuse_way == 2'h1 ? _GEN_594 : _GEN_3284; // @[cache.scala 82:34]
  wire [63:0] _GEN_3669 = unuse_way == 2'h1 ? _GEN_595 : _GEN_3285; // @[cache.scala 82:34]
  wire [63:0] _GEN_3670 = unuse_way == 2'h1 ? _GEN_596 : _GEN_3286; // @[cache.scala 82:34]
  wire [63:0] _GEN_3671 = unuse_way == 2'h1 ? _GEN_597 : _GEN_3287; // @[cache.scala 82:34]
  wire [63:0] _GEN_3672 = unuse_way == 2'h1 ? _GEN_598 : _GEN_3288; // @[cache.scala 82:34]
  wire [63:0] _GEN_3673 = unuse_way == 2'h1 ? _GEN_599 : _GEN_3289; // @[cache.scala 82:34]
  wire [63:0] _GEN_3674 = unuse_way == 2'h1 ? _GEN_600 : _GEN_3290; // @[cache.scala 82:34]
  wire [63:0] _GEN_3675 = unuse_way == 2'h1 ? _GEN_601 : _GEN_3291; // @[cache.scala 82:34]
  wire [63:0] _GEN_3676 = unuse_way == 2'h1 ? _GEN_602 : _GEN_3292; // @[cache.scala 82:34]
  wire [63:0] _GEN_3677 = unuse_way == 2'h1 ? _GEN_603 : _GEN_3293; // @[cache.scala 82:34]
  wire [63:0] _GEN_3678 = unuse_way == 2'h1 ? _GEN_604 : _GEN_3294; // @[cache.scala 82:34]
  wire [63:0] _GEN_3679 = unuse_way == 2'h1 ? _GEN_605 : _GEN_3295; // @[cache.scala 82:34]
  wire [63:0] _GEN_3680 = unuse_way == 2'h1 ? _GEN_606 : _GEN_3296; // @[cache.scala 82:34]
  wire [63:0] _GEN_3681 = unuse_way == 2'h1 ? _GEN_607 : _GEN_3297; // @[cache.scala 82:34]
  wire [63:0] _GEN_3682 = unuse_way == 2'h1 ? _GEN_608 : _GEN_3298; // @[cache.scala 82:34]
  wire [63:0] _GEN_3683 = unuse_way == 2'h1 ? _GEN_609 : _GEN_3299; // @[cache.scala 82:34]
  wire [63:0] _GEN_3684 = unuse_way == 2'h1 ? _GEN_610 : _GEN_3300; // @[cache.scala 82:34]
  wire [63:0] _GEN_3685 = unuse_way == 2'h1 ? _GEN_611 : _GEN_3301; // @[cache.scala 82:34]
  wire [63:0] _GEN_3686 = unuse_way == 2'h1 ? _GEN_612 : _GEN_3302; // @[cache.scala 82:34]
  wire [63:0] _GEN_3687 = unuse_way == 2'h1 ? _GEN_613 : _GEN_3303; // @[cache.scala 82:34]
  wire [63:0] _GEN_3688 = unuse_way == 2'h1 ? _GEN_614 : _GEN_3304; // @[cache.scala 82:34]
  wire [63:0] _GEN_3689 = unuse_way == 2'h1 ? _GEN_615 : _GEN_3305; // @[cache.scala 82:34]
  wire [63:0] _GEN_3690 = unuse_way == 2'h1 ? _GEN_616 : _GEN_3306; // @[cache.scala 82:34]
  wire [63:0] _GEN_3691 = unuse_way == 2'h1 ? _GEN_617 : _GEN_3307; // @[cache.scala 82:34]
  wire [63:0] _GEN_3692 = unuse_way == 2'h1 ? _GEN_618 : _GEN_3308; // @[cache.scala 82:34]
  wire [63:0] _GEN_3693 = unuse_way == 2'h1 ? _GEN_619 : _GEN_3309; // @[cache.scala 82:34]
  wire [63:0] _GEN_3694 = unuse_way == 2'h1 ? _GEN_620 : _GEN_3310; // @[cache.scala 82:34]
  wire [63:0] _GEN_3695 = unuse_way == 2'h1 ? _GEN_621 : _GEN_3311; // @[cache.scala 82:34]
  wire [63:0] _GEN_3696 = unuse_way == 2'h1 ? _GEN_622 : _GEN_3312; // @[cache.scala 82:34]
  wire [63:0] _GEN_3697 = unuse_way == 2'h1 ? _GEN_623 : _GEN_3313; // @[cache.scala 82:34]
  wire [63:0] _GEN_3698 = unuse_way == 2'h1 ? _GEN_624 : _GEN_3314; // @[cache.scala 82:34]
  wire [63:0] _GEN_3699 = unuse_way == 2'h1 ? _GEN_625 : _GEN_3315; // @[cache.scala 82:34]
  wire [63:0] _GEN_3700 = unuse_way == 2'h1 ? _GEN_626 : _GEN_3316; // @[cache.scala 82:34]
  wire [63:0] _GEN_3701 = unuse_way == 2'h1 ? _GEN_627 : _GEN_3317; // @[cache.scala 82:34]
  wire [63:0] _GEN_3702 = unuse_way == 2'h1 ? _GEN_628 : _GEN_3318; // @[cache.scala 82:34]
  wire [63:0] _GEN_3703 = unuse_way == 2'h1 ? _GEN_629 : _GEN_3319; // @[cache.scala 82:34]
  wire [63:0] _GEN_3704 = unuse_way == 2'h1 ? _GEN_630 : _GEN_3320; // @[cache.scala 82:34]
  wire [63:0] _GEN_3705 = unuse_way == 2'h1 ? _GEN_631 : _GEN_3321; // @[cache.scala 82:34]
  wire [63:0] _GEN_3706 = unuse_way == 2'h1 ? _GEN_632 : _GEN_3322; // @[cache.scala 82:34]
  wire [63:0] _GEN_3707 = unuse_way == 2'h1 ? _GEN_633 : _GEN_3323; // @[cache.scala 82:34]
  wire [63:0] _GEN_3708 = unuse_way == 2'h1 ? _GEN_634 : _GEN_3324; // @[cache.scala 82:34]
  wire [63:0] _GEN_3709 = unuse_way == 2'h1 ? _GEN_635 : _GEN_3325; // @[cache.scala 82:34]
  wire [63:0] _GEN_3710 = unuse_way == 2'h1 ? _GEN_636 : _GEN_3326; // @[cache.scala 82:34]
  wire [63:0] _GEN_3711 = unuse_way == 2'h1 ? _GEN_637 : _GEN_3327; // @[cache.scala 82:34]
  wire [63:0] _GEN_3712 = unuse_way == 2'h1 ? _GEN_638 : _GEN_3328; // @[cache.scala 82:34]
  wire [63:0] _GEN_3713 = unuse_way == 2'h1 ? _GEN_639 : _GEN_3329; // @[cache.scala 82:34]
  wire [63:0] _GEN_3714 = unuse_way == 2'h1 ? _GEN_640 : _GEN_3330; // @[cache.scala 82:34]
  wire [63:0] _GEN_3715 = unuse_way == 2'h1 ? _GEN_641 : _GEN_3331; // @[cache.scala 82:34]
  wire [63:0] _GEN_3716 = unuse_way == 2'h1 ? _GEN_642 : _GEN_3332; // @[cache.scala 82:34]
  wire [63:0] _GEN_3717 = unuse_way == 2'h1 ? _GEN_643 : _GEN_3333; // @[cache.scala 82:34]
  wire [63:0] _GEN_3718 = unuse_way == 2'h1 ? _GEN_644 : _GEN_3334; // @[cache.scala 82:34]
  wire [63:0] _GEN_3719 = unuse_way == 2'h1 ? _GEN_645 : _GEN_3335; // @[cache.scala 82:34]
  wire [63:0] _GEN_3720 = unuse_way == 2'h1 ? _GEN_646 : _GEN_3336; // @[cache.scala 82:34]
  wire [63:0] _GEN_3721 = unuse_way == 2'h1 ? _GEN_647 : _GEN_3337; // @[cache.scala 82:34]
  wire [63:0] _GEN_3722 = unuse_way == 2'h1 ? _GEN_648 : _GEN_3338; // @[cache.scala 82:34]
  wire [63:0] _GEN_3723 = unuse_way == 2'h1 ? _GEN_649 : _GEN_3339; // @[cache.scala 82:34]
  wire [31:0] _GEN_3724 = unuse_way == 2'h1 ? _GEN_650 : _GEN_3340; // @[cache.scala 82:34]
  wire [31:0] _GEN_3725 = unuse_way == 2'h1 ? _GEN_651 : _GEN_3341; // @[cache.scala 82:34]
  wire [31:0] _GEN_3726 = unuse_way == 2'h1 ? _GEN_652 : _GEN_3342; // @[cache.scala 82:34]
  wire [31:0] _GEN_3727 = unuse_way == 2'h1 ? _GEN_653 : _GEN_3343; // @[cache.scala 82:34]
  wire [31:0] _GEN_3728 = unuse_way == 2'h1 ? _GEN_654 : _GEN_3344; // @[cache.scala 82:34]
  wire [31:0] _GEN_3729 = unuse_way == 2'h1 ? _GEN_655 : _GEN_3345; // @[cache.scala 82:34]
  wire [31:0] _GEN_3730 = unuse_way == 2'h1 ? _GEN_656 : _GEN_3346; // @[cache.scala 82:34]
  wire [31:0] _GEN_3731 = unuse_way == 2'h1 ? _GEN_657 : _GEN_3347; // @[cache.scala 82:34]
  wire [31:0] _GEN_3732 = unuse_way == 2'h1 ? _GEN_658 : _GEN_3348; // @[cache.scala 82:34]
  wire [31:0] _GEN_3733 = unuse_way == 2'h1 ? _GEN_659 : _GEN_3349; // @[cache.scala 82:34]
  wire [31:0] _GEN_3734 = unuse_way == 2'h1 ? _GEN_660 : _GEN_3350; // @[cache.scala 82:34]
  wire [31:0] _GEN_3735 = unuse_way == 2'h1 ? _GEN_661 : _GEN_3351; // @[cache.scala 82:34]
  wire [31:0] _GEN_3736 = unuse_way == 2'h1 ? _GEN_662 : _GEN_3352; // @[cache.scala 82:34]
  wire [31:0] _GEN_3737 = unuse_way == 2'h1 ? _GEN_663 : _GEN_3353; // @[cache.scala 82:34]
  wire [31:0] _GEN_3738 = unuse_way == 2'h1 ? _GEN_664 : _GEN_3354; // @[cache.scala 82:34]
  wire [31:0] _GEN_3739 = unuse_way == 2'h1 ? _GEN_665 : _GEN_3355; // @[cache.scala 82:34]
  wire [31:0] _GEN_3740 = unuse_way == 2'h1 ? _GEN_666 : _GEN_3356; // @[cache.scala 82:34]
  wire [31:0] _GEN_3741 = unuse_way == 2'h1 ? _GEN_667 : _GEN_3357; // @[cache.scala 82:34]
  wire [31:0] _GEN_3742 = unuse_way == 2'h1 ? _GEN_668 : _GEN_3358; // @[cache.scala 82:34]
  wire [31:0] _GEN_3743 = unuse_way == 2'h1 ? _GEN_669 : _GEN_3359; // @[cache.scala 82:34]
  wire [31:0] _GEN_3744 = unuse_way == 2'h1 ? _GEN_670 : _GEN_3360; // @[cache.scala 82:34]
  wire [31:0] _GEN_3745 = unuse_way == 2'h1 ? _GEN_671 : _GEN_3361; // @[cache.scala 82:34]
  wire [31:0] _GEN_3746 = unuse_way == 2'h1 ? _GEN_672 : _GEN_3362; // @[cache.scala 82:34]
  wire [31:0] _GEN_3747 = unuse_way == 2'h1 ? _GEN_673 : _GEN_3363; // @[cache.scala 82:34]
  wire [31:0] _GEN_3748 = unuse_way == 2'h1 ? _GEN_674 : _GEN_3364; // @[cache.scala 82:34]
  wire [31:0] _GEN_3749 = unuse_way == 2'h1 ? _GEN_675 : _GEN_3365; // @[cache.scala 82:34]
  wire [31:0] _GEN_3750 = unuse_way == 2'h1 ? _GEN_676 : _GEN_3366; // @[cache.scala 82:34]
  wire [31:0] _GEN_3751 = unuse_way == 2'h1 ? _GEN_677 : _GEN_3367; // @[cache.scala 82:34]
  wire [31:0] _GEN_3752 = unuse_way == 2'h1 ? _GEN_678 : _GEN_3368; // @[cache.scala 82:34]
  wire [31:0] _GEN_3753 = unuse_way == 2'h1 ? _GEN_679 : _GEN_3369; // @[cache.scala 82:34]
  wire [31:0] _GEN_3754 = unuse_way == 2'h1 ? _GEN_680 : _GEN_3370; // @[cache.scala 82:34]
  wire [31:0] _GEN_3755 = unuse_way == 2'h1 ? _GEN_681 : _GEN_3371; // @[cache.scala 82:34]
  wire [31:0] _GEN_3756 = unuse_way == 2'h1 ? _GEN_682 : _GEN_3372; // @[cache.scala 82:34]
  wire [31:0] _GEN_3757 = unuse_way == 2'h1 ? _GEN_683 : _GEN_3373; // @[cache.scala 82:34]
  wire [31:0] _GEN_3758 = unuse_way == 2'h1 ? _GEN_684 : _GEN_3374; // @[cache.scala 82:34]
  wire [31:0] _GEN_3759 = unuse_way == 2'h1 ? _GEN_685 : _GEN_3375; // @[cache.scala 82:34]
  wire [31:0] _GEN_3760 = unuse_way == 2'h1 ? _GEN_686 : _GEN_3376; // @[cache.scala 82:34]
  wire [31:0] _GEN_3761 = unuse_way == 2'h1 ? _GEN_687 : _GEN_3377; // @[cache.scala 82:34]
  wire [31:0] _GEN_3762 = unuse_way == 2'h1 ? _GEN_688 : _GEN_3378; // @[cache.scala 82:34]
  wire [31:0] _GEN_3763 = unuse_way == 2'h1 ? _GEN_689 : _GEN_3379; // @[cache.scala 82:34]
  wire [31:0] _GEN_3764 = unuse_way == 2'h1 ? _GEN_690 : _GEN_3380; // @[cache.scala 82:34]
  wire [31:0] _GEN_3765 = unuse_way == 2'h1 ? _GEN_691 : _GEN_3381; // @[cache.scala 82:34]
  wire [31:0] _GEN_3766 = unuse_way == 2'h1 ? _GEN_692 : _GEN_3382; // @[cache.scala 82:34]
  wire [31:0] _GEN_3767 = unuse_way == 2'h1 ? _GEN_693 : _GEN_3383; // @[cache.scala 82:34]
  wire [31:0] _GEN_3768 = unuse_way == 2'h1 ? _GEN_694 : _GEN_3384; // @[cache.scala 82:34]
  wire [31:0] _GEN_3769 = unuse_way == 2'h1 ? _GEN_695 : _GEN_3385; // @[cache.scala 82:34]
  wire [31:0] _GEN_3770 = unuse_way == 2'h1 ? _GEN_696 : _GEN_3386; // @[cache.scala 82:34]
  wire [31:0] _GEN_3771 = unuse_way == 2'h1 ? _GEN_697 : _GEN_3387; // @[cache.scala 82:34]
  wire [31:0] _GEN_3772 = unuse_way == 2'h1 ? _GEN_698 : _GEN_3388; // @[cache.scala 82:34]
  wire [31:0] _GEN_3773 = unuse_way == 2'h1 ? _GEN_699 : _GEN_3389; // @[cache.scala 82:34]
  wire [31:0] _GEN_3774 = unuse_way == 2'h1 ? _GEN_700 : _GEN_3390; // @[cache.scala 82:34]
  wire [31:0] _GEN_3775 = unuse_way == 2'h1 ? _GEN_701 : _GEN_3391; // @[cache.scala 82:34]
  wire [31:0] _GEN_3776 = unuse_way == 2'h1 ? _GEN_702 : _GEN_3392; // @[cache.scala 82:34]
  wire [31:0] _GEN_3777 = unuse_way == 2'h1 ? _GEN_703 : _GEN_3393; // @[cache.scala 82:34]
  wire [31:0] _GEN_3778 = unuse_way == 2'h1 ? _GEN_704 : _GEN_3394; // @[cache.scala 82:34]
  wire [31:0] _GEN_3779 = unuse_way == 2'h1 ? _GEN_705 : _GEN_3395; // @[cache.scala 82:34]
  wire [31:0] _GEN_3780 = unuse_way == 2'h1 ? _GEN_706 : _GEN_3396; // @[cache.scala 82:34]
  wire [31:0] _GEN_3781 = unuse_way == 2'h1 ? _GEN_707 : _GEN_3397; // @[cache.scala 82:34]
  wire [31:0] _GEN_3782 = unuse_way == 2'h1 ? _GEN_708 : _GEN_3398; // @[cache.scala 82:34]
  wire [31:0] _GEN_3783 = unuse_way == 2'h1 ? _GEN_709 : _GEN_3399; // @[cache.scala 82:34]
  wire [31:0] _GEN_3784 = unuse_way == 2'h1 ? _GEN_710 : _GEN_3400; // @[cache.scala 82:34]
  wire [31:0] _GEN_3785 = unuse_way == 2'h1 ? _GEN_711 : _GEN_3401; // @[cache.scala 82:34]
  wire [31:0] _GEN_3786 = unuse_way == 2'h1 ? _GEN_712 : _GEN_3402; // @[cache.scala 82:34]
  wire [31:0] _GEN_3787 = unuse_way == 2'h1 ? _GEN_713 : _GEN_3403; // @[cache.scala 82:34]
  wire [31:0] _GEN_3788 = unuse_way == 2'h1 ? _GEN_714 : _GEN_3404; // @[cache.scala 82:34]
  wire [31:0] _GEN_3789 = unuse_way == 2'h1 ? _GEN_715 : _GEN_3405; // @[cache.scala 82:34]
  wire [31:0] _GEN_3790 = unuse_way == 2'h1 ? _GEN_716 : _GEN_3406; // @[cache.scala 82:34]
  wire [31:0] _GEN_3791 = unuse_way == 2'h1 ? _GEN_717 : _GEN_3407; // @[cache.scala 82:34]
  wire [31:0] _GEN_3792 = unuse_way == 2'h1 ? _GEN_718 : _GEN_3408; // @[cache.scala 82:34]
  wire [31:0] _GEN_3793 = unuse_way == 2'h1 ? _GEN_719 : _GEN_3409; // @[cache.scala 82:34]
  wire [31:0] _GEN_3794 = unuse_way == 2'h1 ? _GEN_720 : _GEN_3410; // @[cache.scala 82:34]
  wire [31:0] _GEN_3795 = unuse_way == 2'h1 ? _GEN_721 : _GEN_3411; // @[cache.scala 82:34]
  wire [31:0] _GEN_3796 = unuse_way == 2'h1 ? _GEN_722 : _GEN_3412; // @[cache.scala 82:34]
  wire [31:0] _GEN_3797 = unuse_way == 2'h1 ? _GEN_723 : _GEN_3413; // @[cache.scala 82:34]
  wire [31:0] _GEN_3798 = unuse_way == 2'h1 ? _GEN_724 : _GEN_3414; // @[cache.scala 82:34]
  wire [31:0] _GEN_3799 = unuse_way == 2'h1 ? _GEN_725 : _GEN_3415; // @[cache.scala 82:34]
  wire [31:0] _GEN_3800 = unuse_way == 2'h1 ? _GEN_726 : _GEN_3416; // @[cache.scala 82:34]
  wire [31:0] _GEN_3801 = unuse_way == 2'h1 ? _GEN_727 : _GEN_3417; // @[cache.scala 82:34]
  wire [31:0] _GEN_3802 = unuse_way == 2'h1 ? _GEN_728 : _GEN_3418; // @[cache.scala 82:34]
  wire [31:0] _GEN_3803 = unuse_way == 2'h1 ? _GEN_729 : _GEN_3419; // @[cache.scala 82:34]
  wire [31:0] _GEN_3804 = unuse_way == 2'h1 ? _GEN_730 : _GEN_3420; // @[cache.scala 82:34]
  wire [31:0] _GEN_3805 = unuse_way == 2'h1 ? _GEN_731 : _GEN_3421; // @[cache.scala 82:34]
  wire [31:0] _GEN_3806 = unuse_way == 2'h1 ? _GEN_732 : _GEN_3422; // @[cache.scala 82:34]
  wire [31:0] _GEN_3807 = unuse_way == 2'h1 ? _GEN_733 : _GEN_3423; // @[cache.scala 82:34]
  wire [31:0] _GEN_3808 = unuse_way == 2'h1 ? _GEN_734 : _GEN_3424; // @[cache.scala 82:34]
  wire [31:0] _GEN_3809 = unuse_way == 2'h1 ? _GEN_735 : _GEN_3425; // @[cache.scala 82:34]
  wire [31:0] _GEN_3810 = unuse_way == 2'h1 ? _GEN_736 : _GEN_3426; // @[cache.scala 82:34]
  wire [31:0] _GEN_3811 = unuse_way == 2'h1 ? _GEN_737 : _GEN_3427; // @[cache.scala 82:34]
  wire [31:0] _GEN_3812 = unuse_way == 2'h1 ? _GEN_738 : _GEN_3428; // @[cache.scala 82:34]
  wire [31:0] _GEN_3813 = unuse_way == 2'h1 ? _GEN_739 : _GEN_3429; // @[cache.scala 82:34]
  wire [31:0] _GEN_3814 = unuse_way == 2'h1 ? _GEN_740 : _GEN_3430; // @[cache.scala 82:34]
  wire [31:0] _GEN_3815 = unuse_way == 2'h1 ? _GEN_741 : _GEN_3431; // @[cache.scala 82:34]
  wire [31:0] _GEN_3816 = unuse_way == 2'h1 ? _GEN_742 : _GEN_3432; // @[cache.scala 82:34]
  wire [31:0] _GEN_3817 = unuse_way == 2'h1 ? _GEN_743 : _GEN_3433; // @[cache.scala 82:34]
  wire [31:0] _GEN_3818 = unuse_way == 2'h1 ? _GEN_744 : _GEN_3434; // @[cache.scala 82:34]
  wire [31:0] _GEN_3819 = unuse_way == 2'h1 ? _GEN_745 : _GEN_3435; // @[cache.scala 82:34]
  wire [31:0] _GEN_3820 = unuse_way == 2'h1 ? _GEN_746 : _GEN_3436; // @[cache.scala 82:34]
  wire [31:0] _GEN_3821 = unuse_way == 2'h1 ? _GEN_747 : _GEN_3437; // @[cache.scala 82:34]
  wire [31:0] _GEN_3822 = unuse_way == 2'h1 ? _GEN_748 : _GEN_3438; // @[cache.scala 82:34]
  wire [31:0] _GEN_3823 = unuse_way == 2'h1 ? _GEN_749 : _GEN_3439; // @[cache.scala 82:34]
  wire [31:0] _GEN_3824 = unuse_way == 2'h1 ? _GEN_750 : _GEN_3440; // @[cache.scala 82:34]
  wire [31:0] _GEN_3825 = unuse_way == 2'h1 ? _GEN_751 : _GEN_3441; // @[cache.scala 82:34]
  wire [31:0] _GEN_3826 = unuse_way == 2'h1 ? _GEN_752 : _GEN_3442; // @[cache.scala 82:34]
  wire [31:0] _GEN_3827 = unuse_way == 2'h1 ? _GEN_753 : _GEN_3443; // @[cache.scala 82:34]
  wire [31:0] _GEN_3828 = unuse_way == 2'h1 ? _GEN_754 : _GEN_3444; // @[cache.scala 82:34]
  wire [31:0] _GEN_3829 = unuse_way == 2'h1 ? _GEN_755 : _GEN_3445; // @[cache.scala 82:34]
  wire [31:0] _GEN_3830 = unuse_way == 2'h1 ? _GEN_756 : _GEN_3446; // @[cache.scala 82:34]
  wire [31:0] _GEN_3831 = unuse_way == 2'h1 ? _GEN_757 : _GEN_3447; // @[cache.scala 82:34]
  wire [31:0] _GEN_3832 = unuse_way == 2'h1 ? _GEN_758 : _GEN_3448; // @[cache.scala 82:34]
  wire [31:0] _GEN_3833 = unuse_way == 2'h1 ? _GEN_759 : _GEN_3449; // @[cache.scala 82:34]
  wire [31:0] _GEN_3834 = unuse_way == 2'h1 ? _GEN_760 : _GEN_3450; // @[cache.scala 82:34]
  wire [31:0] _GEN_3835 = unuse_way == 2'h1 ? _GEN_761 : _GEN_3451; // @[cache.scala 82:34]
  wire [31:0] _GEN_3836 = unuse_way == 2'h1 ? _GEN_762 : _GEN_3452; // @[cache.scala 82:34]
  wire [31:0] _GEN_3837 = unuse_way == 2'h1 ? _GEN_763 : _GEN_3453; // @[cache.scala 82:34]
  wire [31:0] _GEN_3838 = unuse_way == 2'h1 ? _GEN_764 : _GEN_3454; // @[cache.scala 82:34]
  wire [31:0] _GEN_3839 = unuse_way == 2'h1 ? _GEN_765 : _GEN_3455; // @[cache.scala 82:34]
  wire [31:0] _GEN_3840 = unuse_way == 2'h1 ? _GEN_766 : _GEN_3456; // @[cache.scala 82:34]
  wire [31:0] _GEN_3841 = unuse_way == 2'h1 ? _GEN_767 : _GEN_3457; // @[cache.scala 82:34]
  wire [31:0] _GEN_3842 = unuse_way == 2'h1 ? _GEN_768 : _GEN_3458; // @[cache.scala 82:34]
  wire [31:0] _GEN_3843 = unuse_way == 2'h1 ? _GEN_769 : _GEN_3459; // @[cache.scala 82:34]
  wire [31:0] _GEN_3844 = unuse_way == 2'h1 ? _GEN_770 : _GEN_3460; // @[cache.scala 82:34]
  wire [31:0] _GEN_3845 = unuse_way == 2'h1 ? _GEN_771 : _GEN_3461; // @[cache.scala 82:34]
  wire [31:0] _GEN_3846 = unuse_way == 2'h1 ? _GEN_772 : _GEN_3462; // @[cache.scala 82:34]
  wire [31:0] _GEN_3847 = unuse_way == 2'h1 ? _GEN_773 : _GEN_3463; // @[cache.scala 82:34]
  wire [31:0] _GEN_3848 = unuse_way == 2'h1 ? _GEN_774 : _GEN_3464; // @[cache.scala 82:34]
  wire [31:0] _GEN_3849 = unuse_way == 2'h1 ? _GEN_775 : _GEN_3465; // @[cache.scala 82:34]
  wire [31:0] _GEN_3850 = unuse_way == 2'h1 ? _GEN_776 : _GEN_3466; // @[cache.scala 82:34]
  wire [31:0] _GEN_3851 = unuse_way == 2'h1 ? _GEN_777 : _GEN_3467; // @[cache.scala 82:34]
  wire  _GEN_3852 = unuse_way == 2'h1 ? _GEN_778 : _GEN_3468; // @[cache.scala 82:34]
  wire  _GEN_3853 = unuse_way == 2'h1 ? _GEN_779 : _GEN_3469; // @[cache.scala 82:34]
  wire  _GEN_3854 = unuse_way == 2'h1 ? _GEN_780 : _GEN_3470; // @[cache.scala 82:34]
  wire  _GEN_3855 = unuse_way == 2'h1 ? _GEN_781 : _GEN_3471; // @[cache.scala 82:34]
  wire  _GEN_3856 = unuse_way == 2'h1 ? _GEN_782 : _GEN_3472; // @[cache.scala 82:34]
  wire  _GEN_3857 = unuse_way == 2'h1 ? _GEN_783 : _GEN_3473; // @[cache.scala 82:34]
  wire  _GEN_3858 = unuse_way == 2'h1 ? _GEN_784 : _GEN_3474; // @[cache.scala 82:34]
  wire  _GEN_3859 = unuse_way == 2'h1 ? _GEN_785 : _GEN_3475; // @[cache.scala 82:34]
  wire  _GEN_3860 = unuse_way == 2'h1 ? _GEN_786 : _GEN_3476; // @[cache.scala 82:34]
  wire  _GEN_3861 = unuse_way == 2'h1 ? _GEN_787 : _GEN_3477; // @[cache.scala 82:34]
  wire  _GEN_3862 = unuse_way == 2'h1 ? _GEN_788 : _GEN_3478; // @[cache.scala 82:34]
  wire  _GEN_3863 = unuse_way == 2'h1 ? _GEN_789 : _GEN_3479; // @[cache.scala 82:34]
  wire  _GEN_3864 = unuse_way == 2'h1 ? _GEN_790 : _GEN_3480; // @[cache.scala 82:34]
  wire  _GEN_3865 = unuse_way == 2'h1 ? _GEN_791 : _GEN_3481; // @[cache.scala 82:34]
  wire  _GEN_3866 = unuse_way == 2'h1 ? _GEN_792 : _GEN_3482; // @[cache.scala 82:34]
  wire  _GEN_3867 = unuse_way == 2'h1 ? _GEN_793 : _GEN_3483; // @[cache.scala 82:34]
  wire  _GEN_3868 = unuse_way == 2'h1 ? _GEN_794 : _GEN_3484; // @[cache.scala 82:34]
  wire  _GEN_3869 = unuse_way == 2'h1 ? _GEN_795 : _GEN_3485; // @[cache.scala 82:34]
  wire  _GEN_3870 = unuse_way == 2'h1 ? _GEN_796 : _GEN_3486; // @[cache.scala 82:34]
  wire  _GEN_3871 = unuse_way == 2'h1 ? _GEN_797 : _GEN_3487; // @[cache.scala 82:34]
  wire  _GEN_3872 = unuse_way == 2'h1 ? _GEN_798 : _GEN_3488; // @[cache.scala 82:34]
  wire  _GEN_3873 = unuse_way == 2'h1 ? _GEN_799 : _GEN_3489; // @[cache.scala 82:34]
  wire  _GEN_3874 = unuse_way == 2'h1 ? _GEN_800 : _GEN_3490; // @[cache.scala 82:34]
  wire  _GEN_3875 = unuse_way == 2'h1 ? _GEN_801 : _GEN_3491; // @[cache.scala 82:34]
  wire  _GEN_3876 = unuse_way == 2'h1 ? _GEN_802 : _GEN_3492; // @[cache.scala 82:34]
  wire  _GEN_3877 = unuse_way == 2'h1 ? _GEN_803 : _GEN_3493; // @[cache.scala 82:34]
  wire  _GEN_3878 = unuse_way == 2'h1 ? _GEN_804 : _GEN_3494; // @[cache.scala 82:34]
  wire  _GEN_3879 = unuse_way == 2'h1 ? _GEN_805 : _GEN_3495; // @[cache.scala 82:34]
  wire  _GEN_3880 = unuse_way == 2'h1 ? _GEN_806 : _GEN_3496; // @[cache.scala 82:34]
  wire  _GEN_3881 = unuse_way == 2'h1 ? _GEN_807 : _GEN_3497; // @[cache.scala 82:34]
  wire  _GEN_3882 = unuse_way == 2'h1 ? _GEN_808 : _GEN_3498; // @[cache.scala 82:34]
  wire  _GEN_3883 = unuse_way == 2'h1 ? _GEN_809 : _GEN_3499; // @[cache.scala 82:34]
  wire  _GEN_3884 = unuse_way == 2'h1 ? _GEN_810 : _GEN_3500; // @[cache.scala 82:34]
  wire  _GEN_3885 = unuse_way == 2'h1 ? _GEN_811 : _GEN_3501; // @[cache.scala 82:34]
  wire  _GEN_3886 = unuse_way == 2'h1 ? _GEN_812 : _GEN_3502; // @[cache.scala 82:34]
  wire  _GEN_3887 = unuse_way == 2'h1 ? _GEN_813 : _GEN_3503; // @[cache.scala 82:34]
  wire  _GEN_3888 = unuse_way == 2'h1 ? _GEN_814 : _GEN_3504; // @[cache.scala 82:34]
  wire  _GEN_3889 = unuse_way == 2'h1 ? _GEN_815 : _GEN_3505; // @[cache.scala 82:34]
  wire  _GEN_3890 = unuse_way == 2'h1 ? _GEN_816 : _GEN_3506; // @[cache.scala 82:34]
  wire  _GEN_3891 = unuse_way == 2'h1 ? _GEN_817 : _GEN_3507; // @[cache.scala 82:34]
  wire  _GEN_3892 = unuse_way == 2'h1 ? _GEN_818 : _GEN_3508; // @[cache.scala 82:34]
  wire  _GEN_3893 = unuse_way == 2'h1 ? _GEN_819 : _GEN_3509; // @[cache.scala 82:34]
  wire  _GEN_3894 = unuse_way == 2'h1 ? _GEN_820 : _GEN_3510; // @[cache.scala 82:34]
  wire  _GEN_3895 = unuse_way == 2'h1 ? _GEN_821 : _GEN_3511; // @[cache.scala 82:34]
  wire  _GEN_3896 = unuse_way == 2'h1 ? _GEN_822 : _GEN_3512; // @[cache.scala 82:34]
  wire  _GEN_3897 = unuse_way == 2'h1 ? _GEN_823 : _GEN_3513; // @[cache.scala 82:34]
  wire  _GEN_3898 = unuse_way == 2'h1 ? _GEN_824 : _GEN_3514; // @[cache.scala 82:34]
  wire  _GEN_3899 = unuse_way == 2'h1 ? _GEN_825 : _GEN_3515; // @[cache.scala 82:34]
  wire  _GEN_3900 = unuse_way == 2'h1 ? _GEN_826 : _GEN_3516; // @[cache.scala 82:34]
  wire  _GEN_3901 = unuse_way == 2'h1 ? _GEN_827 : _GEN_3517; // @[cache.scala 82:34]
  wire  _GEN_3902 = unuse_way == 2'h1 ? _GEN_828 : _GEN_3518; // @[cache.scala 82:34]
  wire  _GEN_3903 = unuse_way == 2'h1 ? _GEN_829 : _GEN_3519; // @[cache.scala 82:34]
  wire  _GEN_3904 = unuse_way == 2'h1 ? _GEN_830 : _GEN_3520; // @[cache.scala 82:34]
  wire  _GEN_3905 = unuse_way == 2'h1 ? _GEN_831 : _GEN_3521; // @[cache.scala 82:34]
  wire  _GEN_3906 = unuse_way == 2'h1 ? _GEN_832 : _GEN_3522; // @[cache.scala 82:34]
  wire  _GEN_3907 = unuse_way == 2'h1 ? _GEN_833 : _GEN_3523; // @[cache.scala 82:34]
  wire  _GEN_3908 = unuse_way == 2'h1 ? _GEN_834 : _GEN_3524; // @[cache.scala 82:34]
  wire  _GEN_3909 = unuse_way == 2'h1 ? _GEN_835 : _GEN_3525; // @[cache.scala 82:34]
  wire  _GEN_3910 = unuse_way == 2'h1 ? _GEN_836 : _GEN_3526; // @[cache.scala 82:34]
  wire  _GEN_3911 = unuse_way == 2'h1 ? _GEN_837 : _GEN_3527; // @[cache.scala 82:34]
  wire  _GEN_3912 = unuse_way == 2'h1 ? _GEN_838 : _GEN_3528; // @[cache.scala 82:34]
  wire  _GEN_3913 = unuse_way == 2'h1 ? _GEN_839 : _GEN_3529; // @[cache.scala 82:34]
  wire  _GEN_3914 = unuse_way == 2'h1 ? _GEN_840 : _GEN_3530; // @[cache.scala 82:34]
  wire  _GEN_3915 = unuse_way == 2'h1 ? _GEN_841 : _GEN_3531; // @[cache.scala 82:34]
  wire  _GEN_3916 = unuse_way == 2'h1 ? _GEN_842 : _GEN_3532; // @[cache.scala 82:34]
  wire  _GEN_3917 = unuse_way == 2'h1 ? _GEN_843 : _GEN_3533; // @[cache.scala 82:34]
  wire  _GEN_3918 = unuse_way == 2'h1 ? _GEN_844 : _GEN_3534; // @[cache.scala 82:34]
  wire  _GEN_3919 = unuse_way == 2'h1 ? _GEN_845 : _GEN_3535; // @[cache.scala 82:34]
  wire  _GEN_3920 = unuse_way == 2'h1 ? _GEN_846 : _GEN_3536; // @[cache.scala 82:34]
  wire  _GEN_3921 = unuse_way == 2'h1 ? _GEN_847 : _GEN_3537; // @[cache.scala 82:34]
  wire  _GEN_3922 = unuse_way == 2'h1 ? _GEN_848 : _GEN_3538; // @[cache.scala 82:34]
  wire  _GEN_3923 = unuse_way == 2'h1 ? _GEN_849 : _GEN_3539; // @[cache.scala 82:34]
  wire  _GEN_3924 = unuse_way == 2'h1 ? _GEN_850 : _GEN_3540; // @[cache.scala 82:34]
  wire  _GEN_3925 = unuse_way == 2'h1 ? _GEN_851 : _GEN_3541; // @[cache.scala 82:34]
  wire  _GEN_3926 = unuse_way == 2'h1 ? _GEN_852 : _GEN_3542; // @[cache.scala 82:34]
  wire  _GEN_3927 = unuse_way == 2'h1 ? _GEN_853 : _GEN_3543; // @[cache.scala 82:34]
  wire  _GEN_3928 = unuse_way == 2'h1 ? _GEN_854 : _GEN_3544; // @[cache.scala 82:34]
  wire  _GEN_3929 = unuse_way == 2'h1 ? _GEN_855 : _GEN_3545; // @[cache.scala 82:34]
  wire  _GEN_3930 = unuse_way == 2'h1 ? _GEN_856 : _GEN_3546; // @[cache.scala 82:34]
  wire  _GEN_3931 = unuse_way == 2'h1 ? _GEN_857 : _GEN_3547; // @[cache.scala 82:34]
  wire  _GEN_3932 = unuse_way == 2'h1 ? _GEN_858 : _GEN_3548; // @[cache.scala 82:34]
  wire  _GEN_3933 = unuse_way == 2'h1 ? _GEN_859 : _GEN_3549; // @[cache.scala 82:34]
  wire  _GEN_3934 = unuse_way == 2'h1 ? _GEN_860 : _GEN_3550; // @[cache.scala 82:34]
  wire  _GEN_3935 = unuse_way == 2'h1 ? _GEN_861 : _GEN_3551; // @[cache.scala 82:34]
  wire  _GEN_3936 = unuse_way == 2'h1 ? _GEN_862 : _GEN_3552; // @[cache.scala 82:34]
  wire  _GEN_3937 = unuse_way == 2'h1 ? _GEN_863 : _GEN_3553; // @[cache.scala 82:34]
  wire  _GEN_3938 = unuse_way == 2'h1 ? _GEN_864 : _GEN_3554; // @[cache.scala 82:34]
  wire  _GEN_3939 = unuse_way == 2'h1 ? _GEN_865 : _GEN_3555; // @[cache.scala 82:34]
  wire  _GEN_3940 = unuse_way == 2'h1 ? _GEN_866 : _GEN_3556; // @[cache.scala 82:34]
  wire  _GEN_3941 = unuse_way == 2'h1 ? _GEN_867 : _GEN_3557; // @[cache.scala 82:34]
  wire  _GEN_3942 = unuse_way == 2'h1 ? _GEN_868 : _GEN_3558; // @[cache.scala 82:34]
  wire  _GEN_3943 = unuse_way == 2'h1 ? _GEN_869 : _GEN_3559; // @[cache.scala 82:34]
  wire  _GEN_3944 = unuse_way == 2'h1 ? _GEN_870 : _GEN_3560; // @[cache.scala 82:34]
  wire  _GEN_3945 = unuse_way == 2'h1 ? _GEN_871 : _GEN_3561; // @[cache.scala 82:34]
  wire  _GEN_3946 = unuse_way == 2'h1 ? _GEN_872 : _GEN_3562; // @[cache.scala 82:34]
  wire  _GEN_3947 = unuse_way == 2'h1 ? _GEN_873 : _GEN_3563; // @[cache.scala 82:34]
  wire  _GEN_3948 = unuse_way == 2'h1 ? _GEN_874 : _GEN_3564; // @[cache.scala 82:34]
  wire  _GEN_3949 = unuse_way == 2'h1 ? _GEN_875 : _GEN_3565; // @[cache.scala 82:34]
  wire  _GEN_3950 = unuse_way == 2'h1 ? _GEN_876 : _GEN_3566; // @[cache.scala 82:34]
  wire  _GEN_3951 = unuse_way == 2'h1 ? _GEN_877 : _GEN_3567; // @[cache.scala 82:34]
  wire  _GEN_3952 = unuse_way == 2'h1 ? _GEN_878 : _GEN_3568; // @[cache.scala 82:34]
  wire  _GEN_3953 = unuse_way == 2'h1 ? _GEN_879 : _GEN_3569; // @[cache.scala 82:34]
  wire  _GEN_3954 = unuse_way == 2'h1 ? _GEN_880 : _GEN_3570; // @[cache.scala 82:34]
  wire  _GEN_3955 = unuse_way == 2'h1 ? _GEN_881 : _GEN_3571; // @[cache.scala 82:34]
  wire  _GEN_3956 = unuse_way == 2'h1 ? _GEN_882 : _GEN_3572; // @[cache.scala 82:34]
  wire  _GEN_3957 = unuse_way == 2'h1 ? _GEN_883 : _GEN_3573; // @[cache.scala 82:34]
  wire  _GEN_3958 = unuse_way == 2'h1 ? _GEN_884 : _GEN_3574; // @[cache.scala 82:34]
  wire  _GEN_3959 = unuse_way == 2'h1 ? _GEN_885 : _GEN_3575; // @[cache.scala 82:34]
  wire  _GEN_3960 = unuse_way == 2'h1 ? _GEN_886 : _GEN_3576; // @[cache.scala 82:34]
  wire  _GEN_3961 = unuse_way == 2'h1 ? _GEN_887 : _GEN_3577; // @[cache.scala 82:34]
  wire  _GEN_3962 = unuse_way == 2'h1 ? _GEN_888 : _GEN_3578; // @[cache.scala 82:34]
  wire  _GEN_3963 = unuse_way == 2'h1 ? _GEN_889 : _GEN_3579; // @[cache.scala 82:34]
  wire  _GEN_3964 = unuse_way == 2'h1 ? _GEN_890 : _GEN_3580; // @[cache.scala 82:34]
  wire  _GEN_3965 = unuse_way == 2'h1 ? _GEN_891 : _GEN_3581; // @[cache.scala 82:34]
  wire  _GEN_3966 = unuse_way == 2'h1 ? _GEN_892 : _GEN_3582; // @[cache.scala 82:34]
  wire  _GEN_3967 = unuse_way == 2'h1 ? _GEN_893 : _GEN_3583; // @[cache.scala 82:34]
  wire  _GEN_3968 = unuse_way == 2'h1 ? _GEN_894 : _GEN_3584; // @[cache.scala 82:34]
  wire  _GEN_3969 = unuse_way == 2'h1 ? _GEN_895 : _GEN_3585; // @[cache.scala 82:34]
  wire  _GEN_3970 = unuse_way == 2'h1 ? _GEN_896 : _GEN_3586; // @[cache.scala 82:34]
  wire  _GEN_3971 = unuse_way == 2'h1 ? _GEN_897 : _GEN_3587; // @[cache.scala 82:34]
  wire  _GEN_3972 = unuse_way == 2'h1 ? _GEN_898 : _GEN_3588; // @[cache.scala 82:34]
  wire  _GEN_3973 = unuse_way == 2'h1 ? _GEN_899 : _GEN_3589; // @[cache.scala 82:34]
  wire  _GEN_3974 = unuse_way == 2'h1 ? _GEN_900 : _GEN_3590; // @[cache.scala 82:34]
  wire  _GEN_3975 = unuse_way == 2'h1 ? _GEN_901 : _GEN_3591; // @[cache.scala 82:34]
  wire  _GEN_3976 = unuse_way == 2'h1 ? _GEN_902 : _GEN_3592; // @[cache.scala 82:34]
  wire  _GEN_3977 = unuse_way == 2'h1 ? _GEN_903 : _GEN_3593; // @[cache.scala 82:34]
  wire  _GEN_3978 = unuse_way == 2'h1 ? _GEN_904 : _GEN_3594; // @[cache.scala 82:34]
  wire  _GEN_3979 = unuse_way == 2'h1 ? _GEN_905 : _GEN_3595; // @[cache.scala 82:34]
  wire  _GEN_3980 = unuse_way == 2'h1 | _GEN_3211; // @[cache.scala 82:34 86:23]
  wire [63:0] _GEN_3981 = unuse_way == 2'h1 ? ram_1_0 : _GEN_2827; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3982 = unuse_way == 2'h1 ? ram_1_1 : _GEN_2828; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3983 = unuse_way == 2'h1 ? ram_1_2 : _GEN_2829; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3984 = unuse_way == 2'h1 ? ram_1_3 : _GEN_2830; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3985 = unuse_way == 2'h1 ? ram_1_4 : _GEN_2831; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3986 = unuse_way == 2'h1 ? ram_1_5 : _GEN_2832; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3987 = unuse_way == 2'h1 ? ram_1_6 : _GEN_2833; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3988 = unuse_way == 2'h1 ? ram_1_7 : _GEN_2834; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3989 = unuse_way == 2'h1 ? ram_1_8 : _GEN_2835; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3990 = unuse_way == 2'h1 ? ram_1_9 : _GEN_2836; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3991 = unuse_way == 2'h1 ? ram_1_10 : _GEN_2837; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3992 = unuse_way == 2'h1 ? ram_1_11 : _GEN_2838; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3993 = unuse_way == 2'h1 ? ram_1_12 : _GEN_2839; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3994 = unuse_way == 2'h1 ? ram_1_13 : _GEN_2840; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3995 = unuse_way == 2'h1 ? ram_1_14 : _GEN_2841; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3996 = unuse_way == 2'h1 ? ram_1_15 : _GEN_2842; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3997 = unuse_way == 2'h1 ? ram_1_16 : _GEN_2843; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3998 = unuse_way == 2'h1 ? ram_1_17 : _GEN_2844; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_3999 = unuse_way == 2'h1 ? ram_1_18 : _GEN_2845; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4000 = unuse_way == 2'h1 ? ram_1_19 : _GEN_2846; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4001 = unuse_way == 2'h1 ? ram_1_20 : _GEN_2847; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4002 = unuse_way == 2'h1 ? ram_1_21 : _GEN_2848; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4003 = unuse_way == 2'h1 ? ram_1_22 : _GEN_2849; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4004 = unuse_way == 2'h1 ? ram_1_23 : _GEN_2850; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4005 = unuse_way == 2'h1 ? ram_1_24 : _GEN_2851; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4006 = unuse_way == 2'h1 ? ram_1_25 : _GEN_2852; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4007 = unuse_way == 2'h1 ? ram_1_26 : _GEN_2853; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4008 = unuse_way == 2'h1 ? ram_1_27 : _GEN_2854; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4009 = unuse_way == 2'h1 ? ram_1_28 : _GEN_2855; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4010 = unuse_way == 2'h1 ? ram_1_29 : _GEN_2856; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4011 = unuse_way == 2'h1 ? ram_1_30 : _GEN_2857; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4012 = unuse_way == 2'h1 ? ram_1_31 : _GEN_2858; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4013 = unuse_way == 2'h1 ? ram_1_32 : _GEN_2859; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4014 = unuse_way == 2'h1 ? ram_1_33 : _GEN_2860; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4015 = unuse_way == 2'h1 ? ram_1_34 : _GEN_2861; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4016 = unuse_way == 2'h1 ? ram_1_35 : _GEN_2862; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4017 = unuse_way == 2'h1 ? ram_1_36 : _GEN_2863; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4018 = unuse_way == 2'h1 ? ram_1_37 : _GEN_2864; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4019 = unuse_way == 2'h1 ? ram_1_38 : _GEN_2865; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4020 = unuse_way == 2'h1 ? ram_1_39 : _GEN_2866; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4021 = unuse_way == 2'h1 ? ram_1_40 : _GEN_2867; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4022 = unuse_way == 2'h1 ? ram_1_41 : _GEN_2868; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4023 = unuse_way == 2'h1 ? ram_1_42 : _GEN_2869; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4024 = unuse_way == 2'h1 ? ram_1_43 : _GEN_2870; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4025 = unuse_way == 2'h1 ? ram_1_44 : _GEN_2871; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4026 = unuse_way == 2'h1 ? ram_1_45 : _GEN_2872; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4027 = unuse_way == 2'h1 ? ram_1_46 : _GEN_2873; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4028 = unuse_way == 2'h1 ? ram_1_47 : _GEN_2874; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4029 = unuse_way == 2'h1 ? ram_1_48 : _GEN_2875; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4030 = unuse_way == 2'h1 ? ram_1_49 : _GEN_2876; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4031 = unuse_way == 2'h1 ? ram_1_50 : _GEN_2877; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4032 = unuse_way == 2'h1 ? ram_1_51 : _GEN_2878; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4033 = unuse_way == 2'h1 ? ram_1_52 : _GEN_2879; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4034 = unuse_way == 2'h1 ? ram_1_53 : _GEN_2880; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4035 = unuse_way == 2'h1 ? ram_1_54 : _GEN_2881; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4036 = unuse_way == 2'h1 ? ram_1_55 : _GEN_2882; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4037 = unuse_way == 2'h1 ? ram_1_56 : _GEN_2883; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4038 = unuse_way == 2'h1 ? ram_1_57 : _GEN_2884; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4039 = unuse_way == 2'h1 ? ram_1_58 : _GEN_2885; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4040 = unuse_way == 2'h1 ? ram_1_59 : _GEN_2886; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4041 = unuse_way == 2'h1 ? ram_1_60 : _GEN_2887; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4042 = unuse_way == 2'h1 ? ram_1_61 : _GEN_2888; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4043 = unuse_way == 2'h1 ? ram_1_62 : _GEN_2889; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4044 = unuse_way == 2'h1 ? ram_1_63 : _GEN_2890; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4045 = unuse_way == 2'h1 ? ram_1_64 : _GEN_2891; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4046 = unuse_way == 2'h1 ? ram_1_65 : _GEN_2892; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4047 = unuse_way == 2'h1 ? ram_1_66 : _GEN_2893; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4048 = unuse_way == 2'h1 ? ram_1_67 : _GEN_2894; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4049 = unuse_way == 2'h1 ? ram_1_68 : _GEN_2895; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4050 = unuse_way == 2'h1 ? ram_1_69 : _GEN_2896; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4051 = unuse_way == 2'h1 ? ram_1_70 : _GEN_2897; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4052 = unuse_way == 2'h1 ? ram_1_71 : _GEN_2898; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4053 = unuse_way == 2'h1 ? ram_1_72 : _GEN_2899; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4054 = unuse_way == 2'h1 ? ram_1_73 : _GEN_2900; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4055 = unuse_way == 2'h1 ? ram_1_74 : _GEN_2901; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4056 = unuse_way == 2'h1 ? ram_1_75 : _GEN_2902; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4057 = unuse_way == 2'h1 ? ram_1_76 : _GEN_2903; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4058 = unuse_way == 2'h1 ? ram_1_77 : _GEN_2904; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4059 = unuse_way == 2'h1 ? ram_1_78 : _GEN_2905; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4060 = unuse_way == 2'h1 ? ram_1_79 : _GEN_2906; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4061 = unuse_way == 2'h1 ? ram_1_80 : _GEN_2907; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4062 = unuse_way == 2'h1 ? ram_1_81 : _GEN_2908; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4063 = unuse_way == 2'h1 ? ram_1_82 : _GEN_2909; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4064 = unuse_way == 2'h1 ? ram_1_83 : _GEN_2910; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4065 = unuse_way == 2'h1 ? ram_1_84 : _GEN_2911; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4066 = unuse_way == 2'h1 ? ram_1_85 : _GEN_2912; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4067 = unuse_way == 2'h1 ? ram_1_86 : _GEN_2913; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4068 = unuse_way == 2'h1 ? ram_1_87 : _GEN_2914; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4069 = unuse_way == 2'h1 ? ram_1_88 : _GEN_2915; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4070 = unuse_way == 2'h1 ? ram_1_89 : _GEN_2916; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4071 = unuse_way == 2'h1 ? ram_1_90 : _GEN_2917; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4072 = unuse_way == 2'h1 ? ram_1_91 : _GEN_2918; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4073 = unuse_way == 2'h1 ? ram_1_92 : _GEN_2919; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4074 = unuse_way == 2'h1 ? ram_1_93 : _GEN_2920; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4075 = unuse_way == 2'h1 ? ram_1_94 : _GEN_2921; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4076 = unuse_way == 2'h1 ? ram_1_95 : _GEN_2922; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4077 = unuse_way == 2'h1 ? ram_1_96 : _GEN_2923; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4078 = unuse_way == 2'h1 ? ram_1_97 : _GEN_2924; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4079 = unuse_way == 2'h1 ? ram_1_98 : _GEN_2925; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4080 = unuse_way == 2'h1 ? ram_1_99 : _GEN_2926; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4081 = unuse_way == 2'h1 ? ram_1_100 : _GEN_2927; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4082 = unuse_way == 2'h1 ? ram_1_101 : _GEN_2928; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4083 = unuse_way == 2'h1 ? ram_1_102 : _GEN_2929; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4084 = unuse_way == 2'h1 ? ram_1_103 : _GEN_2930; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4085 = unuse_way == 2'h1 ? ram_1_104 : _GEN_2931; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4086 = unuse_way == 2'h1 ? ram_1_105 : _GEN_2932; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4087 = unuse_way == 2'h1 ? ram_1_106 : _GEN_2933; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4088 = unuse_way == 2'h1 ? ram_1_107 : _GEN_2934; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4089 = unuse_way == 2'h1 ? ram_1_108 : _GEN_2935; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4090 = unuse_way == 2'h1 ? ram_1_109 : _GEN_2936; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4091 = unuse_way == 2'h1 ? ram_1_110 : _GEN_2937; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4092 = unuse_way == 2'h1 ? ram_1_111 : _GEN_2938; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4093 = unuse_way == 2'h1 ? ram_1_112 : _GEN_2939; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4094 = unuse_way == 2'h1 ? ram_1_113 : _GEN_2940; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4095 = unuse_way == 2'h1 ? ram_1_114 : _GEN_2941; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4096 = unuse_way == 2'h1 ? ram_1_115 : _GEN_2942; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4097 = unuse_way == 2'h1 ? ram_1_116 : _GEN_2943; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4098 = unuse_way == 2'h1 ? ram_1_117 : _GEN_2944; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4099 = unuse_way == 2'h1 ? ram_1_118 : _GEN_2945; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4100 = unuse_way == 2'h1 ? ram_1_119 : _GEN_2946; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4101 = unuse_way == 2'h1 ? ram_1_120 : _GEN_2947; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4102 = unuse_way == 2'h1 ? ram_1_121 : _GEN_2948; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4103 = unuse_way == 2'h1 ? ram_1_122 : _GEN_2949; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4104 = unuse_way == 2'h1 ? ram_1_123 : _GEN_2950; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4105 = unuse_way == 2'h1 ? ram_1_124 : _GEN_2951; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4106 = unuse_way == 2'h1 ? ram_1_125 : _GEN_2952; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4107 = unuse_way == 2'h1 ? ram_1_126 : _GEN_2953; // @[cache.scala 18:24 82:34]
  wire [63:0] _GEN_4108 = unuse_way == 2'h1 ? ram_1_127 : _GEN_2954; // @[cache.scala 18:24 82:34]
  wire [31:0] _GEN_4109 = unuse_way == 2'h1 ? tag_1_0 : _GEN_2955; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4110 = unuse_way == 2'h1 ? tag_1_1 : _GEN_2956; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4111 = unuse_way == 2'h1 ? tag_1_2 : _GEN_2957; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4112 = unuse_way == 2'h1 ? tag_1_3 : _GEN_2958; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4113 = unuse_way == 2'h1 ? tag_1_4 : _GEN_2959; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4114 = unuse_way == 2'h1 ? tag_1_5 : _GEN_2960; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4115 = unuse_way == 2'h1 ? tag_1_6 : _GEN_2961; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4116 = unuse_way == 2'h1 ? tag_1_7 : _GEN_2962; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4117 = unuse_way == 2'h1 ? tag_1_8 : _GEN_2963; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4118 = unuse_way == 2'h1 ? tag_1_9 : _GEN_2964; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4119 = unuse_way == 2'h1 ? tag_1_10 : _GEN_2965; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4120 = unuse_way == 2'h1 ? tag_1_11 : _GEN_2966; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4121 = unuse_way == 2'h1 ? tag_1_12 : _GEN_2967; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4122 = unuse_way == 2'h1 ? tag_1_13 : _GEN_2968; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4123 = unuse_way == 2'h1 ? tag_1_14 : _GEN_2969; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4124 = unuse_way == 2'h1 ? tag_1_15 : _GEN_2970; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4125 = unuse_way == 2'h1 ? tag_1_16 : _GEN_2971; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4126 = unuse_way == 2'h1 ? tag_1_17 : _GEN_2972; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4127 = unuse_way == 2'h1 ? tag_1_18 : _GEN_2973; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4128 = unuse_way == 2'h1 ? tag_1_19 : _GEN_2974; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4129 = unuse_way == 2'h1 ? tag_1_20 : _GEN_2975; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4130 = unuse_way == 2'h1 ? tag_1_21 : _GEN_2976; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4131 = unuse_way == 2'h1 ? tag_1_22 : _GEN_2977; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4132 = unuse_way == 2'h1 ? tag_1_23 : _GEN_2978; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4133 = unuse_way == 2'h1 ? tag_1_24 : _GEN_2979; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4134 = unuse_way == 2'h1 ? tag_1_25 : _GEN_2980; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4135 = unuse_way == 2'h1 ? tag_1_26 : _GEN_2981; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4136 = unuse_way == 2'h1 ? tag_1_27 : _GEN_2982; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4137 = unuse_way == 2'h1 ? tag_1_28 : _GEN_2983; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4138 = unuse_way == 2'h1 ? tag_1_29 : _GEN_2984; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4139 = unuse_way == 2'h1 ? tag_1_30 : _GEN_2985; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4140 = unuse_way == 2'h1 ? tag_1_31 : _GEN_2986; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4141 = unuse_way == 2'h1 ? tag_1_32 : _GEN_2987; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4142 = unuse_way == 2'h1 ? tag_1_33 : _GEN_2988; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4143 = unuse_way == 2'h1 ? tag_1_34 : _GEN_2989; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4144 = unuse_way == 2'h1 ? tag_1_35 : _GEN_2990; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4145 = unuse_way == 2'h1 ? tag_1_36 : _GEN_2991; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4146 = unuse_way == 2'h1 ? tag_1_37 : _GEN_2992; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4147 = unuse_way == 2'h1 ? tag_1_38 : _GEN_2993; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4148 = unuse_way == 2'h1 ? tag_1_39 : _GEN_2994; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4149 = unuse_way == 2'h1 ? tag_1_40 : _GEN_2995; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4150 = unuse_way == 2'h1 ? tag_1_41 : _GEN_2996; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4151 = unuse_way == 2'h1 ? tag_1_42 : _GEN_2997; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4152 = unuse_way == 2'h1 ? tag_1_43 : _GEN_2998; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4153 = unuse_way == 2'h1 ? tag_1_44 : _GEN_2999; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4154 = unuse_way == 2'h1 ? tag_1_45 : _GEN_3000; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4155 = unuse_way == 2'h1 ? tag_1_46 : _GEN_3001; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4156 = unuse_way == 2'h1 ? tag_1_47 : _GEN_3002; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4157 = unuse_way == 2'h1 ? tag_1_48 : _GEN_3003; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4158 = unuse_way == 2'h1 ? tag_1_49 : _GEN_3004; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4159 = unuse_way == 2'h1 ? tag_1_50 : _GEN_3005; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4160 = unuse_way == 2'h1 ? tag_1_51 : _GEN_3006; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4161 = unuse_way == 2'h1 ? tag_1_52 : _GEN_3007; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4162 = unuse_way == 2'h1 ? tag_1_53 : _GEN_3008; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4163 = unuse_way == 2'h1 ? tag_1_54 : _GEN_3009; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4164 = unuse_way == 2'h1 ? tag_1_55 : _GEN_3010; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4165 = unuse_way == 2'h1 ? tag_1_56 : _GEN_3011; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4166 = unuse_way == 2'h1 ? tag_1_57 : _GEN_3012; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4167 = unuse_way == 2'h1 ? tag_1_58 : _GEN_3013; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4168 = unuse_way == 2'h1 ? tag_1_59 : _GEN_3014; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4169 = unuse_way == 2'h1 ? tag_1_60 : _GEN_3015; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4170 = unuse_way == 2'h1 ? tag_1_61 : _GEN_3016; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4171 = unuse_way == 2'h1 ? tag_1_62 : _GEN_3017; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4172 = unuse_way == 2'h1 ? tag_1_63 : _GEN_3018; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4173 = unuse_way == 2'h1 ? tag_1_64 : _GEN_3019; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4174 = unuse_way == 2'h1 ? tag_1_65 : _GEN_3020; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4175 = unuse_way == 2'h1 ? tag_1_66 : _GEN_3021; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4176 = unuse_way == 2'h1 ? tag_1_67 : _GEN_3022; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4177 = unuse_way == 2'h1 ? tag_1_68 : _GEN_3023; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4178 = unuse_way == 2'h1 ? tag_1_69 : _GEN_3024; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4179 = unuse_way == 2'h1 ? tag_1_70 : _GEN_3025; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4180 = unuse_way == 2'h1 ? tag_1_71 : _GEN_3026; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4181 = unuse_way == 2'h1 ? tag_1_72 : _GEN_3027; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4182 = unuse_way == 2'h1 ? tag_1_73 : _GEN_3028; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4183 = unuse_way == 2'h1 ? tag_1_74 : _GEN_3029; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4184 = unuse_way == 2'h1 ? tag_1_75 : _GEN_3030; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4185 = unuse_way == 2'h1 ? tag_1_76 : _GEN_3031; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4186 = unuse_way == 2'h1 ? tag_1_77 : _GEN_3032; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4187 = unuse_way == 2'h1 ? tag_1_78 : _GEN_3033; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4188 = unuse_way == 2'h1 ? tag_1_79 : _GEN_3034; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4189 = unuse_way == 2'h1 ? tag_1_80 : _GEN_3035; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4190 = unuse_way == 2'h1 ? tag_1_81 : _GEN_3036; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4191 = unuse_way == 2'h1 ? tag_1_82 : _GEN_3037; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4192 = unuse_way == 2'h1 ? tag_1_83 : _GEN_3038; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4193 = unuse_way == 2'h1 ? tag_1_84 : _GEN_3039; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4194 = unuse_way == 2'h1 ? tag_1_85 : _GEN_3040; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4195 = unuse_way == 2'h1 ? tag_1_86 : _GEN_3041; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4196 = unuse_way == 2'h1 ? tag_1_87 : _GEN_3042; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4197 = unuse_way == 2'h1 ? tag_1_88 : _GEN_3043; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4198 = unuse_way == 2'h1 ? tag_1_89 : _GEN_3044; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4199 = unuse_way == 2'h1 ? tag_1_90 : _GEN_3045; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4200 = unuse_way == 2'h1 ? tag_1_91 : _GEN_3046; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4201 = unuse_way == 2'h1 ? tag_1_92 : _GEN_3047; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4202 = unuse_way == 2'h1 ? tag_1_93 : _GEN_3048; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4203 = unuse_way == 2'h1 ? tag_1_94 : _GEN_3049; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4204 = unuse_way == 2'h1 ? tag_1_95 : _GEN_3050; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4205 = unuse_way == 2'h1 ? tag_1_96 : _GEN_3051; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4206 = unuse_way == 2'h1 ? tag_1_97 : _GEN_3052; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4207 = unuse_way == 2'h1 ? tag_1_98 : _GEN_3053; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4208 = unuse_way == 2'h1 ? tag_1_99 : _GEN_3054; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4209 = unuse_way == 2'h1 ? tag_1_100 : _GEN_3055; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4210 = unuse_way == 2'h1 ? tag_1_101 : _GEN_3056; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4211 = unuse_way == 2'h1 ? tag_1_102 : _GEN_3057; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4212 = unuse_way == 2'h1 ? tag_1_103 : _GEN_3058; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4213 = unuse_way == 2'h1 ? tag_1_104 : _GEN_3059; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4214 = unuse_way == 2'h1 ? tag_1_105 : _GEN_3060; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4215 = unuse_way == 2'h1 ? tag_1_106 : _GEN_3061; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4216 = unuse_way == 2'h1 ? tag_1_107 : _GEN_3062; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4217 = unuse_way == 2'h1 ? tag_1_108 : _GEN_3063; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4218 = unuse_way == 2'h1 ? tag_1_109 : _GEN_3064; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4219 = unuse_way == 2'h1 ? tag_1_110 : _GEN_3065; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4220 = unuse_way == 2'h1 ? tag_1_111 : _GEN_3066; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4221 = unuse_way == 2'h1 ? tag_1_112 : _GEN_3067; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4222 = unuse_way == 2'h1 ? tag_1_113 : _GEN_3068; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4223 = unuse_way == 2'h1 ? tag_1_114 : _GEN_3069; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4224 = unuse_way == 2'h1 ? tag_1_115 : _GEN_3070; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4225 = unuse_way == 2'h1 ? tag_1_116 : _GEN_3071; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4226 = unuse_way == 2'h1 ? tag_1_117 : _GEN_3072; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4227 = unuse_way == 2'h1 ? tag_1_118 : _GEN_3073; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4228 = unuse_way == 2'h1 ? tag_1_119 : _GEN_3074; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4229 = unuse_way == 2'h1 ? tag_1_120 : _GEN_3075; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4230 = unuse_way == 2'h1 ? tag_1_121 : _GEN_3076; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4231 = unuse_way == 2'h1 ? tag_1_122 : _GEN_3077; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4232 = unuse_way == 2'h1 ? tag_1_123 : _GEN_3078; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4233 = unuse_way == 2'h1 ? tag_1_124 : _GEN_3079; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4234 = unuse_way == 2'h1 ? tag_1_125 : _GEN_3080; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4235 = unuse_way == 2'h1 ? tag_1_126 : _GEN_3081; // @[cache.scala 20:24 82:34]
  wire [31:0] _GEN_4236 = unuse_way == 2'h1 ? tag_1_127 : _GEN_3082; // @[cache.scala 20:24 82:34]
  wire  _GEN_4237 = unuse_way == 2'h1 ? valid_1_0 : _GEN_3083; // @[cache.scala 22:26 82:34]
  wire  _GEN_4238 = unuse_way == 2'h1 ? valid_1_1 : _GEN_3084; // @[cache.scala 22:26 82:34]
  wire  _GEN_4239 = unuse_way == 2'h1 ? valid_1_2 : _GEN_3085; // @[cache.scala 22:26 82:34]
  wire  _GEN_4240 = unuse_way == 2'h1 ? valid_1_3 : _GEN_3086; // @[cache.scala 22:26 82:34]
  wire  _GEN_4241 = unuse_way == 2'h1 ? valid_1_4 : _GEN_3087; // @[cache.scala 22:26 82:34]
  wire  _GEN_4242 = unuse_way == 2'h1 ? valid_1_5 : _GEN_3088; // @[cache.scala 22:26 82:34]
  wire  _GEN_4243 = unuse_way == 2'h1 ? valid_1_6 : _GEN_3089; // @[cache.scala 22:26 82:34]
  wire  _GEN_4244 = unuse_way == 2'h1 ? valid_1_7 : _GEN_3090; // @[cache.scala 22:26 82:34]
  wire  _GEN_4245 = unuse_way == 2'h1 ? valid_1_8 : _GEN_3091; // @[cache.scala 22:26 82:34]
  wire  _GEN_4246 = unuse_way == 2'h1 ? valid_1_9 : _GEN_3092; // @[cache.scala 22:26 82:34]
  wire  _GEN_4247 = unuse_way == 2'h1 ? valid_1_10 : _GEN_3093; // @[cache.scala 22:26 82:34]
  wire  _GEN_4248 = unuse_way == 2'h1 ? valid_1_11 : _GEN_3094; // @[cache.scala 22:26 82:34]
  wire  _GEN_4249 = unuse_way == 2'h1 ? valid_1_12 : _GEN_3095; // @[cache.scala 22:26 82:34]
  wire  _GEN_4250 = unuse_way == 2'h1 ? valid_1_13 : _GEN_3096; // @[cache.scala 22:26 82:34]
  wire  _GEN_4251 = unuse_way == 2'h1 ? valid_1_14 : _GEN_3097; // @[cache.scala 22:26 82:34]
  wire  _GEN_4252 = unuse_way == 2'h1 ? valid_1_15 : _GEN_3098; // @[cache.scala 22:26 82:34]
  wire  _GEN_4253 = unuse_way == 2'h1 ? valid_1_16 : _GEN_3099; // @[cache.scala 22:26 82:34]
  wire  _GEN_4254 = unuse_way == 2'h1 ? valid_1_17 : _GEN_3100; // @[cache.scala 22:26 82:34]
  wire  _GEN_4255 = unuse_way == 2'h1 ? valid_1_18 : _GEN_3101; // @[cache.scala 22:26 82:34]
  wire  _GEN_4256 = unuse_way == 2'h1 ? valid_1_19 : _GEN_3102; // @[cache.scala 22:26 82:34]
  wire  _GEN_4257 = unuse_way == 2'h1 ? valid_1_20 : _GEN_3103; // @[cache.scala 22:26 82:34]
  wire  _GEN_4258 = unuse_way == 2'h1 ? valid_1_21 : _GEN_3104; // @[cache.scala 22:26 82:34]
  wire  _GEN_4259 = unuse_way == 2'h1 ? valid_1_22 : _GEN_3105; // @[cache.scala 22:26 82:34]
  wire  _GEN_4260 = unuse_way == 2'h1 ? valid_1_23 : _GEN_3106; // @[cache.scala 22:26 82:34]
  wire  _GEN_4261 = unuse_way == 2'h1 ? valid_1_24 : _GEN_3107; // @[cache.scala 22:26 82:34]
  wire  _GEN_4262 = unuse_way == 2'h1 ? valid_1_25 : _GEN_3108; // @[cache.scala 22:26 82:34]
  wire  _GEN_4263 = unuse_way == 2'h1 ? valid_1_26 : _GEN_3109; // @[cache.scala 22:26 82:34]
  wire  _GEN_4264 = unuse_way == 2'h1 ? valid_1_27 : _GEN_3110; // @[cache.scala 22:26 82:34]
  wire  _GEN_4265 = unuse_way == 2'h1 ? valid_1_28 : _GEN_3111; // @[cache.scala 22:26 82:34]
  wire  _GEN_4266 = unuse_way == 2'h1 ? valid_1_29 : _GEN_3112; // @[cache.scala 22:26 82:34]
  wire  _GEN_4267 = unuse_way == 2'h1 ? valid_1_30 : _GEN_3113; // @[cache.scala 22:26 82:34]
  wire  _GEN_4268 = unuse_way == 2'h1 ? valid_1_31 : _GEN_3114; // @[cache.scala 22:26 82:34]
  wire  _GEN_4269 = unuse_way == 2'h1 ? valid_1_32 : _GEN_3115; // @[cache.scala 22:26 82:34]
  wire  _GEN_4270 = unuse_way == 2'h1 ? valid_1_33 : _GEN_3116; // @[cache.scala 22:26 82:34]
  wire  _GEN_4271 = unuse_way == 2'h1 ? valid_1_34 : _GEN_3117; // @[cache.scala 22:26 82:34]
  wire  _GEN_4272 = unuse_way == 2'h1 ? valid_1_35 : _GEN_3118; // @[cache.scala 22:26 82:34]
  wire  _GEN_4273 = unuse_way == 2'h1 ? valid_1_36 : _GEN_3119; // @[cache.scala 22:26 82:34]
  wire  _GEN_4274 = unuse_way == 2'h1 ? valid_1_37 : _GEN_3120; // @[cache.scala 22:26 82:34]
  wire  _GEN_4275 = unuse_way == 2'h1 ? valid_1_38 : _GEN_3121; // @[cache.scala 22:26 82:34]
  wire  _GEN_4276 = unuse_way == 2'h1 ? valid_1_39 : _GEN_3122; // @[cache.scala 22:26 82:34]
  wire  _GEN_4277 = unuse_way == 2'h1 ? valid_1_40 : _GEN_3123; // @[cache.scala 22:26 82:34]
  wire  _GEN_4278 = unuse_way == 2'h1 ? valid_1_41 : _GEN_3124; // @[cache.scala 22:26 82:34]
  wire  _GEN_4279 = unuse_way == 2'h1 ? valid_1_42 : _GEN_3125; // @[cache.scala 22:26 82:34]
  wire  _GEN_4280 = unuse_way == 2'h1 ? valid_1_43 : _GEN_3126; // @[cache.scala 22:26 82:34]
  wire  _GEN_4281 = unuse_way == 2'h1 ? valid_1_44 : _GEN_3127; // @[cache.scala 22:26 82:34]
  wire  _GEN_4282 = unuse_way == 2'h1 ? valid_1_45 : _GEN_3128; // @[cache.scala 22:26 82:34]
  wire  _GEN_4283 = unuse_way == 2'h1 ? valid_1_46 : _GEN_3129; // @[cache.scala 22:26 82:34]
  wire  _GEN_4284 = unuse_way == 2'h1 ? valid_1_47 : _GEN_3130; // @[cache.scala 22:26 82:34]
  wire  _GEN_4285 = unuse_way == 2'h1 ? valid_1_48 : _GEN_3131; // @[cache.scala 22:26 82:34]
  wire  _GEN_4286 = unuse_way == 2'h1 ? valid_1_49 : _GEN_3132; // @[cache.scala 22:26 82:34]
  wire  _GEN_4287 = unuse_way == 2'h1 ? valid_1_50 : _GEN_3133; // @[cache.scala 22:26 82:34]
  wire  _GEN_4288 = unuse_way == 2'h1 ? valid_1_51 : _GEN_3134; // @[cache.scala 22:26 82:34]
  wire  _GEN_4289 = unuse_way == 2'h1 ? valid_1_52 : _GEN_3135; // @[cache.scala 22:26 82:34]
  wire  _GEN_4290 = unuse_way == 2'h1 ? valid_1_53 : _GEN_3136; // @[cache.scala 22:26 82:34]
  wire  _GEN_4291 = unuse_way == 2'h1 ? valid_1_54 : _GEN_3137; // @[cache.scala 22:26 82:34]
  wire  _GEN_4292 = unuse_way == 2'h1 ? valid_1_55 : _GEN_3138; // @[cache.scala 22:26 82:34]
  wire  _GEN_4293 = unuse_way == 2'h1 ? valid_1_56 : _GEN_3139; // @[cache.scala 22:26 82:34]
  wire  _GEN_4294 = unuse_way == 2'h1 ? valid_1_57 : _GEN_3140; // @[cache.scala 22:26 82:34]
  wire  _GEN_4295 = unuse_way == 2'h1 ? valid_1_58 : _GEN_3141; // @[cache.scala 22:26 82:34]
  wire  _GEN_4296 = unuse_way == 2'h1 ? valid_1_59 : _GEN_3142; // @[cache.scala 22:26 82:34]
  wire  _GEN_4297 = unuse_way == 2'h1 ? valid_1_60 : _GEN_3143; // @[cache.scala 22:26 82:34]
  wire  _GEN_4298 = unuse_way == 2'h1 ? valid_1_61 : _GEN_3144; // @[cache.scala 22:26 82:34]
  wire  _GEN_4299 = unuse_way == 2'h1 ? valid_1_62 : _GEN_3145; // @[cache.scala 22:26 82:34]
  wire  _GEN_4300 = unuse_way == 2'h1 ? valid_1_63 : _GEN_3146; // @[cache.scala 22:26 82:34]
  wire  _GEN_4301 = unuse_way == 2'h1 ? valid_1_64 : _GEN_3147; // @[cache.scala 22:26 82:34]
  wire  _GEN_4302 = unuse_way == 2'h1 ? valid_1_65 : _GEN_3148; // @[cache.scala 22:26 82:34]
  wire  _GEN_4303 = unuse_way == 2'h1 ? valid_1_66 : _GEN_3149; // @[cache.scala 22:26 82:34]
  wire  _GEN_4304 = unuse_way == 2'h1 ? valid_1_67 : _GEN_3150; // @[cache.scala 22:26 82:34]
  wire  _GEN_4305 = unuse_way == 2'h1 ? valid_1_68 : _GEN_3151; // @[cache.scala 22:26 82:34]
  wire  _GEN_4306 = unuse_way == 2'h1 ? valid_1_69 : _GEN_3152; // @[cache.scala 22:26 82:34]
  wire  _GEN_4307 = unuse_way == 2'h1 ? valid_1_70 : _GEN_3153; // @[cache.scala 22:26 82:34]
  wire  _GEN_4308 = unuse_way == 2'h1 ? valid_1_71 : _GEN_3154; // @[cache.scala 22:26 82:34]
  wire  _GEN_4309 = unuse_way == 2'h1 ? valid_1_72 : _GEN_3155; // @[cache.scala 22:26 82:34]
  wire  _GEN_4310 = unuse_way == 2'h1 ? valid_1_73 : _GEN_3156; // @[cache.scala 22:26 82:34]
  wire  _GEN_4311 = unuse_way == 2'h1 ? valid_1_74 : _GEN_3157; // @[cache.scala 22:26 82:34]
  wire  _GEN_4312 = unuse_way == 2'h1 ? valid_1_75 : _GEN_3158; // @[cache.scala 22:26 82:34]
  wire  _GEN_4313 = unuse_way == 2'h1 ? valid_1_76 : _GEN_3159; // @[cache.scala 22:26 82:34]
  wire  _GEN_4314 = unuse_way == 2'h1 ? valid_1_77 : _GEN_3160; // @[cache.scala 22:26 82:34]
  wire  _GEN_4315 = unuse_way == 2'h1 ? valid_1_78 : _GEN_3161; // @[cache.scala 22:26 82:34]
  wire  _GEN_4316 = unuse_way == 2'h1 ? valid_1_79 : _GEN_3162; // @[cache.scala 22:26 82:34]
  wire  _GEN_4317 = unuse_way == 2'h1 ? valid_1_80 : _GEN_3163; // @[cache.scala 22:26 82:34]
  wire  _GEN_4318 = unuse_way == 2'h1 ? valid_1_81 : _GEN_3164; // @[cache.scala 22:26 82:34]
  wire  _GEN_4319 = unuse_way == 2'h1 ? valid_1_82 : _GEN_3165; // @[cache.scala 22:26 82:34]
  wire  _GEN_4320 = unuse_way == 2'h1 ? valid_1_83 : _GEN_3166; // @[cache.scala 22:26 82:34]
  wire  _GEN_4321 = unuse_way == 2'h1 ? valid_1_84 : _GEN_3167; // @[cache.scala 22:26 82:34]
  wire  _GEN_4322 = unuse_way == 2'h1 ? valid_1_85 : _GEN_3168; // @[cache.scala 22:26 82:34]
  wire  _GEN_4323 = unuse_way == 2'h1 ? valid_1_86 : _GEN_3169; // @[cache.scala 22:26 82:34]
  wire  _GEN_4324 = unuse_way == 2'h1 ? valid_1_87 : _GEN_3170; // @[cache.scala 22:26 82:34]
  wire  _GEN_4325 = unuse_way == 2'h1 ? valid_1_88 : _GEN_3171; // @[cache.scala 22:26 82:34]
  wire  _GEN_4326 = unuse_way == 2'h1 ? valid_1_89 : _GEN_3172; // @[cache.scala 22:26 82:34]
  wire  _GEN_4327 = unuse_way == 2'h1 ? valid_1_90 : _GEN_3173; // @[cache.scala 22:26 82:34]
  wire  _GEN_4328 = unuse_way == 2'h1 ? valid_1_91 : _GEN_3174; // @[cache.scala 22:26 82:34]
  wire  _GEN_4329 = unuse_way == 2'h1 ? valid_1_92 : _GEN_3175; // @[cache.scala 22:26 82:34]
  wire  _GEN_4330 = unuse_way == 2'h1 ? valid_1_93 : _GEN_3176; // @[cache.scala 22:26 82:34]
  wire  _GEN_4331 = unuse_way == 2'h1 ? valid_1_94 : _GEN_3177; // @[cache.scala 22:26 82:34]
  wire  _GEN_4332 = unuse_way == 2'h1 ? valid_1_95 : _GEN_3178; // @[cache.scala 22:26 82:34]
  wire  _GEN_4333 = unuse_way == 2'h1 ? valid_1_96 : _GEN_3179; // @[cache.scala 22:26 82:34]
  wire  _GEN_4334 = unuse_way == 2'h1 ? valid_1_97 : _GEN_3180; // @[cache.scala 22:26 82:34]
  wire  _GEN_4335 = unuse_way == 2'h1 ? valid_1_98 : _GEN_3181; // @[cache.scala 22:26 82:34]
  wire  _GEN_4336 = unuse_way == 2'h1 ? valid_1_99 : _GEN_3182; // @[cache.scala 22:26 82:34]
  wire  _GEN_4337 = unuse_way == 2'h1 ? valid_1_100 : _GEN_3183; // @[cache.scala 22:26 82:34]
  wire  _GEN_4338 = unuse_way == 2'h1 ? valid_1_101 : _GEN_3184; // @[cache.scala 22:26 82:34]
  wire  _GEN_4339 = unuse_way == 2'h1 ? valid_1_102 : _GEN_3185; // @[cache.scala 22:26 82:34]
  wire  _GEN_4340 = unuse_way == 2'h1 ? valid_1_103 : _GEN_3186; // @[cache.scala 22:26 82:34]
  wire  _GEN_4341 = unuse_way == 2'h1 ? valid_1_104 : _GEN_3187; // @[cache.scala 22:26 82:34]
  wire  _GEN_4342 = unuse_way == 2'h1 ? valid_1_105 : _GEN_3188; // @[cache.scala 22:26 82:34]
  wire  _GEN_4343 = unuse_way == 2'h1 ? valid_1_106 : _GEN_3189; // @[cache.scala 22:26 82:34]
  wire  _GEN_4344 = unuse_way == 2'h1 ? valid_1_107 : _GEN_3190; // @[cache.scala 22:26 82:34]
  wire  _GEN_4345 = unuse_way == 2'h1 ? valid_1_108 : _GEN_3191; // @[cache.scala 22:26 82:34]
  wire  _GEN_4346 = unuse_way == 2'h1 ? valid_1_109 : _GEN_3192; // @[cache.scala 22:26 82:34]
  wire  _GEN_4347 = unuse_way == 2'h1 ? valid_1_110 : _GEN_3193; // @[cache.scala 22:26 82:34]
  wire  _GEN_4348 = unuse_way == 2'h1 ? valid_1_111 : _GEN_3194; // @[cache.scala 22:26 82:34]
  wire  _GEN_4349 = unuse_way == 2'h1 ? valid_1_112 : _GEN_3195; // @[cache.scala 22:26 82:34]
  wire  _GEN_4350 = unuse_way == 2'h1 ? valid_1_113 : _GEN_3196; // @[cache.scala 22:26 82:34]
  wire  _GEN_4351 = unuse_way == 2'h1 ? valid_1_114 : _GEN_3197; // @[cache.scala 22:26 82:34]
  wire  _GEN_4352 = unuse_way == 2'h1 ? valid_1_115 : _GEN_3198; // @[cache.scala 22:26 82:34]
  wire  _GEN_4353 = unuse_way == 2'h1 ? valid_1_116 : _GEN_3199; // @[cache.scala 22:26 82:34]
  wire  _GEN_4354 = unuse_way == 2'h1 ? valid_1_117 : _GEN_3200; // @[cache.scala 22:26 82:34]
  wire  _GEN_4355 = unuse_way == 2'h1 ? valid_1_118 : _GEN_3201; // @[cache.scala 22:26 82:34]
  wire  _GEN_4356 = unuse_way == 2'h1 ? valid_1_119 : _GEN_3202; // @[cache.scala 22:26 82:34]
  wire  _GEN_4357 = unuse_way == 2'h1 ? valid_1_120 : _GEN_3203; // @[cache.scala 22:26 82:34]
  wire  _GEN_4358 = unuse_way == 2'h1 ? valid_1_121 : _GEN_3204; // @[cache.scala 22:26 82:34]
  wire  _GEN_4359 = unuse_way == 2'h1 ? valid_1_122 : _GEN_3205; // @[cache.scala 22:26 82:34]
  wire  _GEN_4360 = unuse_way == 2'h1 ? valid_1_123 : _GEN_3206; // @[cache.scala 22:26 82:34]
  wire  _GEN_4361 = unuse_way == 2'h1 ? valid_1_124 : _GEN_3207; // @[cache.scala 22:26 82:34]
  wire  _GEN_4362 = unuse_way == 2'h1 ? valid_1_125 : _GEN_3208; // @[cache.scala 22:26 82:34]
  wire  _GEN_4363 = unuse_way == 2'h1 ? valid_1_126 : _GEN_3209; // @[cache.scala 22:26 82:34]
  wire  _GEN_4364 = unuse_way == 2'h1 ? valid_1_127 : _GEN_3210; // @[cache.scala 22:26 82:34]
  wire [1:0] _GEN_4365 = 2'h3 == state ? 2'h0 : state; // @[cache.scala 51:18 81:19 49:24]
  wire [63:0] _GEN_4366 = 2'h3 == state ? _GEN_3596 : ram_0_0; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4367 = 2'h3 == state ? _GEN_3597 : ram_0_1; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4368 = 2'h3 == state ? _GEN_3598 : ram_0_2; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4369 = 2'h3 == state ? _GEN_3599 : ram_0_3; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4370 = 2'h3 == state ? _GEN_3600 : ram_0_4; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4371 = 2'h3 == state ? _GEN_3601 : ram_0_5; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4372 = 2'h3 == state ? _GEN_3602 : ram_0_6; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4373 = 2'h3 == state ? _GEN_3603 : ram_0_7; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4374 = 2'h3 == state ? _GEN_3604 : ram_0_8; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4375 = 2'h3 == state ? _GEN_3605 : ram_0_9; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4376 = 2'h3 == state ? _GEN_3606 : ram_0_10; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4377 = 2'h3 == state ? _GEN_3607 : ram_0_11; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4378 = 2'h3 == state ? _GEN_3608 : ram_0_12; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4379 = 2'h3 == state ? _GEN_3609 : ram_0_13; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4380 = 2'h3 == state ? _GEN_3610 : ram_0_14; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4381 = 2'h3 == state ? _GEN_3611 : ram_0_15; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4382 = 2'h3 == state ? _GEN_3612 : ram_0_16; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4383 = 2'h3 == state ? _GEN_3613 : ram_0_17; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4384 = 2'h3 == state ? _GEN_3614 : ram_0_18; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4385 = 2'h3 == state ? _GEN_3615 : ram_0_19; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4386 = 2'h3 == state ? _GEN_3616 : ram_0_20; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4387 = 2'h3 == state ? _GEN_3617 : ram_0_21; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4388 = 2'h3 == state ? _GEN_3618 : ram_0_22; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4389 = 2'h3 == state ? _GEN_3619 : ram_0_23; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4390 = 2'h3 == state ? _GEN_3620 : ram_0_24; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4391 = 2'h3 == state ? _GEN_3621 : ram_0_25; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4392 = 2'h3 == state ? _GEN_3622 : ram_0_26; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4393 = 2'h3 == state ? _GEN_3623 : ram_0_27; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4394 = 2'h3 == state ? _GEN_3624 : ram_0_28; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4395 = 2'h3 == state ? _GEN_3625 : ram_0_29; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4396 = 2'h3 == state ? _GEN_3626 : ram_0_30; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4397 = 2'h3 == state ? _GEN_3627 : ram_0_31; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4398 = 2'h3 == state ? _GEN_3628 : ram_0_32; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4399 = 2'h3 == state ? _GEN_3629 : ram_0_33; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4400 = 2'h3 == state ? _GEN_3630 : ram_0_34; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4401 = 2'h3 == state ? _GEN_3631 : ram_0_35; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4402 = 2'h3 == state ? _GEN_3632 : ram_0_36; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4403 = 2'h3 == state ? _GEN_3633 : ram_0_37; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4404 = 2'h3 == state ? _GEN_3634 : ram_0_38; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4405 = 2'h3 == state ? _GEN_3635 : ram_0_39; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4406 = 2'h3 == state ? _GEN_3636 : ram_0_40; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4407 = 2'h3 == state ? _GEN_3637 : ram_0_41; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4408 = 2'h3 == state ? _GEN_3638 : ram_0_42; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4409 = 2'h3 == state ? _GEN_3639 : ram_0_43; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4410 = 2'h3 == state ? _GEN_3640 : ram_0_44; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4411 = 2'h3 == state ? _GEN_3641 : ram_0_45; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4412 = 2'h3 == state ? _GEN_3642 : ram_0_46; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4413 = 2'h3 == state ? _GEN_3643 : ram_0_47; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4414 = 2'h3 == state ? _GEN_3644 : ram_0_48; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4415 = 2'h3 == state ? _GEN_3645 : ram_0_49; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4416 = 2'h3 == state ? _GEN_3646 : ram_0_50; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4417 = 2'h3 == state ? _GEN_3647 : ram_0_51; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4418 = 2'h3 == state ? _GEN_3648 : ram_0_52; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4419 = 2'h3 == state ? _GEN_3649 : ram_0_53; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4420 = 2'h3 == state ? _GEN_3650 : ram_0_54; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4421 = 2'h3 == state ? _GEN_3651 : ram_0_55; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4422 = 2'h3 == state ? _GEN_3652 : ram_0_56; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4423 = 2'h3 == state ? _GEN_3653 : ram_0_57; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4424 = 2'h3 == state ? _GEN_3654 : ram_0_58; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4425 = 2'h3 == state ? _GEN_3655 : ram_0_59; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4426 = 2'h3 == state ? _GEN_3656 : ram_0_60; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4427 = 2'h3 == state ? _GEN_3657 : ram_0_61; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4428 = 2'h3 == state ? _GEN_3658 : ram_0_62; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4429 = 2'h3 == state ? _GEN_3659 : ram_0_63; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4430 = 2'h3 == state ? _GEN_3660 : ram_0_64; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4431 = 2'h3 == state ? _GEN_3661 : ram_0_65; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4432 = 2'h3 == state ? _GEN_3662 : ram_0_66; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4433 = 2'h3 == state ? _GEN_3663 : ram_0_67; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4434 = 2'h3 == state ? _GEN_3664 : ram_0_68; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4435 = 2'h3 == state ? _GEN_3665 : ram_0_69; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4436 = 2'h3 == state ? _GEN_3666 : ram_0_70; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4437 = 2'h3 == state ? _GEN_3667 : ram_0_71; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4438 = 2'h3 == state ? _GEN_3668 : ram_0_72; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4439 = 2'h3 == state ? _GEN_3669 : ram_0_73; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4440 = 2'h3 == state ? _GEN_3670 : ram_0_74; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4441 = 2'h3 == state ? _GEN_3671 : ram_0_75; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4442 = 2'h3 == state ? _GEN_3672 : ram_0_76; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4443 = 2'h3 == state ? _GEN_3673 : ram_0_77; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4444 = 2'h3 == state ? _GEN_3674 : ram_0_78; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4445 = 2'h3 == state ? _GEN_3675 : ram_0_79; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4446 = 2'h3 == state ? _GEN_3676 : ram_0_80; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4447 = 2'h3 == state ? _GEN_3677 : ram_0_81; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4448 = 2'h3 == state ? _GEN_3678 : ram_0_82; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4449 = 2'h3 == state ? _GEN_3679 : ram_0_83; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4450 = 2'h3 == state ? _GEN_3680 : ram_0_84; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4451 = 2'h3 == state ? _GEN_3681 : ram_0_85; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4452 = 2'h3 == state ? _GEN_3682 : ram_0_86; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4453 = 2'h3 == state ? _GEN_3683 : ram_0_87; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4454 = 2'h3 == state ? _GEN_3684 : ram_0_88; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4455 = 2'h3 == state ? _GEN_3685 : ram_0_89; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4456 = 2'h3 == state ? _GEN_3686 : ram_0_90; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4457 = 2'h3 == state ? _GEN_3687 : ram_0_91; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4458 = 2'h3 == state ? _GEN_3688 : ram_0_92; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4459 = 2'h3 == state ? _GEN_3689 : ram_0_93; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4460 = 2'h3 == state ? _GEN_3690 : ram_0_94; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4461 = 2'h3 == state ? _GEN_3691 : ram_0_95; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4462 = 2'h3 == state ? _GEN_3692 : ram_0_96; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4463 = 2'h3 == state ? _GEN_3693 : ram_0_97; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4464 = 2'h3 == state ? _GEN_3694 : ram_0_98; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4465 = 2'h3 == state ? _GEN_3695 : ram_0_99; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4466 = 2'h3 == state ? _GEN_3696 : ram_0_100; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4467 = 2'h3 == state ? _GEN_3697 : ram_0_101; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4468 = 2'h3 == state ? _GEN_3698 : ram_0_102; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4469 = 2'h3 == state ? _GEN_3699 : ram_0_103; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4470 = 2'h3 == state ? _GEN_3700 : ram_0_104; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4471 = 2'h3 == state ? _GEN_3701 : ram_0_105; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4472 = 2'h3 == state ? _GEN_3702 : ram_0_106; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4473 = 2'h3 == state ? _GEN_3703 : ram_0_107; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4474 = 2'h3 == state ? _GEN_3704 : ram_0_108; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4475 = 2'h3 == state ? _GEN_3705 : ram_0_109; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4476 = 2'h3 == state ? _GEN_3706 : ram_0_110; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4477 = 2'h3 == state ? _GEN_3707 : ram_0_111; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4478 = 2'h3 == state ? _GEN_3708 : ram_0_112; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4479 = 2'h3 == state ? _GEN_3709 : ram_0_113; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4480 = 2'h3 == state ? _GEN_3710 : ram_0_114; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4481 = 2'h3 == state ? _GEN_3711 : ram_0_115; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4482 = 2'h3 == state ? _GEN_3712 : ram_0_116; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4483 = 2'h3 == state ? _GEN_3713 : ram_0_117; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4484 = 2'h3 == state ? _GEN_3714 : ram_0_118; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4485 = 2'h3 == state ? _GEN_3715 : ram_0_119; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4486 = 2'h3 == state ? _GEN_3716 : ram_0_120; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4487 = 2'h3 == state ? _GEN_3717 : ram_0_121; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4488 = 2'h3 == state ? _GEN_3718 : ram_0_122; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4489 = 2'h3 == state ? _GEN_3719 : ram_0_123; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4490 = 2'h3 == state ? _GEN_3720 : ram_0_124; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4491 = 2'h3 == state ? _GEN_3721 : ram_0_125; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4492 = 2'h3 == state ? _GEN_3722 : ram_0_126; // @[cache.scala 51:18 17:24]
  wire [63:0] _GEN_4493 = 2'h3 == state ? _GEN_3723 : ram_0_127; // @[cache.scala 51:18 17:24]
  wire [31:0] _GEN_4494 = 2'h3 == state ? _GEN_3724 : tag_0_0; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4495 = 2'h3 == state ? _GEN_3725 : tag_0_1; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4496 = 2'h3 == state ? _GEN_3726 : tag_0_2; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4497 = 2'h3 == state ? _GEN_3727 : tag_0_3; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4498 = 2'h3 == state ? _GEN_3728 : tag_0_4; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4499 = 2'h3 == state ? _GEN_3729 : tag_0_5; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4500 = 2'h3 == state ? _GEN_3730 : tag_0_6; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4501 = 2'h3 == state ? _GEN_3731 : tag_0_7; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4502 = 2'h3 == state ? _GEN_3732 : tag_0_8; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4503 = 2'h3 == state ? _GEN_3733 : tag_0_9; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4504 = 2'h3 == state ? _GEN_3734 : tag_0_10; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4505 = 2'h3 == state ? _GEN_3735 : tag_0_11; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4506 = 2'h3 == state ? _GEN_3736 : tag_0_12; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4507 = 2'h3 == state ? _GEN_3737 : tag_0_13; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4508 = 2'h3 == state ? _GEN_3738 : tag_0_14; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4509 = 2'h3 == state ? _GEN_3739 : tag_0_15; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4510 = 2'h3 == state ? _GEN_3740 : tag_0_16; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4511 = 2'h3 == state ? _GEN_3741 : tag_0_17; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4512 = 2'h3 == state ? _GEN_3742 : tag_0_18; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4513 = 2'h3 == state ? _GEN_3743 : tag_0_19; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4514 = 2'h3 == state ? _GEN_3744 : tag_0_20; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4515 = 2'h3 == state ? _GEN_3745 : tag_0_21; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4516 = 2'h3 == state ? _GEN_3746 : tag_0_22; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4517 = 2'h3 == state ? _GEN_3747 : tag_0_23; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4518 = 2'h3 == state ? _GEN_3748 : tag_0_24; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4519 = 2'h3 == state ? _GEN_3749 : tag_0_25; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4520 = 2'h3 == state ? _GEN_3750 : tag_0_26; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4521 = 2'h3 == state ? _GEN_3751 : tag_0_27; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4522 = 2'h3 == state ? _GEN_3752 : tag_0_28; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4523 = 2'h3 == state ? _GEN_3753 : tag_0_29; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4524 = 2'h3 == state ? _GEN_3754 : tag_0_30; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4525 = 2'h3 == state ? _GEN_3755 : tag_0_31; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4526 = 2'h3 == state ? _GEN_3756 : tag_0_32; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4527 = 2'h3 == state ? _GEN_3757 : tag_0_33; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4528 = 2'h3 == state ? _GEN_3758 : tag_0_34; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4529 = 2'h3 == state ? _GEN_3759 : tag_0_35; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4530 = 2'h3 == state ? _GEN_3760 : tag_0_36; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4531 = 2'h3 == state ? _GEN_3761 : tag_0_37; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4532 = 2'h3 == state ? _GEN_3762 : tag_0_38; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4533 = 2'h3 == state ? _GEN_3763 : tag_0_39; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4534 = 2'h3 == state ? _GEN_3764 : tag_0_40; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4535 = 2'h3 == state ? _GEN_3765 : tag_0_41; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4536 = 2'h3 == state ? _GEN_3766 : tag_0_42; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4537 = 2'h3 == state ? _GEN_3767 : tag_0_43; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4538 = 2'h3 == state ? _GEN_3768 : tag_0_44; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4539 = 2'h3 == state ? _GEN_3769 : tag_0_45; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4540 = 2'h3 == state ? _GEN_3770 : tag_0_46; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4541 = 2'h3 == state ? _GEN_3771 : tag_0_47; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4542 = 2'h3 == state ? _GEN_3772 : tag_0_48; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4543 = 2'h3 == state ? _GEN_3773 : tag_0_49; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4544 = 2'h3 == state ? _GEN_3774 : tag_0_50; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4545 = 2'h3 == state ? _GEN_3775 : tag_0_51; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4546 = 2'h3 == state ? _GEN_3776 : tag_0_52; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4547 = 2'h3 == state ? _GEN_3777 : tag_0_53; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4548 = 2'h3 == state ? _GEN_3778 : tag_0_54; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4549 = 2'h3 == state ? _GEN_3779 : tag_0_55; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4550 = 2'h3 == state ? _GEN_3780 : tag_0_56; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4551 = 2'h3 == state ? _GEN_3781 : tag_0_57; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4552 = 2'h3 == state ? _GEN_3782 : tag_0_58; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4553 = 2'h3 == state ? _GEN_3783 : tag_0_59; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4554 = 2'h3 == state ? _GEN_3784 : tag_0_60; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4555 = 2'h3 == state ? _GEN_3785 : tag_0_61; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4556 = 2'h3 == state ? _GEN_3786 : tag_0_62; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4557 = 2'h3 == state ? _GEN_3787 : tag_0_63; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4558 = 2'h3 == state ? _GEN_3788 : tag_0_64; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4559 = 2'h3 == state ? _GEN_3789 : tag_0_65; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4560 = 2'h3 == state ? _GEN_3790 : tag_0_66; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4561 = 2'h3 == state ? _GEN_3791 : tag_0_67; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4562 = 2'h3 == state ? _GEN_3792 : tag_0_68; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4563 = 2'h3 == state ? _GEN_3793 : tag_0_69; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4564 = 2'h3 == state ? _GEN_3794 : tag_0_70; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4565 = 2'h3 == state ? _GEN_3795 : tag_0_71; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4566 = 2'h3 == state ? _GEN_3796 : tag_0_72; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4567 = 2'h3 == state ? _GEN_3797 : tag_0_73; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4568 = 2'h3 == state ? _GEN_3798 : tag_0_74; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4569 = 2'h3 == state ? _GEN_3799 : tag_0_75; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4570 = 2'h3 == state ? _GEN_3800 : tag_0_76; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4571 = 2'h3 == state ? _GEN_3801 : tag_0_77; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4572 = 2'h3 == state ? _GEN_3802 : tag_0_78; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4573 = 2'h3 == state ? _GEN_3803 : tag_0_79; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4574 = 2'h3 == state ? _GEN_3804 : tag_0_80; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4575 = 2'h3 == state ? _GEN_3805 : tag_0_81; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4576 = 2'h3 == state ? _GEN_3806 : tag_0_82; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4577 = 2'h3 == state ? _GEN_3807 : tag_0_83; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4578 = 2'h3 == state ? _GEN_3808 : tag_0_84; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4579 = 2'h3 == state ? _GEN_3809 : tag_0_85; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4580 = 2'h3 == state ? _GEN_3810 : tag_0_86; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4581 = 2'h3 == state ? _GEN_3811 : tag_0_87; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4582 = 2'h3 == state ? _GEN_3812 : tag_0_88; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4583 = 2'h3 == state ? _GEN_3813 : tag_0_89; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4584 = 2'h3 == state ? _GEN_3814 : tag_0_90; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4585 = 2'h3 == state ? _GEN_3815 : tag_0_91; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4586 = 2'h3 == state ? _GEN_3816 : tag_0_92; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4587 = 2'h3 == state ? _GEN_3817 : tag_0_93; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4588 = 2'h3 == state ? _GEN_3818 : tag_0_94; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4589 = 2'h3 == state ? _GEN_3819 : tag_0_95; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4590 = 2'h3 == state ? _GEN_3820 : tag_0_96; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4591 = 2'h3 == state ? _GEN_3821 : tag_0_97; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4592 = 2'h3 == state ? _GEN_3822 : tag_0_98; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4593 = 2'h3 == state ? _GEN_3823 : tag_0_99; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4594 = 2'h3 == state ? _GEN_3824 : tag_0_100; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4595 = 2'h3 == state ? _GEN_3825 : tag_0_101; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4596 = 2'h3 == state ? _GEN_3826 : tag_0_102; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4597 = 2'h3 == state ? _GEN_3827 : tag_0_103; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4598 = 2'h3 == state ? _GEN_3828 : tag_0_104; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4599 = 2'h3 == state ? _GEN_3829 : tag_0_105; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4600 = 2'h3 == state ? _GEN_3830 : tag_0_106; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4601 = 2'h3 == state ? _GEN_3831 : tag_0_107; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4602 = 2'h3 == state ? _GEN_3832 : tag_0_108; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4603 = 2'h3 == state ? _GEN_3833 : tag_0_109; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4604 = 2'h3 == state ? _GEN_3834 : tag_0_110; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4605 = 2'h3 == state ? _GEN_3835 : tag_0_111; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4606 = 2'h3 == state ? _GEN_3836 : tag_0_112; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4607 = 2'h3 == state ? _GEN_3837 : tag_0_113; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4608 = 2'h3 == state ? _GEN_3838 : tag_0_114; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4609 = 2'h3 == state ? _GEN_3839 : tag_0_115; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4610 = 2'h3 == state ? _GEN_3840 : tag_0_116; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4611 = 2'h3 == state ? _GEN_3841 : tag_0_117; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4612 = 2'h3 == state ? _GEN_3842 : tag_0_118; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4613 = 2'h3 == state ? _GEN_3843 : tag_0_119; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4614 = 2'h3 == state ? _GEN_3844 : tag_0_120; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4615 = 2'h3 == state ? _GEN_3845 : tag_0_121; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4616 = 2'h3 == state ? _GEN_3846 : tag_0_122; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4617 = 2'h3 == state ? _GEN_3847 : tag_0_123; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4618 = 2'h3 == state ? _GEN_3848 : tag_0_124; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4619 = 2'h3 == state ? _GEN_3849 : tag_0_125; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4620 = 2'h3 == state ? _GEN_3850 : tag_0_126; // @[cache.scala 51:18 19:24]
  wire [31:0] _GEN_4621 = 2'h3 == state ? _GEN_3851 : tag_0_127; // @[cache.scala 51:18 19:24]
  wire  _GEN_4622 = 2'h3 == state ? _GEN_3852 : valid_0_0; // @[cache.scala 51:18 21:26]
  wire  _GEN_4623 = 2'h3 == state ? _GEN_3853 : valid_0_1; // @[cache.scala 51:18 21:26]
  wire  _GEN_4624 = 2'h3 == state ? _GEN_3854 : valid_0_2; // @[cache.scala 51:18 21:26]
  wire  _GEN_4625 = 2'h3 == state ? _GEN_3855 : valid_0_3; // @[cache.scala 51:18 21:26]
  wire  _GEN_4626 = 2'h3 == state ? _GEN_3856 : valid_0_4; // @[cache.scala 51:18 21:26]
  wire  _GEN_4627 = 2'h3 == state ? _GEN_3857 : valid_0_5; // @[cache.scala 51:18 21:26]
  wire  _GEN_4628 = 2'h3 == state ? _GEN_3858 : valid_0_6; // @[cache.scala 51:18 21:26]
  wire  _GEN_4629 = 2'h3 == state ? _GEN_3859 : valid_0_7; // @[cache.scala 51:18 21:26]
  wire  _GEN_4630 = 2'h3 == state ? _GEN_3860 : valid_0_8; // @[cache.scala 51:18 21:26]
  wire  _GEN_4631 = 2'h3 == state ? _GEN_3861 : valid_0_9; // @[cache.scala 51:18 21:26]
  wire  _GEN_4632 = 2'h3 == state ? _GEN_3862 : valid_0_10; // @[cache.scala 51:18 21:26]
  wire  _GEN_4633 = 2'h3 == state ? _GEN_3863 : valid_0_11; // @[cache.scala 51:18 21:26]
  wire  _GEN_4634 = 2'h3 == state ? _GEN_3864 : valid_0_12; // @[cache.scala 51:18 21:26]
  wire  _GEN_4635 = 2'h3 == state ? _GEN_3865 : valid_0_13; // @[cache.scala 51:18 21:26]
  wire  _GEN_4636 = 2'h3 == state ? _GEN_3866 : valid_0_14; // @[cache.scala 51:18 21:26]
  wire  _GEN_4637 = 2'h3 == state ? _GEN_3867 : valid_0_15; // @[cache.scala 51:18 21:26]
  wire  _GEN_4638 = 2'h3 == state ? _GEN_3868 : valid_0_16; // @[cache.scala 51:18 21:26]
  wire  _GEN_4639 = 2'h3 == state ? _GEN_3869 : valid_0_17; // @[cache.scala 51:18 21:26]
  wire  _GEN_4640 = 2'h3 == state ? _GEN_3870 : valid_0_18; // @[cache.scala 51:18 21:26]
  wire  _GEN_4641 = 2'h3 == state ? _GEN_3871 : valid_0_19; // @[cache.scala 51:18 21:26]
  wire  _GEN_4642 = 2'h3 == state ? _GEN_3872 : valid_0_20; // @[cache.scala 51:18 21:26]
  wire  _GEN_4643 = 2'h3 == state ? _GEN_3873 : valid_0_21; // @[cache.scala 51:18 21:26]
  wire  _GEN_4644 = 2'h3 == state ? _GEN_3874 : valid_0_22; // @[cache.scala 51:18 21:26]
  wire  _GEN_4645 = 2'h3 == state ? _GEN_3875 : valid_0_23; // @[cache.scala 51:18 21:26]
  wire  _GEN_4646 = 2'h3 == state ? _GEN_3876 : valid_0_24; // @[cache.scala 51:18 21:26]
  wire  _GEN_4647 = 2'h3 == state ? _GEN_3877 : valid_0_25; // @[cache.scala 51:18 21:26]
  wire  _GEN_4648 = 2'h3 == state ? _GEN_3878 : valid_0_26; // @[cache.scala 51:18 21:26]
  wire  _GEN_4649 = 2'h3 == state ? _GEN_3879 : valid_0_27; // @[cache.scala 51:18 21:26]
  wire  _GEN_4650 = 2'h3 == state ? _GEN_3880 : valid_0_28; // @[cache.scala 51:18 21:26]
  wire  _GEN_4651 = 2'h3 == state ? _GEN_3881 : valid_0_29; // @[cache.scala 51:18 21:26]
  wire  _GEN_4652 = 2'h3 == state ? _GEN_3882 : valid_0_30; // @[cache.scala 51:18 21:26]
  wire  _GEN_4653 = 2'h3 == state ? _GEN_3883 : valid_0_31; // @[cache.scala 51:18 21:26]
  wire  _GEN_4654 = 2'h3 == state ? _GEN_3884 : valid_0_32; // @[cache.scala 51:18 21:26]
  wire  _GEN_4655 = 2'h3 == state ? _GEN_3885 : valid_0_33; // @[cache.scala 51:18 21:26]
  wire  _GEN_4656 = 2'h3 == state ? _GEN_3886 : valid_0_34; // @[cache.scala 51:18 21:26]
  wire  _GEN_4657 = 2'h3 == state ? _GEN_3887 : valid_0_35; // @[cache.scala 51:18 21:26]
  wire  _GEN_4658 = 2'h3 == state ? _GEN_3888 : valid_0_36; // @[cache.scala 51:18 21:26]
  wire  _GEN_4659 = 2'h3 == state ? _GEN_3889 : valid_0_37; // @[cache.scala 51:18 21:26]
  wire  _GEN_4660 = 2'h3 == state ? _GEN_3890 : valid_0_38; // @[cache.scala 51:18 21:26]
  wire  _GEN_4661 = 2'h3 == state ? _GEN_3891 : valid_0_39; // @[cache.scala 51:18 21:26]
  wire  _GEN_4662 = 2'h3 == state ? _GEN_3892 : valid_0_40; // @[cache.scala 51:18 21:26]
  wire  _GEN_4663 = 2'h3 == state ? _GEN_3893 : valid_0_41; // @[cache.scala 51:18 21:26]
  wire  _GEN_4664 = 2'h3 == state ? _GEN_3894 : valid_0_42; // @[cache.scala 51:18 21:26]
  wire  _GEN_4665 = 2'h3 == state ? _GEN_3895 : valid_0_43; // @[cache.scala 51:18 21:26]
  wire  _GEN_4666 = 2'h3 == state ? _GEN_3896 : valid_0_44; // @[cache.scala 51:18 21:26]
  wire  _GEN_4667 = 2'h3 == state ? _GEN_3897 : valid_0_45; // @[cache.scala 51:18 21:26]
  wire  _GEN_4668 = 2'h3 == state ? _GEN_3898 : valid_0_46; // @[cache.scala 51:18 21:26]
  wire  _GEN_4669 = 2'h3 == state ? _GEN_3899 : valid_0_47; // @[cache.scala 51:18 21:26]
  wire  _GEN_4670 = 2'h3 == state ? _GEN_3900 : valid_0_48; // @[cache.scala 51:18 21:26]
  wire  _GEN_4671 = 2'h3 == state ? _GEN_3901 : valid_0_49; // @[cache.scala 51:18 21:26]
  wire  _GEN_4672 = 2'h3 == state ? _GEN_3902 : valid_0_50; // @[cache.scala 51:18 21:26]
  wire  _GEN_4673 = 2'h3 == state ? _GEN_3903 : valid_0_51; // @[cache.scala 51:18 21:26]
  wire  _GEN_4674 = 2'h3 == state ? _GEN_3904 : valid_0_52; // @[cache.scala 51:18 21:26]
  wire  _GEN_4675 = 2'h3 == state ? _GEN_3905 : valid_0_53; // @[cache.scala 51:18 21:26]
  wire  _GEN_4676 = 2'h3 == state ? _GEN_3906 : valid_0_54; // @[cache.scala 51:18 21:26]
  wire  _GEN_4677 = 2'h3 == state ? _GEN_3907 : valid_0_55; // @[cache.scala 51:18 21:26]
  wire  _GEN_4678 = 2'h3 == state ? _GEN_3908 : valid_0_56; // @[cache.scala 51:18 21:26]
  wire  _GEN_4679 = 2'h3 == state ? _GEN_3909 : valid_0_57; // @[cache.scala 51:18 21:26]
  wire  _GEN_4680 = 2'h3 == state ? _GEN_3910 : valid_0_58; // @[cache.scala 51:18 21:26]
  wire  _GEN_4681 = 2'h3 == state ? _GEN_3911 : valid_0_59; // @[cache.scala 51:18 21:26]
  wire  _GEN_4682 = 2'h3 == state ? _GEN_3912 : valid_0_60; // @[cache.scala 51:18 21:26]
  wire  _GEN_4683 = 2'h3 == state ? _GEN_3913 : valid_0_61; // @[cache.scala 51:18 21:26]
  wire  _GEN_4684 = 2'h3 == state ? _GEN_3914 : valid_0_62; // @[cache.scala 51:18 21:26]
  wire  _GEN_4685 = 2'h3 == state ? _GEN_3915 : valid_0_63; // @[cache.scala 51:18 21:26]
  wire  _GEN_4686 = 2'h3 == state ? _GEN_3916 : valid_0_64; // @[cache.scala 51:18 21:26]
  wire  _GEN_4687 = 2'h3 == state ? _GEN_3917 : valid_0_65; // @[cache.scala 51:18 21:26]
  wire  _GEN_4688 = 2'h3 == state ? _GEN_3918 : valid_0_66; // @[cache.scala 51:18 21:26]
  wire  _GEN_4689 = 2'h3 == state ? _GEN_3919 : valid_0_67; // @[cache.scala 51:18 21:26]
  wire  _GEN_4690 = 2'h3 == state ? _GEN_3920 : valid_0_68; // @[cache.scala 51:18 21:26]
  wire  _GEN_4691 = 2'h3 == state ? _GEN_3921 : valid_0_69; // @[cache.scala 51:18 21:26]
  wire  _GEN_4692 = 2'h3 == state ? _GEN_3922 : valid_0_70; // @[cache.scala 51:18 21:26]
  wire  _GEN_4693 = 2'h3 == state ? _GEN_3923 : valid_0_71; // @[cache.scala 51:18 21:26]
  wire  _GEN_4694 = 2'h3 == state ? _GEN_3924 : valid_0_72; // @[cache.scala 51:18 21:26]
  wire  _GEN_4695 = 2'h3 == state ? _GEN_3925 : valid_0_73; // @[cache.scala 51:18 21:26]
  wire  _GEN_4696 = 2'h3 == state ? _GEN_3926 : valid_0_74; // @[cache.scala 51:18 21:26]
  wire  _GEN_4697 = 2'h3 == state ? _GEN_3927 : valid_0_75; // @[cache.scala 51:18 21:26]
  wire  _GEN_4698 = 2'h3 == state ? _GEN_3928 : valid_0_76; // @[cache.scala 51:18 21:26]
  wire  _GEN_4699 = 2'h3 == state ? _GEN_3929 : valid_0_77; // @[cache.scala 51:18 21:26]
  wire  _GEN_4700 = 2'h3 == state ? _GEN_3930 : valid_0_78; // @[cache.scala 51:18 21:26]
  wire  _GEN_4701 = 2'h3 == state ? _GEN_3931 : valid_0_79; // @[cache.scala 51:18 21:26]
  wire  _GEN_4702 = 2'h3 == state ? _GEN_3932 : valid_0_80; // @[cache.scala 51:18 21:26]
  wire  _GEN_4703 = 2'h3 == state ? _GEN_3933 : valid_0_81; // @[cache.scala 51:18 21:26]
  wire  _GEN_4704 = 2'h3 == state ? _GEN_3934 : valid_0_82; // @[cache.scala 51:18 21:26]
  wire  _GEN_4705 = 2'h3 == state ? _GEN_3935 : valid_0_83; // @[cache.scala 51:18 21:26]
  wire  _GEN_4706 = 2'h3 == state ? _GEN_3936 : valid_0_84; // @[cache.scala 51:18 21:26]
  wire  _GEN_4707 = 2'h3 == state ? _GEN_3937 : valid_0_85; // @[cache.scala 51:18 21:26]
  wire  _GEN_4708 = 2'h3 == state ? _GEN_3938 : valid_0_86; // @[cache.scala 51:18 21:26]
  wire  _GEN_4709 = 2'h3 == state ? _GEN_3939 : valid_0_87; // @[cache.scala 51:18 21:26]
  wire  _GEN_4710 = 2'h3 == state ? _GEN_3940 : valid_0_88; // @[cache.scala 51:18 21:26]
  wire  _GEN_4711 = 2'h3 == state ? _GEN_3941 : valid_0_89; // @[cache.scala 51:18 21:26]
  wire  _GEN_4712 = 2'h3 == state ? _GEN_3942 : valid_0_90; // @[cache.scala 51:18 21:26]
  wire  _GEN_4713 = 2'h3 == state ? _GEN_3943 : valid_0_91; // @[cache.scala 51:18 21:26]
  wire  _GEN_4714 = 2'h3 == state ? _GEN_3944 : valid_0_92; // @[cache.scala 51:18 21:26]
  wire  _GEN_4715 = 2'h3 == state ? _GEN_3945 : valid_0_93; // @[cache.scala 51:18 21:26]
  wire  _GEN_4716 = 2'h3 == state ? _GEN_3946 : valid_0_94; // @[cache.scala 51:18 21:26]
  wire  _GEN_4717 = 2'h3 == state ? _GEN_3947 : valid_0_95; // @[cache.scala 51:18 21:26]
  wire  _GEN_4718 = 2'h3 == state ? _GEN_3948 : valid_0_96; // @[cache.scala 51:18 21:26]
  wire  _GEN_4719 = 2'h3 == state ? _GEN_3949 : valid_0_97; // @[cache.scala 51:18 21:26]
  wire  _GEN_4720 = 2'h3 == state ? _GEN_3950 : valid_0_98; // @[cache.scala 51:18 21:26]
  wire  _GEN_4721 = 2'h3 == state ? _GEN_3951 : valid_0_99; // @[cache.scala 51:18 21:26]
  wire  _GEN_4722 = 2'h3 == state ? _GEN_3952 : valid_0_100; // @[cache.scala 51:18 21:26]
  wire  _GEN_4723 = 2'h3 == state ? _GEN_3953 : valid_0_101; // @[cache.scala 51:18 21:26]
  wire  _GEN_4724 = 2'h3 == state ? _GEN_3954 : valid_0_102; // @[cache.scala 51:18 21:26]
  wire  _GEN_4725 = 2'h3 == state ? _GEN_3955 : valid_0_103; // @[cache.scala 51:18 21:26]
  wire  _GEN_4726 = 2'h3 == state ? _GEN_3956 : valid_0_104; // @[cache.scala 51:18 21:26]
  wire  _GEN_4727 = 2'h3 == state ? _GEN_3957 : valid_0_105; // @[cache.scala 51:18 21:26]
  wire  _GEN_4728 = 2'h3 == state ? _GEN_3958 : valid_0_106; // @[cache.scala 51:18 21:26]
  wire  _GEN_4729 = 2'h3 == state ? _GEN_3959 : valid_0_107; // @[cache.scala 51:18 21:26]
  wire  _GEN_4730 = 2'h3 == state ? _GEN_3960 : valid_0_108; // @[cache.scala 51:18 21:26]
  wire  _GEN_4731 = 2'h3 == state ? _GEN_3961 : valid_0_109; // @[cache.scala 51:18 21:26]
  wire  _GEN_4732 = 2'h3 == state ? _GEN_3962 : valid_0_110; // @[cache.scala 51:18 21:26]
  wire  _GEN_4733 = 2'h3 == state ? _GEN_3963 : valid_0_111; // @[cache.scala 51:18 21:26]
  wire  _GEN_4734 = 2'h3 == state ? _GEN_3964 : valid_0_112; // @[cache.scala 51:18 21:26]
  wire  _GEN_4735 = 2'h3 == state ? _GEN_3965 : valid_0_113; // @[cache.scala 51:18 21:26]
  wire  _GEN_4736 = 2'h3 == state ? _GEN_3966 : valid_0_114; // @[cache.scala 51:18 21:26]
  wire  _GEN_4737 = 2'h3 == state ? _GEN_3967 : valid_0_115; // @[cache.scala 51:18 21:26]
  wire  _GEN_4738 = 2'h3 == state ? _GEN_3968 : valid_0_116; // @[cache.scala 51:18 21:26]
  wire  _GEN_4739 = 2'h3 == state ? _GEN_3969 : valid_0_117; // @[cache.scala 51:18 21:26]
  wire  _GEN_4740 = 2'h3 == state ? _GEN_3970 : valid_0_118; // @[cache.scala 51:18 21:26]
  wire  _GEN_4741 = 2'h3 == state ? _GEN_3971 : valid_0_119; // @[cache.scala 51:18 21:26]
  wire  _GEN_4742 = 2'h3 == state ? _GEN_3972 : valid_0_120; // @[cache.scala 51:18 21:26]
  wire  _GEN_4743 = 2'h3 == state ? _GEN_3973 : valid_0_121; // @[cache.scala 51:18 21:26]
  wire  _GEN_4744 = 2'h3 == state ? _GEN_3974 : valid_0_122; // @[cache.scala 51:18 21:26]
  wire  _GEN_4745 = 2'h3 == state ? _GEN_3975 : valid_0_123; // @[cache.scala 51:18 21:26]
  wire  _GEN_4746 = 2'h3 == state ? _GEN_3976 : valid_0_124; // @[cache.scala 51:18 21:26]
  wire  _GEN_4747 = 2'h3 == state ? _GEN_3977 : valid_0_125; // @[cache.scala 51:18 21:26]
  wire  _GEN_4748 = 2'h3 == state ? _GEN_3978 : valid_0_126; // @[cache.scala 51:18 21:26]
  wire  _GEN_4749 = 2'h3 == state ? _GEN_3979 : valid_0_127; // @[cache.scala 51:18 21:26]
  wire  _GEN_4750 = 2'h3 == state ? _GEN_3980 : quene; // @[cache.scala 51:18 28:24]
  wire [63:0] _GEN_4751 = 2'h3 == state ? _GEN_3981 : ram_1_0; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4752 = 2'h3 == state ? _GEN_3982 : ram_1_1; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4753 = 2'h3 == state ? _GEN_3983 : ram_1_2; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4754 = 2'h3 == state ? _GEN_3984 : ram_1_3; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4755 = 2'h3 == state ? _GEN_3985 : ram_1_4; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4756 = 2'h3 == state ? _GEN_3986 : ram_1_5; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4757 = 2'h3 == state ? _GEN_3987 : ram_1_6; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4758 = 2'h3 == state ? _GEN_3988 : ram_1_7; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4759 = 2'h3 == state ? _GEN_3989 : ram_1_8; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4760 = 2'h3 == state ? _GEN_3990 : ram_1_9; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4761 = 2'h3 == state ? _GEN_3991 : ram_1_10; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4762 = 2'h3 == state ? _GEN_3992 : ram_1_11; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4763 = 2'h3 == state ? _GEN_3993 : ram_1_12; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4764 = 2'h3 == state ? _GEN_3994 : ram_1_13; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4765 = 2'h3 == state ? _GEN_3995 : ram_1_14; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4766 = 2'h3 == state ? _GEN_3996 : ram_1_15; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4767 = 2'h3 == state ? _GEN_3997 : ram_1_16; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4768 = 2'h3 == state ? _GEN_3998 : ram_1_17; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4769 = 2'h3 == state ? _GEN_3999 : ram_1_18; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4770 = 2'h3 == state ? _GEN_4000 : ram_1_19; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4771 = 2'h3 == state ? _GEN_4001 : ram_1_20; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4772 = 2'h3 == state ? _GEN_4002 : ram_1_21; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4773 = 2'h3 == state ? _GEN_4003 : ram_1_22; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4774 = 2'h3 == state ? _GEN_4004 : ram_1_23; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4775 = 2'h3 == state ? _GEN_4005 : ram_1_24; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4776 = 2'h3 == state ? _GEN_4006 : ram_1_25; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4777 = 2'h3 == state ? _GEN_4007 : ram_1_26; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4778 = 2'h3 == state ? _GEN_4008 : ram_1_27; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4779 = 2'h3 == state ? _GEN_4009 : ram_1_28; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4780 = 2'h3 == state ? _GEN_4010 : ram_1_29; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4781 = 2'h3 == state ? _GEN_4011 : ram_1_30; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4782 = 2'h3 == state ? _GEN_4012 : ram_1_31; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4783 = 2'h3 == state ? _GEN_4013 : ram_1_32; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4784 = 2'h3 == state ? _GEN_4014 : ram_1_33; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4785 = 2'h3 == state ? _GEN_4015 : ram_1_34; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4786 = 2'h3 == state ? _GEN_4016 : ram_1_35; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4787 = 2'h3 == state ? _GEN_4017 : ram_1_36; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4788 = 2'h3 == state ? _GEN_4018 : ram_1_37; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4789 = 2'h3 == state ? _GEN_4019 : ram_1_38; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4790 = 2'h3 == state ? _GEN_4020 : ram_1_39; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4791 = 2'h3 == state ? _GEN_4021 : ram_1_40; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4792 = 2'h3 == state ? _GEN_4022 : ram_1_41; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4793 = 2'h3 == state ? _GEN_4023 : ram_1_42; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4794 = 2'h3 == state ? _GEN_4024 : ram_1_43; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4795 = 2'h3 == state ? _GEN_4025 : ram_1_44; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4796 = 2'h3 == state ? _GEN_4026 : ram_1_45; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4797 = 2'h3 == state ? _GEN_4027 : ram_1_46; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4798 = 2'h3 == state ? _GEN_4028 : ram_1_47; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4799 = 2'h3 == state ? _GEN_4029 : ram_1_48; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4800 = 2'h3 == state ? _GEN_4030 : ram_1_49; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4801 = 2'h3 == state ? _GEN_4031 : ram_1_50; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4802 = 2'h3 == state ? _GEN_4032 : ram_1_51; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4803 = 2'h3 == state ? _GEN_4033 : ram_1_52; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4804 = 2'h3 == state ? _GEN_4034 : ram_1_53; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4805 = 2'h3 == state ? _GEN_4035 : ram_1_54; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4806 = 2'h3 == state ? _GEN_4036 : ram_1_55; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4807 = 2'h3 == state ? _GEN_4037 : ram_1_56; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4808 = 2'h3 == state ? _GEN_4038 : ram_1_57; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4809 = 2'h3 == state ? _GEN_4039 : ram_1_58; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4810 = 2'h3 == state ? _GEN_4040 : ram_1_59; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4811 = 2'h3 == state ? _GEN_4041 : ram_1_60; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4812 = 2'h3 == state ? _GEN_4042 : ram_1_61; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4813 = 2'h3 == state ? _GEN_4043 : ram_1_62; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4814 = 2'h3 == state ? _GEN_4044 : ram_1_63; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4815 = 2'h3 == state ? _GEN_4045 : ram_1_64; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4816 = 2'h3 == state ? _GEN_4046 : ram_1_65; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4817 = 2'h3 == state ? _GEN_4047 : ram_1_66; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4818 = 2'h3 == state ? _GEN_4048 : ram_1_67; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4819 = 2'h3 == state ? _GEN_4049 : ram_1_68; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4820 = 2'h3 == state ? _GEN_4050 : ram_1_69; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4821 = 2'h3 == state ? _GEN_4051 : ram_1_70; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4822 = 2'h3 == state ? _GEN_4052 : ram_1_71; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4823 = 2'h3 == state ? _GEN_4053 : ram_1_72; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4824 = 2'h3 == state ? _GEN_4054 : ram_1_73; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4825 = 2'h3 == state ? _GEN_4055 : ram_1_74; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4826 = 2'h3 == state ? _GEN_4056 : ram_1_75; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4827 = 2'h3 == state ? _GEN_4057 : ram_1_76; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4828 = 2'h3 == state ? _GEN_4058 : ram_1_77; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4829 = 2'h3 == state ? _GEN_4059 : ram_1_78; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4830 = 2'h3 == state ? _GEN_4060 : ram_1_79; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4831 = 2'h3 == state ? _GEN_4061 : ram_1_80; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4832 = 2'h3 == state ? _GEN_4062 : ram_1_81; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4833 = 2'h3 == state ? _GEN_4063 : ram_1_82; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4834 = 2'h3 == state ? _GEN_4064 : ram_1_83; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4835 = 2'h3 == state ? _GEN_4065 : ram_1_84; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4836 = 2'h3 == state ? _GEN_4066 : ram_1_85; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4837 = 2'h3 == state ? _GEN_4067 : ram_1_86; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4838 = 2'h3 == state ? _GEN_4068 : ram_1_87; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4839 = 2'h3 == state ? _GEN_4069 : ram_1_88; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4840 = 2'h3 == state ? _GEN_4070 : ram_1_89; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4841 = 2'h3 == state ? _GEN_4071 : ram_1_90; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4842 = 2'h3 == state ? _GEN_4072 : ram_1_91; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4843 = 2'h3 == state ? _GEN_4073 : ram_1_92; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4844 = 2'h3 == state ? _GEN_4074 : ram_1_93; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4845 = 2'h3 == state ? _GEN_4075 : ram_1_94; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4846 = 2'h3 == state ? _GEN_4076 : ram_1_95; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4847 = 2'h3 == state ? _GEN_4077 : ram_1_96; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4848 = 2'h3 == state ? _GEN_4078 : ram_1_97; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4849 = 2'h3 == state ? _GEN_4079 : ram_1_98; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4850 = 2'h3 == state ? _GEN_4080 : ram_1_99; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4851 = 2'h3 == state ? _GEN_4081 : ram_1_100; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4852 = 2'h3 == state ? _GEN_4082 : ram_1_101; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4853 = 2'h3 == state ? _GEN_4083 : ram_1_102; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4854 = 2'h3 == state ? _GEN_4084 : ram_1_103; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4855 = 2'h3 == state ? _GEN_4085 : ram_1_104; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4856 = 2'h3 == state ? _GEN_4086 : ram_1_105; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4857 = 2'h3 == state ? _GEN_4087 : ram_1_106; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4858 = 2'h3 == state ? _GEN_4088 : ram_1_107; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4859 = 2'h3 == state ? _GEN_4089 : ram_1_108; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4860 = 2'h3 == state ? _GEN_4090 : ram_1_109; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4861 = 2'h3 == state ? _GEN_4091 : ram_1_110; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4862 = 2'h3 == state ? _GEN_4092 : ram_1_111; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4863 = 2'h3 == state ? _GEN_4093 : ram_1_112; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4864 = 2'h3 == state ? _GEN_4094 : ram_1_113; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4865 = 2'h3 == state ? _GEN_4095 : ram_1_114; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4866 = 2'h3 == state ? _GEN_4096 : ram_1_115; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4867 = 2'h3 == state ? _GEN_4097 : ram_1_116; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4868 = 2'h3 == state ? _GEN_4098 : ram_1_117; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4869 = 2'h3 == state ? _GEN_4099 : ram_1_118; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4870 = 2'h3 == state ? _GEN_4100 : ram_1_119; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4871 = 2'h3 == state ? _GEN_4101 : ram_1_120; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4872 = 2'h3 == state ? _GEN_4102 : ram_1_121; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4873 = 2'h3 == state ? _GEN_4103 : ram_1_122; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4874 = 2'h3 == state ? _GEN_4104 : ram_1_123; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4875 = 2'h3 == state ? _GEN_4105 : ram_1_124; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4876 = 2'h3 == state ? _GEN_4106 : ram_1_125; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4877 = 2'h3 == state ? _GEN_4107 : ram_1_126; // @[cache.scala 51:18 18:24]
  wire [63:0] _GEN_4878 = 2'h3 == state ? _GEN_4108 : ram_1_127; // @[cache.scala 51:18 18:24]
  wire [31:0] _GEN_4879 = 2'h3 == state ? _GEN_4109 : tag_1_0; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4880 = 2'h3 == state ? _GEN_4110 : tag_1_1; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4881 = 2'h3 == state ? _GEN_4111 : tag_1_2; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4882 = 2'h3 == state ? _GEN_4112 : tag_1_3; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4883 = 2'h3 == state ? _GEN_4113 : tag_1_4; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4884 = 2'h3 == state ? _GEN_4114 : tag_1_5; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4885 = 2'h3 == state ? _GEN_4115 : tag_1_6; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4886 = 2'h3 == state ? _GEN_4116 : tag_1_7; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4887 = 2'h3 == state ? _GEN_4117 : tag_1_8; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4888 = 2'h3 == state ? _GEN_4118 : tag_1_9; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4889 = 2'h3 == state ? _GEN_4119 : tag_1_10; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4890 = 2'h3 == state ? _GEN_4120 : tag_1_11; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4891 = 2'h3 == state ? _GEN_4121 : tag_1_12; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4892 = 2'h3 == state ? _GEN_4122 : tag_1_13; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4893 = 2'h3 == state ? _GEN_4123 : tag_1_14; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4894 = 2'h3 == state ? _GEN_4124 : tag_1_15; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4895 = 2'h3 == state ? _GEN_4125 : tag_1_16; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4896 = 2'h3 == state ? _GEN_4126 : tag_1_17; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4897 = 2'h3 == state ? _GEN_4127 : tag_1_18; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4898 = 2'h3 == state ? _GEN_4128 : tag_1_19; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4899 = 2'h3 == state ? _GEN_4129 : tag_1_20; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4900 = 2'h3 == state ? _GEN_4130 : tag_1_21; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4901 = 2'h3 == state ? _GEN_4131 : tag_1_22; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4902 = 2'h3 == state ? _GEN_4132 : tag_1_23; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4903 = 2'h3 == state ? _GEN_4133 : tag_1_24; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4904 = 2'h3 == state ? _GEN_4134 : tag_1_25; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4905 = 2'h3 == state ? _GEN_4135 : tag_1_26; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4906 = 2'h3 == state ? _GEN_4136 : tag_1_27; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4907 = 2'h3 == state ? _GEN_4137 : tag_1_28; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4908 = 2'h3 == state ? _GEN_4138 : tag_1_29; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4909 = 2'h3 == state ? _GEN_4139 : tag_1_30; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4910 = 2'h3 == state ? _GEN_4140 : tag_1_31; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4911 = 2'h3 == state ? _GEN_4141 : tag_1_32; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4912 = 2'h3 == state ? _GEN_4142 : tag_1_33; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4913 = 2'h3 == state ? _GEN_4143 : tag_1_34; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4914 = 2'h3 == state ? _GEN_4144 : tag_1_35; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4915 = 2'h3 == state ? _GEN_4145 : tag_1_36; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4916 = 2'h3 == state ? _GEN_4146 : tag_1_37; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4917 = 2'h3 == state ? _GEN_4147 : tag_1_38; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4918 = 2'h3 == state ? _GEN_4148 : tag_1_39; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4919 = 2'h3 == state ? _GEN_4149 : tag_1_40; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4920 = 2'h3 == state ? _GEN_4150 : tag_1_41; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4921 = 2'h3 == state ? _GEN_4151 : tag_1_42; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4922 = 2'h3 == state ? _GEN_4152 : tag_1_43; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4923 = 2'h3 == state ? _GEN_4153 : tag_1_44; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4924 = 2'h3 == state ? _GEN_4154 : tag_1_45; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4925 = 2'h3 == state ? _GEN_4155 : tag_1_46; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4926 = 2'h3 == state ? _GEN_4156 : tag_1_47; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4927 = 2'h3 == state ? _GEN_4157 : tag_1_48; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4928 = 2'h3 == state ? _GEN_4158 : tag_1_49; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4929 = 2'h3 == state ? _GEN_4159 : tag_1_50; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4930 = 2'h3 == state ? _GEN_4160 : tag_1_51; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4931 = 2'h3 == state ? _GEN_4161 : tag_1_52; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4932 = 2'h3 == state ? _GEN_4162 : tag_1_53; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4933 = 2'h3 == state ? _GEN_4163 : tag_1_54; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4934 = 2'h3 == state ? _GEN_4164 : tag_1_55; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4935 = 2'h3 == state ? _GEN_4165 : tag_1_56; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4936 = 2'h3 == state ? _GEN_4166 : tag_1_57; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4937 = 2'h3 == state ? _GEN_4167 : tag_1_58; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4938 = 2'h3 == state ? _GEN_4168 : tag_1_59; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4939 = 2'h3 == state ? _GEN_4169 : tag_1_60; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4940 = 2'h3 == state ? _GEN_4170 : tag_1_61; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4941 = 2'h3 == state ? _GEN_4171 : tag_1_62; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4942 = 2'h3 == state ? _GEN_4172 : tag_1_63; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4943 = 2'h3 == state ? _GEN_4173 : tag_1_64; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4944 = 2'h3 == state ? _GEN_4174 : tag_1_65; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4945 = 2'h3 == state ? _GEN_4175 : tag_1_66; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4946 = 2'h3 == state ? _GEN_4176 : tag_1_67; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4947 = 2'h3 == state ? _GEN_4177 : tag_1_68; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4948 = 2'h3 == state ? _GEN_4178 : tag_1_69; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4949 = 2'h3 == state ? _GEN_4179 : tag_1_70; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4950 = 2'h3 == state ? _GEN_4180 : tag_1_71; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4951 = 2'h3 == state ? _GEN_4181 : tag_1_72; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4952 = 2'h3 == state ? _GEN_4182 : tag_1_73; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4953 = 2'h3 == state ? _GEN_4183 : tag_1_74; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4954 = 2'h3 == state ? _GEN_4184 : tag_1_75; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4955 = 2'h3 == state ? _GEN_4185 : tag_1_76; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4956 = 2'h3 == state ? _GEN_4186 : tag_1_77; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4957 = 2'h3 == state ? _GEN_4187 : tag_1_78; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4958 = 2'h3 == state ? _GEN_4188 : tag_1_79; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4959 = 2'h3 == state ? _GEN_4189 : tag_1_80; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4960 = 2'h3 == state ? _GEN_4190 : tag_1_81; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4961 = 2'h3 == state ? _GEN_4191 : tag_1_82; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4962 = 2'h3 == state ? _GEN_4192 : tag_1_83; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4963 = 2'h3 == state ? _GEN_4193 : tag_1_84; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4964 = 2'h3 == state ? _GEN_4194 : tag_1_85; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4965 = 2'h3 == state ? _GEN_4195 : tag_1_86; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4966 = 2'h3 == state ? _GEN_4196 : tag_1_87; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4967 = 2'h3 == state ? _GEN_4197 : tag_1_88; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4968 = 2'h3 == state ? _GEN_4198 : tag_1_89; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4969 = 2'h3 == state ? _GEN_4199 : tag_1_90; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4970 = 2'h3 == state ? _GEN_4200 : tag_1_91; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4971 = 2'h3 == state ? _GEN_4201 : tag_1_92; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4972 = 2'h3 == state ? _GEN_4202 : tag_1_93; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4973 = 2'h3 == state ? _GEN_4203 : tag_1_94; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4974 = 2'h3 == state ? _GEN_4204 : tag_1_95; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4975 = 2'h3 == state ? _GEN_4205 : tag_1_96; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4976 = 2'h3 == state ? _GEN_4206 : tag_1_97; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4977 = 2'h3 == state ? _GEN_4207 : tag_1_98; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4978 = 2'h3 == state ? _GEN_4208 : tag_1_99; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4979 = 2'h3 == state ? _GEN_4209 : tag_1_100; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4980 = 2'h3 == state ? _GEN_4210 : tag_1_101; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4981 = 2'h3 == state ? _GEN_4211 : tag_1_102; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4982 = 2'h3 == state ? _GEN_4212 : tag_1_103; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4983 = 2'h3 == state ? _GEN_4213 : tag_1_104; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4984 = 2'h3 == state ? _GEN_4214 : tag_1_105; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4985 = 2'h3 == state ? _GEN_4215 : tag_1_106; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4986 = 2'h3 == state ? _GEN_4216 : tag_1_107; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4987 = 2'h3 == state ? _GEN_4217 : tag_1_108; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4988 = 2'h3 == state ? _GEN_4218 : tag_1_109; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4989 = 2'h3 == state ? _GEN_4219 : tag_1_110; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4990 = 2'h3 == state ? _GEN_4220 : tag_1_111; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4991 = 2'h3 == state ? _GEN_4221 : tag_1_112; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4992 = 2'h3 == state ? _GEN_4222 : tag_1_113; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4993 = 2'h3 == state ? _GEN_4223 : tag_1_114; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4994 = 2'h3 == state ? _GEN_4224 : tag_1_115; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4995 = 2'h3 == state ? _GEN_4225 : tag_1_116; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4996 = 2'h3 == state ? _GEN_4226 : tag_1_117; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4997 = 2'h3 == state ? _GEN_4227 : tag_1_118; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4998 = 2'h3 == state ? _GEN_4228 : tag_1_119; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_4999 = 2'h3 == state ? _GEN_4229 : tag_1_120; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_5000 = 2'h3 == state ? _GEN_4230 : tag_1_121; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_5001 = 2'h3 == state ? _GEN_4231 : tag_1_122; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_5002 = 2'h3 == state ? _GEN_4232 : tag_1_123; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_5003 = 2'h3 == state ? _GEN_4233 : tag_1_124; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_5004 = 2'h3 == state ? _GEN_4234 : tag_1_125; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_5005 = 2'h3 == state ? _GEN_4235 : tag_1_126; // @[cache.scala 51:18 20:24]
  wire [31:0] _GEN_5006 = 2'h3 == state ? _GEN_4236 : tag_1_127; // @[cache.scala 51:18 20:24]
  wire  _GEN_5007 = 2'h3 == state ? _GEN_4237 : valid_1_0; // @[cache.scala 51:18 22:26]
  wire  _GEN_5008 = 2'h3 == state ? _GEN_4238 : valid_1_1; // @[cache.scala 51:18 22:26]
  wire  _GEN_5009 = 2'h3 == state ? _GEN_4239 : valid_1_2; // @[cache.scala 51:18 22:26]
  wire  _GEN_5010 = 2'h3 == state ? _GEN_4240 : valid_1_3; // @[cache.scala 51:18 22:26]
  wire  _GEN_5011 = 2'h3 == state ? _GEN_4241 : valid_1_4; // @[cache.scala 51:18 22:26]
  wire  _GEN_5012 = 2'h3 == state ? _GEN_4242 : valid_1_5; // @[cache.scala 51:18 22:26]
  wire  _GEN_5013 = 2'h3 == state ? _GEN_4243 : valid_1_6; // @[cache.scala 51:18 22:26]
  wire  _GEN_5014 = 2'h3 == state ? _GEN_4244 : valid_1_7; // @[cache.scala 51:18 22:26]
  wire  _GEN_5015 = 2'h3 == state ? _GEN_4245 : valid_1_8; // @[cache.scala 51:18 22:26]
  wire  _GEN_5016 = 2'h3 == state ? _GEN_4246 : valid_1_9; // @[cache.scala 51:18 22:26]
  wire  _GEN_5017 = 2'h3 == state ? _GEN_4247 : valid_1_10; // @[cache.scala 51:18 22:26]
  wire  _GEN_5018 = 2'h3 == state ? _GEN_4248 : valid_1_11; // @[cache.scala 51:18 22:26]
  wire  _GEN_5019 = 2'h3 == state ? _GEN_4249 : valid_1_12; // @[cache.scala 51:18 22:26]
  wire  _GEN_5020 = 2'h3 == state ? _GEN_4250 : valid_1_13; // @[cache.scala 51:18 22:26]
  wire  _GEN_5021 = 2'h3 == state ? _GEN_4251 : valid_1_14; // @[cache.scala 51:18 22:26]
  wire  _GEN_5022 = 2'h3 == state ? _GEN_4252 : valid_1_15; // @[cache.scala 51:18 22:26]
  wire  _GEN_5023 = 2'h3 == state ? _GEN_4253 : valid_1_16; // @[cache.scala 51:18 22:26]
  wire  _GEN_5024 = 2'h3 == state ? _GEN_4254 : valid_1_17; // @[cache.scala 51:18 22:26]
  wire  _GEN_5025 = 2'h3 == state ? _GEN_4255 : valid_1_18; // @[cache.scala 51:18 22:26]
  wire  _GEN_5026 = 2'h3 == state ? _GEN_4256 : valid_1_19; // @[cache.scala 51:18 22:26]
  wire  _GEN_5027 = 2'h3 == state ? _GEN_4257 : valid_1_20; // @[cache.scala 51:18 22:26]
  wire  _GEN_5028 = 2'h3 == state ? _GEN_4258 : valid_1_21; // @[cache.scala 51:18 22:26]
  wire  _GEN_5029 = 2'h3 == state ? _GEN_4259 : valid_1_22; // @[cache.scala 51:18 22:26]
  wire  _GEN_5030 = 2'h3 == state ? _GEN_4260 : valid_1_23; // @[cache.scala 51:18 22:26]
  wire  _GEN_5031 = 2'h3 == state ? _GEN_4261 : valid_1_24; // @[cache.scala 51:18 22:26]
  wire  _GEN_5032 = 2'h3 == state ? _GEN_4262 : valid_1_25; // @[cache.scala 51:18 22:26]
  wire  _GEN_5033 = 2'h3 == state ? _GEN_4263 : valid_1_26; // @[cache.scala 51:18 22:26]
  wire  _GEN_5034 = 2'h3 == state ? _GEN_4264 : valid_1_27; // @[cache.scala 51:18 22:26]
  wire  _GEN_5035 = 2'h3 == state ? _GEN_4265 : valid_1_28; // @[cache.scala 51:18 22:26]
  wire  _GEN_5036 = 2'h3 == state ? _GEN_4266 : valid_1_29; // @[cache.scala 51:18 22:26]
  wire  _GEN_5037 = 2'h3 == state ? _GEN_4267 : valid_1_30; // @[cache.scala 51:18 22:26]
  wire  _GEN_5038 = 2'h3 == state ? _GEN_4268 : valid_1_31; // @[cache.scala 51:18 22:26]
  wire  _GEN_5039 = 2'h3 == state ? _GEN_4269 : valid_1_32; // @[cache.scala 51:18 22:26]
  wire  _GEN_5040 = 2'h3 == state ? _GEN_4270 : valid_1_33; // @[cache.scala 51:18 22:26]
  wire  _GEN_5041 = 2'h3 == state ? _GEN_4271 : valid_1_34; // @[cache.scala 51:18 22:26]
  wire  _GEN_5042 = 2'h3 == state ? _GEN_4272 : valid_1_35; // @[cache.scala 51:18 22:26]
  wire  _GEN_5043 = 2'h3 == state ? _GEN_4273 : valid_1_36; // @[cache.scala 51:18 22:26]
  wire  _GEN_5044 = 2'h3 == state ? _GEN_4274 : valid_1_37; // @[cache.scala 51:18 22:26]
  wire  _GEN_5045 = 2'h3 == state ? _GEN_4275 : valid_1_38; // @[cache.scala 51:18 22:26]
  wire  _GEN_5046 = 2'h3 == state ? _GEN_4276 : valid_1_39; // @[cache.scala 51:18 22:26]
  wire  _GEN_5047 = 2'h3 == state ? _GEN_4277 : valid_1_40; // @[cache.scala 51:18 22:26]
  wire  _GEN_5048 = 2'h3 == state ? _GEN_4278 : valid_1_41; // @[cache.scala 51:18 22:26]
  wire  _GEN_5049 = 2'h3 == state ? _GEN_4279 : valid_1_42; // @[cache.scala 51:18 22:26]
  wire  _GEN_5050 = 2'h3 == state ? _GEN_4280 : valid_1_43; // @[cache.scala 51:18 22:26]
  wire  _GEN_5051 = 2'h3 == state ? _GEN_4281 : valid_1_44; // @[cache.scala 51:18 22:26]
  wire  _GEN_5052 = 2'h3 == state ? _GEN_4282 : valid_1_45; // @[cache.scala 51:18 22:26]
  wire  _GEN_5053 = 2'h3 == state ? _GEN_4283 : valid_1_46; // @[cache.scala 51:18 22:26]
  wire  _GEN_5054 = 2'h3 == state ? _GEN_4284 : valid_1_47; // @[cache.scala 51:18 22:26]
  wire  _GEN_5055 = 2'h3 == state ? _GEN_4285 : valid_1_48; // @[cache.scala 51:18 22:26]
  wire  _GEN_5056 = 2'h3 == state ? _GEN_4286 : valid_1_49; // @[cache.scala 51:18 22:26]
  wire  _GEN_5057 = 2'h3 == state ? _GEN_4287 : valid_1_50; // @[cache.scala 51:18 22:26]
  wire  _GEN_5058 = 2'h3 == state ? _GEN_4288 : valid_1_51; // @[cache.scala 51:18 22:26]
  wire  _GEN_5059 = 2'h3 == state ? _GEN_4289 : valid_1_52; // @[cache.scala 51:18 22:26]
  wire  _GEN_5060 = 2'h3 == state ? _GEN_4290 : valid_1_53; // @[cache.scala 51:18 22:26]
  wire  _GEN_5061 = 2'h3 == state ? _GEN_4291 : valid_1_54; // @[cache.scala 51:18 22:26]
  wire  _GEN_5062 = 2'h3 == state ? _GEN_4292 : valid_1_55; // @[cache.scala 51:18 22:26]
  wire  _GEN_5063 = 2'h3 == state ? _GEN_4293 : valid_1_56; // @[cache.scala 51:18 22:26]
  wire  _GEN_5064 = 2'h3 == state ? _GEN_4294 : valid_1_57; // @[cache.scala 51:18 22:26]
  wire  _GEN_5065 = 2'h3 == state ? _GEN_4295 : valid_1_58; // @[cache.scala 51:18 22:26]
  wire  _GEN_5066 = 2'h3 == state ? _GEN_4296 : valid_1_59; // @[cache.scala 51:18 22:26]
  wire  _GEN_5067 = 2'h3 == state ? _GEN_4297 : valid_1_60; // @[cache.scala 51:18 22:26]
  wire  _GEN_5068 = 2'h3 == state ? _GEN_4298 : valid_1_61; // @[cache.scala 51:18 22:26]
  wire  _GEN_5069 = 2'h3 == state ? _GEN_4299 : valid_1_62; // @[cache.scala 51:18 22:26]
  wire  _GEN_5070 = 2'h3 == state ? _GEN_4300 : valid_1_63; // @[cache.scala 51:18 22:26]
  wire  _GEN_5071 = 2'h3 == state ? _GEN_4301 : valid_1_64; // @[cache.scala 51:18 22:26]
  wire  _GEN_5072 = 2'h3 == state ? _GEN_4302 : valid_1_65; // @[cache.scala 51:18 22:26]
  wire  _GEN_5073 = 2'h3 == state ? _GEN_4303 : valid_1_66; // @[cache.scala 51:18 22:26]
  wire  _GEN_5074 = 2'h3 == state ? _GEN_4304 : valid_1_67; // @[cache.scala 51:18 22:26]
  wire  _GEN_5075 = 2'h3 == state ? _GEN_4305 : valid_1_68; // @[cache.scala 51:18 22:26]
  wire  _GEN_5076 = 2'h3 == state ? _GEN_4306 : valid_1_69; // @[cache.scala 51:18 22:26]
  wire  _GEN_5077 = 2'h3 == state ? _GEN_4307 : valid_1_70; // @[cache.scala 51:18 22:26]
  wire  _GEN_5078 = 2'h3 == state ? _GEN_4308 : valid_1_71; // @[cache.scala 51:18 22:26]
  wire  _GEN_5079 = 2'h3 == state ? _GEN_4309 : valid_1_72; // @[cache.scala 51:18 22:26]
  wire  _GEN_5080 = 2'h3 == state ? _GEN_4310 : valid_1_73; // @[cache.scala 51:18 22:26]
  wire  _GEN_5081 = 2'h3 == state ? _GEN_4311 : valid_1_74; // @[cache.scala 51:18 22:26]
  wire  _GEN_5082 = 2'h3 == state ? _GEN_4312 : valid_1_75; // @[cache.scala 51:18 22:26]
  wire  _GEN_5083 = 2'h3 == state ? _GEN_4313 : valid_1_76; // @[cache.scala 51:18 22:26]
  wire  _GEN_5084 = 2'h3 == state ? _GEN_4314 : valid_1_77; // @[cache.scala 51:18 22:26]
  wire  _GEN_5085 = 2'h3 == state ? _GEN_4315 : valid_1_78; // @[cache.scala 51:18 22:26]
  wire  _GEN_5086 = 2'h3 == state ? _GEN_4316 : valid_1_79; // @[cache.scala 51:18 22:26]
  wire  _GEN_5087 = 2'h3 == state ? _GEN_4317 : valid_1_80; // @[cache.scala 51:18 22:26]
  wire  _GEN_5088 = 2'h3 == state ? _GEN_4318 : valid_1_81; // @[cache.scala 51:18 22:26]
  wire  _GEN_5089 = 2'h3 == state ? _GEN_4319 : valid_1_82; // @[cache.scala 51:18 22:26]
  wire  _GEN_5090 = 2'h3 == state ? _GEN_4320 : valid_1_83; // @[cache.scala 51:18 22:26]
  wire  _GEN_5091 = 2'h3 == state ? _GEN_4321 : valid_1_84; // @[cache.scala 51:18 22:26]
  wire  _GEN_5092 = 2'h3 == state ? _GEN_4322 : valid_1_85; // @[cache.scala 51:18 22:26]
  wire  _GEN_5093 = 2'h3 == state ? _GEN_4323 : valid_1_86; // @[cache.scala 51:18 22:26]
  wire  _GEN_5094 = 2'h3 == state ? _GEN_4324 : valid_1_87; // @[cache.scala 51:18 22:26]
  wire  _GEN_5095 = 2'h3 == state ? _GEN_4325 : valid_1_88; // @[cache.scala 51:18 22:26]
  wire  _GEN_5096 = 2'h3 == state ? _GEN_4326 : valid_1_89; // @[cache.scala 51:18 22:26]
  wire  _GEN_5097 = 2'h3 == state ? _GEN_4327 : valid_1_90; // @[cache.scala 51:18 22:26]
  wire  _GEN_5098 = 2'h3 == state ? _GEN_4328 : valid_1_91; // @[cache.scala 51:18 22:26]
  wire  _GEN_5099 = 2'h3 == state ? _GEN_4329 : valid_1_92; // @[cache.scala 51:18 22:26]
  wire  _GEN_5100 = 2'h3 == state ? _GEN_4330 : valid_1_93; // @[cache.scala 51:18 22:26]
  wire  _GEN_5101 = 2'h3 == state ? _GEN_4331 : valid_1_94; // @[cache.scala 51:18 22:26]
  wire  _GEN_5102 = 2'h3 == state ? _GEN_4332 : valid_1_95; // @[cache.scala 51:18 22:26]
  wire  _GEN_5103 = 2'h3 == state ? _GEN_4333 : valid_1_96; // @[cache.scala 51:18 22:26]
  wire  _GEN_5104 = 2'h3 == state ? _GEN_4334 : valid_1_97; // @[cache.scala 51:18 22:26]
  wire  _GEN_5105 = 2'h3 == state ? _GEN_4335 : valid_1_98; // @[cache.scala 51:18 22:26]
  wire  _GEN_5106 = 2'h3 == state ? _GEN_4336 : valid_1_99; // @[cache.scala 51:18 22:26]
  wire  _GEN_5107 = 2'h3 == state ? _GEN_4337 : valid_1_100; // @[cache.scala 51:18 22:26]
  wire  _GEN_5108 = 2'h3 == state ? _GEN_4338 : valid_1_101; // @[cache.scala 51:18 22:26]
  wire  _GEN_5109 = 2'h3 == state ? _GEN_4339 : valid_1_102; // @[cache.scala 51:18 22:26]
  wire  _GEN_5110 = 2'h3 == state ? _GEN_4340 : valid_1_103; // @[cache.scala 51:18 22:26]
  wire  _GEN_5111 = 2'h3 == state ? _GEN_4341 : valid_1_104; // @[cache.scala 51:18 22:26]
  wire  _GEN_5112 = 2'h3 == state ? _GEN_4342 : valid_1_105; // @[cache.scala 51:18 22:26]
  wire  _GEN_5113 = 2'h3 == state ? _GEN_4343 : valid_1_106; // @[cache.scala 51:18 22:26]
  wire  _GEN_5114 = 2'h3 == state ? _GEN_4344 : valid_1_107; // @[cache.scala 51:18 22:26]
  wire  _GEN_5115 = 2'h3 == state ? _GEN_4345 : valid_1_108; // @[cache.scala 51:18 22:26]
  wire  _GEN_5116 = 2'h3 == state ? _GEN_4346 : valid_1_109; // @[cache.scala 51:18 22:26]
  wire  _GEN_5117 = 2'h3 == state ? _GEN_4347 : valid_1_110; // @[cache.scala 51:18 22:26]
  wire  _GEN_5118 = 2'h3 == state ? _GEN_4348 : valid_1_111; // @[cache.scala 51:18 22:26]
  wire  _GEN_5119 = 2'h3 == state ? _GEN_4349 : valid_1_112; // @[cache.scala 51:18 22:26]
  wire  _GEN_5120 = 2'h3 == state ? _GEN_4350 : valid_1_113; // @[cache.scala 51:18 22:26]
  wire  _GEN_5121 = 2'h3 == state ? _GEN_4351 : valid_1_114; // @[cache.scala 51:18 22:26]
  wire  _GEN_5122 = 2'h3 == state ? _GEN_4352 : valid_1_115; // @[cache.scala 51:18 22:26]
  wire  _GEN_5123 = 2'h3 == state ? _GEN_4353 : valid_1_116; // @[cache.scala 51:18 22:26]
  wire  _GEN_5124 = 2'h3 == state ? _GEN_4354 : valid_1_117; // @[cache.scala 51:18 22:26]
  wire  _GEN_5125 = 2'h3 == state ? _GEN_4355 : valid_1_118; // @[cache.scala 51:18 22:26]
  wire  _GEN_5126 = 2'h3 == state ? _GEN_4356 : valid_1_119; // @[cache.scala 51:18 22:26]
  wire  _GEN_5127 = 2'h3 == state ? _GEN_4357 : valid_1_120; // @[cache.scala 51:18 22:26]
  wire  _GEN_5128 = 2'h3 == state ? _GEN_4358 : valid_1_121; // @[cache.scala 51:18 22:26]
  wire  _GEN_5129 = 2'h3 == state ? _GEN_4359 : valid_1_122; // @[cache.scala 51:18 22:26]
  wire  _GEN_5130 = 2'h3 == state ? _GEN_4360 : valid_1_123; // @[cache.scala 51:18 22:26]
  wire  _GEN_5131 = 2'h3 == state ? _GEN_4361 : valid_1_124; // @[cache.scala 51:18 22:26]
  wire  _GEN_5132 = 2'h3 == state ? _GEN_4362 : valid_1_125; // @[cache.scala 51:18 22:26]
  wire  _GEN_5133 = 2'h3 == state ? _GEN_4363 : valid_1_126; // @[cache.scala 51:18 22:26]
  wire  _GEN_5134 = 2'h3 == state ? _GEN_4364 : valid_1_127; // @[cache.scala 51:18 22:26]
  wire [63:0] _GEN_7449 = 7'h1 == index ? ram_0_1 : ram_0_0; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7450 = 7'h2 == index ? ram_0_2 : _GEN_7449; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7451 = 7'h3 == index ? ram_0_3 : _GEN_7450; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7452 = 7'h4 == index ? ram_0_4 : _GEN_7451; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7453 = 7'h5 == index ? ram_0_5 : _GEN_7452; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7454 = 7'h6 == index ? ram_0_6 : _GEN_7453; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7455 = 7'h7 == index ? ram_0_7 : _GEN_7454; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7456 = 7'h8 == index ? ram_0_8 : _GEN_7455; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7457 = 7'h9 == index ? ram_0_9 : _GEN_7456; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7458 = 7'ha == index ? ram_0_10 : _GEN_7457; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7459 = 7'hb == index ? ram_0_11 : _GEN_7458; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7460 = 7'hc == index ? ram_0_12 : _GEN_7459; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7461 = 7'hd == index ? ram_0_13 : _GEN_7460; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7462 = 7'he == index ? ram_0_14 : _GEN_7461; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7463 = 7'hf == index ? ram_0_15 : _GEN_7462; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7464 = 7'h10 == index ? ram_0_16 : _GEN_7463; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7465 = 7'h11 == index ? ram_0_17 : _GEN_7464; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7466 = 7'h12 == index ? ram_0_18 : _GEN_7465; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7467 = 7'h13 == index ? ram_0_19 : _GEN_7466; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7468 = 7'h14 == index ? ram_0_20 : _GEN_7467; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7469 = 7'h15 == index ? ram_0_21 : _GEN_7468; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7470 = 7'h16 == index ? ram_0_22 : _GEN_7469; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7471 = 7'h17 == index ? ram_0_23 : _GEN_7470; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7472 = 7'h18 == index ? ram_0_24 : _GEN_7471; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7473 = 7'h19 == index ? ram_0_25 : _GEN_7472; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7474 = 7'h1a == index ? ram_0_26 : _GEN_7473; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7475 = 7'h1b == index ? ram_0_27 : _GEN_7474; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7476 = 7'h1c == index ? ram_0_28 : _GEN_7475; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7477 = 7'h1d == index ? ram_0_29 : _GEN_7476; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7478 = 7'h1e == index ? ram_0_30 : _GEN_7477; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7479 = 7'h1f == index ? ram_0_31 : _GEN_7478; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7480 = 7'h20 == index ? ram_0_32 : _GEN_7479; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7481 = 7'h21 == index ? ram_0_33 : _GEN_7480; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7482 = 7'h22 == index ? ram_0_34 : _GEN_7481; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7483 = 7'h23 == index ? ram_0_35 : _GEN_7482; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7484 = 7'h24 == index ? ram_0_36 : _GEN_7483; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7485 = 7'h25 == index ? ram_0_37 : _GEN_7484; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7486 = 7'h26 == index ? ram_0_38 : _GEN_7485; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7487 = 7'h27 == index ? ram_0_39 : _GEN_7486; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7488 = 7'h28 == index ? ram_0_40 : _GEN_7487; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7489 = 7'h29 == index ? ram_0_41 : _GEN_7488; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7490 = 7'h2a == index ? ram_0_42 : _GEN_7489; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7491 = 7'h2b == index ? ram_0_43 : _GEN_7490; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7492 = 7'h2c == index ? ram_0_44 : _GEN_7491; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7493 = 7'h2d == index ? ram_0_45 : _GEN_7492; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7494 = 7'h2e == index ? ram_0_46 : _GEN_7493; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7495 = 7'h2f == index ? ram_0_47 : _GEN_7494; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7496 = 7'h30 == index ? ram_0_48 : _GEN_7495; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7497 = 7'h31 == index ? ram_0_49 : _GEN_7496; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7498 = 7'h32 == index ? ram_0_50 : _GEN_7497; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7499 = 7'h33 == index ? ram_0_51 : _GEN_7498; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7500 = 7'h34 == index ? ram_0_52 : _GEN_7499; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7501 = 7'h35 == index ? ram_0_53 : _GEN_7500; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7502 = 7'h36 == index ? ram_0_54 : _GEN_7501; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7503 = 7'h37 == index ? ram_0_55 : _GEN_7502; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7504 = 7'h38 == index ? ram_0_56 : _GEN_7503; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7505 = 7'h39 == index ? ram_0_57 : _GEN_7504; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7506 = 7'h3a == index ? ram_0_58 : _GEN_7505; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7507 = 7'h3b == index ? ram_0_59 : _GEN_7506; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7508 = 7'h3c == index ? ram_0_60 : _GEN_7507; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7509 = 7'h3d == index ? ram_0_61 : _GEN_7508; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7510 = 7'h3e == index ? ram_0_62 : _GEN_7509; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7511 = 7'h3f == index ? ram_0_63 : _GEN_7510; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7512 = 7'h40 == index ? ram_0_64 : _GEN_7511; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7513 = 7'h41 == index ? ram_0_65 : _GEN_7512; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7514 = 7'h42 == index ? ram_0_66 : _GEN_7513; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7515 = 7'h43 == index ? ram_0_67 : _GEN_7514; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7516 = 7'h44 == index ? ram_0_68 : _GEN_7515; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7517 = 7'h45 == index ? ram_0_69 : _GEN_7516; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7518 = 7'h46 == index ? ram_0_70 : _GEN_7517; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7519 = 7'h47 == index ? ram_0_71 : _GEN_7518; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7520 = 7'h48 == index ? ram_0_72 : _GEN_7519; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7521 = 7'h49 == index ? ram_0_73 : _GEN_7520; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7522 = 7'h4a == index ? ram_0_74 : _GEN_7521; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7523 = 7'h4b == index ? ram_0_75 : _GEN_7522; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7524 = 7'h4c == index ? ram_0_76 : _GEN_7523; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7525 = 7'h4d == index ? ram_0_77 : _GEN_7524; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7526 = 7'h4e == index ? ram_0_78 : _GEN_7525; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7527 = 7'h4f == index ? ram_0_79 : _GEN_7526; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7528 = 7'h50 == index ? ram_0_80 : _GEN_7527; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7529 = 7'h51 == index ? ram_0_81 : _GEN_7528; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7530 = 7'h52 == index ? ram_0_82 : _GEN_7529; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7531 = 7'h53 == index ? ram_0_83 : _GEN_7530; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7532 = 7'h54 == index ? ram_0_84 : _GEN_7531; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7533 = 7'h55 == index ? ram_0_85 : _GEN_7532; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7534 = 7'h56 == index ? ram_0_86 : _GEN_7533; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7535 = 7'h57 == index ? ram_0_87 : _GEN_7534; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7536 = 7'h58 == index ? ram_0_88 : _GEN_7535; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7537 = 7'h59 == index ? ram_0_89 : _GEN_7536; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7538 = 7'h5a == index ? ram_0_90 : _GEN_7537; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7539 = 7'h5b == index ? ram_0_91 : _GEN_7538; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7540 = 7'h5c == index ? ram_0_92 : _GEN_7539; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7541 = 7'h5d == index ? ram_0_93 : _GEN_7540; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7542 = 7'h5e == index ? ram_0_94 : _GEN_7541; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7543 = 7'h5f == index ? ram_0_95 : _GEN_7542; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7544 = 7'h60 == index ? ram_0_96 : _GEN_7543; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7545 = 7'h61 == index ? ram_0_97 : _GEN_7544; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7546 = 7'h62 == index ? ram_0_98 : _GEN_7545; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7547 = 7'h63 == index ? ram_0_99 : _GEN_7546; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7548 = 7'h64 == index ? ram_0_100 : _GEN_7547; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7549 = 7'h65 == index ? ram_0_101 : _GEN_7548; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7550 = 7'h66 == index ? ram_0_102 : _GEN_7549; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7551 = 7'h67 == index ? ram_0_103 : _GEN_7550; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7552 = 7'h68 == index ? ram_0_104 : _GEN_7551; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7553 = 7'h69 == index ? ram_0_105 : _GEN_7552; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7554 = 7'h6a == index ? ram_0_106 : _GEN_7553; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7555 = 7'h6b == index ? ram_0_107 : _GEN_7554; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7556 = 7'h6c == index ? ram_0_108 : _GEN_7555; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7557 = 7'h6d == index ? ram_0_109 : _GEN_7556; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7558 = 7'h6e == index ? ram_0_110 : _GEN_7557; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7559 = 7'h6f == index ? ram_0_111 : _GEN_7558; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7560 = 7'h70 == index ? ram_0_112 : _GEN_7559; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7561 = 7'h71 == index ? ram_0_113 : _GEN_7560; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7562 = 7'h72 == index ? ram_0_114 : _GEN_7561; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7563 = 7'h73 == index ? ram_0_115 : _GEN_7562; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7564 = 7'h74 == index ? ram_0_116 : _GEN_7563; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7565 = 7'h75 == index ? ram_0_117 : _GEN_7564; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7566 = 7'h76 == index ? ram_0_118 : _GEN_7565; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7567 = 7'h77 == index ? ram_0_119 : _GEN_7566; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7568 = 7'h78 == index ? ram_0_120 : _GEN_7567; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7569 = 7'h79 == index ? ram_0_121 : _GEN_7568; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7570 = 7'h7a == index ? ram_0_122 : _GEN_7569; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7571 = 7'h7b == index ? ram_0_123 : _GEN_7570; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7572 = 7'h7c == index ? ram_0_124 : _GEN_7571; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7573 = 7'h7d == index ? ram_0_125 : _GEN_7572; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7574 = 7'h7e == index ? ram_0_126 : _GEN_7573; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7575 = 7'h7f == index ? ram_0_127 : _GEN_7574; // @[cache.scala 134:{33,33}]
  wire [63:0] _GEN_7577 = 7'h1 == index ? ram_1_1 : ram_1_0; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7578 = 7'h2 == index ? ram_1_2 : _GEN_7577; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7579 = 7'h3 == index ? ram_1_3 : _GEN_7578; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7580 = 7'h4 == index ? ram_1_4 : _GEN_7579; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7581 = 7'h5 == index ? ram_1_5 : _GEN_7580; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7582 = 7'h6 == index ? ram_1_6 : _GEN_7581; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7583 = 7'h7 == index ? ram_1_7 : _GEN_7582; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7584 = 7'h8 == index ? ram_1_8 : _GEN_7583; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7585 = 7'h9 == index ? ram_1_9 : _GEN_7584; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7586 = 7'ha == index ? ram_1_10 : _GEN_7585; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7587 = 7'hb == index ? ram_1_11 : _GEN_7586; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7588 = 7'hc == index ? ram_1_12 : _GEN_7587; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7589 = 7'hd == index ? ram_1_13 : _GEN_7588; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7590 = 7'he == index ? ram_1_14 : _GEN_7589; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7591 = 7'hf == index ? ram_1_15 : _GEN_7590; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7592 = 7'h10 == index ? ram_1_16 : _GEN_7591; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7593 = 7'h11 == index ? ram_1_17 : _GEN_7592; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7594 = 7'h12 == index ? ram_1_18 : _GEN_7593; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7595 = 7'h13 == index ? ram_1_19 : _GEN_7594; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7596 = 7'h14 == index ? ram_1_20 : _GEN_7595; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7597 = 7'h15 == index ? ram_1_21 : _GEN_7596; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7598 = 7'h16 == index ? ram_1_22 : _GEN_7597; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7599 = 7'h17 == index ? ram_1_23 : _GEN_7598; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7600 = 7'h18 == index ? ram_1_24 : _GEN_7599; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7601 = 7'h19 == index ? ram_1_25 : _GEN_7600; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7602 = 7'h1a == index ? ram_1_26 : _GEN_7601; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7603 = 7'h1b == index ? ram_1_27 : _GEN_7602; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7604 = 7'h1c == index ? ram_1_28 : _GEN_7603; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7605 = 7'h1d == index ? ram_1_29 : _GEN_7604; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7606 = 7'h1e == index ? ram_1_30 : _GEN_7605; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7607 = 7'h1f == index ? ram_1_31 : _GEN_7606; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7608 = 7'h20 == index ? ram_1_32 : _GEN_7607; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7609 = 7'h21 == index ? ram_1_33 : _GEN_7608; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7610 = 7'h22 == index ? ram_1_34 : _GEN_7609; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7611 = 7'h23 == index ? ram_1_35 : _GEN_7610; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7612 = 7'h24 == index ? ram_1_36 : _GEN_7611; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7613 = 7'h25 == index ? ram_1_37 : _GEN_7612; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7614 = 7'h26 == index ? ram_1_38 : _GEN_7613; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7615 = 7'h27 == index ? ram_1_39 : _GEN_7614; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7616 = 7'h28 == index ? ram_1_40 : _GEN_7615; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7617 = 7'h29 == index ? ram_1_41 : _GEN_7616; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7618 = 7'h2a == index ? ram_1_42 : _GEN_7617; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7619 = 7'h2b == index ? ram_1_43 : _GEN_7618; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7620 = 7'h2c == index ? ram_1_44 : _GEN_7619; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7621 = 7'h2d == index ? ram_1_45 : _GEN_7620; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7622 = 7'h2e == index ? ram_1_46 : _GEN_7621; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7623 = 7'h2f == index ? ram_1_47 : _GEN_7622; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7624 = 7'h30 == index ? ram_1_48 : _GEN_7623; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7625 = 7'h31 == index ? ram_1_49 : _GEN_7624; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7626 = 7'h32 == index ? ram_1_50 : _GEN_7625; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7627 = 7'h33 == index ? ram_1_51 : _GEN_7626; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7628 = 7'h34 == index ? ram_1_52 : _GEN_7627; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7629 = 7'h35 == index ? ram_1_53 : _GEN_7628; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7630 = 7'h36 == index ? ram_1_54 : _GEN_7629; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7631 = 7'h37 == index ? ram_1_55 : _GEN_7630; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7632 = 7'h38 == index ? ram_1_56 : _GEN_7631; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7633 = 7'h39 == index ? ram_1_57 : _GEN_7632; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7634 = 7'h3a == index ? ram_1_58 : _GEN_7633; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7635 = 7'h3b == index ? ram_1_59 : _GEN_7634; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7636 = 7'h3c == index ? ram_1_60 : _GEN_7635; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7637 = 7'h3d == index ? ram_1_61 : _GEN_7636; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7638 = 7'h3e == index ? ram_1_62 : _GEN_7637; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7639 = 7'h3f == index ? ram_1_63 : _GEN_7638; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7640 = 7'h40 == index ? ram_1_64 : _GEN_7639; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7641 = 7'h41 == index ? ram_1_65 : _GEN_7640; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7642 = 7'h42 == index ? ram_1_66 : _GEN_7641; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7643 = 7'h43 == index ? ram_1_67 : _GEN_7642; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7644 = 7'h44 == index ? ram_1_68 : _GEN_7643; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7645 = 7'h45 == index ? ram_1_69 : _GEN_7644; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7646 = 7'h46 == index ? ram_1_70 : _GEN_7645; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7647 = 7'h47 == index ? ram_1_71 : _GEN_7646; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7648 = 7'h48 == index ? ram_1_72 : _GEN_7647; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7649 = 7'h49 == index ? ram_1_73 : _GEN_7648; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7650 = 7'h4a == index ? ram_1_74 : _GEN_7649; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7651 = 7'h4b == index ? ram_1_75 : _GEN_7650; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7652 = 7'h4c == index ? ram_1_76 : _GEN_7651; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7653 = 7'h4d == index ? ram_1_77 : _GEN_7652; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7654 = 7'h4e == index ? ram_1_78 : _GEN_7653; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7655 = 7'h4f == index ? ram_1_79 : _GEN_7654; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7656 = 7'h50 == index ? ram_1_80 : _GEN_7655; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7657 = 7'h51 == index ? ram_1_81 : _GEN_7656; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7658 = 7'h52 == index ? ram_1_82 : _GEN_7657; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7659 = 7'h53 == index ? ram_1_83 : _GEN_7658; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7660 = 7'h54 == index ? ram_1_84 : _GEN_7659; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7661 = 7'h55 == index ? ram_1_85 : _GEN_7660; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7662 = 7'h56 == index ? ram_1_86 : _GEN_7661; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7663 = 7'h57 == index ? ram_1_87 : _GEN_7662; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7664 = 7'h58 == index ? ram_1_88 : _GEN_7663; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7665 = 7'h59 == index ? ram_1_89 : _GEN_7664; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7666 = 7'h5a == index ? ram_1_90 : _GEN_7665; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7667 = 7'h5b == index ? ram_1_91 : _GEN_7666; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7668 = 7'h5c == index ? ram_1_92 : _GEN_7667; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7669 = 7'h5d == index ? ram_1_93 : _GEN_7668; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7670 = 7'h5e == index ? ram_1_94 : _GEN_7669; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7671 = 7'h5f == index ? ram_1_95 : _GEN_7670; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7672 = 7'h60 == index ? ram_1_96 : _GEN_7671; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7673 = 7'h61 == index ? ram_1_97 : _GEN_7672; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7674 = 7'h62 == index ? ram_1_98 : _GEN_7673; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7675 = 7'h63 == index ? ram_1_99 : _GEN_7674; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7676 = 7'h64 == index ? ram_1_100 : _GEN_7675; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7677 = 7'h65 == index ? ram_1_101 : _GEN_7676; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7678 = 7'h66 == index ? ram_1_102 : _GEN_7677; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7679 = 7'h67 == index ? ram_1_103 : _GEN_7678; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7680 = 7'h68 == index ? ram_1_104 : _GEN_7679; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7681 = 7'h69 == index ? ram_1_105 : _GEN_7680; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7682 = 7'h6a == index ? ram_1_106 : _GEN_7681; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7683 = 7'h6b == index ? ram_1_107 : _GEN_7682; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7684 = 7'h6c == index ? ram_1_108 : _GEN_7683; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7685 = 7'h6d == index ? ram_1_109 : _GEN_7684; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7686 = 7'h6e == index ? ram_1_110 : _GEN_7685; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7687 = 7'h6f == index ? ram_1_111 : _GEN_7686; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7688 = 7'h70 == index ? ram_1_112 : _GEN_7687; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7689 = 7'h71 == index ? ram_1_113 : _GEN_7688; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7690 = 7'h72 == index ? ram_1_114 : _GEN_7689; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7691 = 7'h73 == index ? ram_1_115 : _GEN_7690; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7692 = 7'h74 == index ? ram_1_116 : _GEN_7691; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7693 = 7'h75 == index ? ram_1_117 : _GEN_7692; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7694 = 7'h76 == index ? ram_1_118 : _GEN_7693; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7695 = 7'h77 == index ? ram_1_119 : _GEN_7694; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7696 = 7'h78 == index ? ram_1_120 : _GEN_7695; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7697 = 7'h79 == index ? ram_1_121 : _GEN_7696; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7698 = 7'h7a == index ? ram_1_122 : _GEN_7697; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7699 = 7'h7b == index ? ram_1_123 : _GEN_7698; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7700 = 7'h7c == index ? ram_1_124 : _GEN_7699; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7701 = 7'h7d == index ? ram_1_125 : _GEN_7700; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7702 = 7'h7e == index ? ram_1_126 : _GEN_7701; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7703 = 7'h7f == index ? ram_1_127 : _GEN_7702; // @[cache.scala 142:{33,33}]
  wire [63:0] _GEN_7704 = way1_hit ? _GEN_7703 : 64'h0; // @[cache.scala 141:33 142:33 149:33]
  wire [63:0] _GEN_7708 = way0_hit ? _GEN_7575 : _GEN_7704; // @[cache.scala 133:23 134:33]
  wire  _GEN_7710 = way0_hit | way1_hit; // @[cache.scala 133:23 136:34]
  wire  _T_21 = state == 2'h2; // @[cache.scala 156:21]
  wire  _GEN_7721 = state == 2'h1 ? 1'h0 : _T_21; // @[cache.scala 123:31 124:27]
  wire  _GEN_7723 = state == 2'h1 ? 1'h0 : io_from_ifu_rready; // @[cache.scala 123:31 126:26]
  wire [63:0] _GEN_7725 = state == 2'h1 ? _GEN_7708 : 64'h0; // @[cache.scala 123:31]
  wire  _GEN_7727 = state == 2'h1 & _GEN_7710; // @[cache.scala 123:31]
  assign io_to_ifu_rdata = state == 2'h0 ? 64'h0 : _GEN_7725; // @[cache.scala 107:23 108:25]
  assign io_to_ifu_rvalid = state == 2'h0 ? 1'h0 : _GEN_7727; // @[cache.scala 107:23 110:26]
  assign io_to_axi_araddr = io_from_ifu_araddr; // @[cache.scala 107:23 115:26]
  assign io_to_axi_arvalid = state == 2'h0 ? 1'h0 : _GEN_7721; // @[cache.scala 107:23 114:27]
  assign io_to_axi_rready = state == 2'h0 ? io_from_ifu_rready : _GEN_7723; // @[cache.scala 107:23 116:26]
  always @(posedge clock) begin
    if (reset) begin // @[cache.scala 17:24]
      ram_0_0 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_0 <= _GEN_4366;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_1 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_1 <= _GEN_4367;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_2 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_2 <= _GEN_4368;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_3 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_3 <= _GEN_4369;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_4 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_4 <= _GEN_4370;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_5 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_5 <= _GEN_4371;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_6 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_6 <= _GEN_4372;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_7 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_7 <= _GEN_4373;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_8 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_8 <= _GEN_4374;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_9 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_9 <= _GEN_4375;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_10 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_10 <= _GEN_4376;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_11 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_11 <= _GEN_4377;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_12 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_12 <= _GEN_4378;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_13 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_13 <= _GEN_4379;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_14 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_14 <= _GEN_4380;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_15 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_15 <= _GEN_4381;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_16 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_16 <= _GEN_4382;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_17 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_17 <= _GEN_4383;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_18 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_18 <= _GEN_4384;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_19 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_19 <= _GEN_4385;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_20 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_20 <= _GEN_4386;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_21 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_21 <= _GEN_4387;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_22 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_22 <= _GEN_4388;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_23 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_23 <= _GEN_4389;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_24 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_24 <= _GEN_4390;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_25 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_25 <= _GEN_4391;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_26 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_26 <= _GEN_4392;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_27 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_27 <= _GEN_4393;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_28 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_28 <= _GEN_4394;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_29 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_29 <= _GEN_4395;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_30 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_30 <= _GEN_4396;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_31 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_31 <= _GEN_4397;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_32 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_32 <= _GEN_4398;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_33 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_33 <= _GEN_4399;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_34 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_34 <= _GEN_4400;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_35 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_35 <= _GEN_4401;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_36 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_36 <= _GEN_4402;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_37 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_37 <= _GEN_4403;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_38 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_38 <= _GEN_4404;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_39 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_39 <= _GEN_4405;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_40 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_40 <= _GEN_4406;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_41 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_41 <= _GEN_4407;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_42 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_42 <= _GEN_4408;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_43 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_43 <= _GEN_4409;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_44 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_44 <= _GEN_4410;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_45 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_45 <= _GEN_4411;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_46 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_46 <= _GEN_4412;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_47 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_47 <= _GEN_4413;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_48 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_48 <= _GEN_4414;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_49 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_49 <= _GEN_4415;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_50 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_50 <= _GEN_4416;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_51 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_51 <= _GEN_4417;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_52 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_52 <= _GEN_4418;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_53 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_53 <= _GEN_4419;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_54 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_54 <= _GEN_4420;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_55 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_55 <= _GEN_4421;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_56 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_56 <= _GEN_4422;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_57 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_57 <= _GEN_4423;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_58 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_58 <= _GEN_4424;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_59 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_59 <= _GEN_4425;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_60 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_60 <= _GEN_4426;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_61 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_61 <= _GEN_4427;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_62 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_62 <= _GEN_4428;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_63 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_63 <= _GEN_4429;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_64 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_64 <= _GEN_4430;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_65 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_65 <= _GEN_4431;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_66 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_66 <= _GEN_4432;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_67 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_67 <= _GEN_4433;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_68 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_68 <= _GEN_4434;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_69 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_69 <= _GEN_4435;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_70 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_70 <= _GEN_4436;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_71 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_71 <= _GEN_4437;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_72 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_72 <= _GEN_4438;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_73 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_73 <= _GEN_4439;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_74 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_74 <= _GEN_4440;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_75 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_75 <= _GEN_4441;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_76 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_76 <= _GEN_4442;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_77 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_77 <= _GEN_4443;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_78 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_78 <= _GEN_4444;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_79 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_79 <= _GEN_4445;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_80 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_80 <= _GEN_4446;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_81 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_81 <= _GEN_4447;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_82 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_82 <= _GEN_4448;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_83 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_83 <= _GEN_4449;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_84 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_84 <= _GEN_4450;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_85 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_85 <= _GEN_4451;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_86 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_86 <= _GEN_4452;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_87 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_87 <= _GEN_4453;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_88 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_88 <= _GEN_4454;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_89 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_89 <= _GEN_4455;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_90 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_90 <= _GEN_4456;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_91 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_91 <= _GEN_4457;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_92 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_92 <= _GEN_4458;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_93 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_93 <= _GEN_4459;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_94 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_94 <= _GEN_4460;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_95 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_95 <= _GEN_4461;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_96 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_96 <= _GEN_4462;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_97 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_97 <= _GEN_4463;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_98 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_98 <= _GEN_4464;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_99 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_99 <= _GEN_4465;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_100 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_100 <= _GEN_4466;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_101 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_101 <= _GEN_4467;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_102 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_102 <= _GEN_4468;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_103 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_103 <= _GEN_4469;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_104 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_104 <= _GEN_4470;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_105 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_105 <= _GEN_4471;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_106 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_106 <= _GEN_4472;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_107 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_107 <= _GEN_4473;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_108 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_108 <= _GEN_4474;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_109 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_109 <= _GEN_4475;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_110 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_110 <= _GEN_4476;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_111 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_111 <= _GEN_4477;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_112 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_112 <= _GEN_4478;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_113 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_113 <= _GEN_4479;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_114 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_114 <= _GEN_4480;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_115 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_115 <= _GEN_4481;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_116 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_116 <= _GEN_4482;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_117 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_117 <= _GEN_4483;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_118 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_118 <= _GEN_4484;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_119 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_119 <= _GEN_4485;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_120 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_120 <= _GEN_4486;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_121 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_121 <= _GEN_4487;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_122 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_122 <= _GEN_4488;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_123 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_123 <= _GEN_4489;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_124 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_124 <= _GEN_4490;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_125 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_125 <= _GEN_4491;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_126 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_126 <= _GEN_4492;
        end
      end
    end
    if (reset) begin // @[cache.scala 17:24]
      ram_0_127 <= 64'h0; // @[cache.scala 17:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_0_127 <= _GEN_4493;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_0 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_0 <= _GEN_4751;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_1 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_1 <= _GEN_4752;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_2 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_2 <= _GEN_4753;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_3 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_3 <= _GEN_4754;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_4 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_4 <= _GEN_4755;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_5 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_5 <= _GEN_4756;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_6 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_6 <= _GEN_4757;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_7 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_7 <= _GEN_4758;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_8 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_8 <= _GEN_4759;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_9 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_9 <= _GEN_4760;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_10 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_10 <= _GEN_4761;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_11 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_11 <= _GEN_4762;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_12 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_12 <= _GEN_4763;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_13 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_13 <= _GEN_4764;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_14 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_14 <= _GEN_4765;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_15 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_15 <= _GEN_4766;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_16 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_16 <= _GEN_4767;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_17 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_17 <= _GEN_4768;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_18 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_18 <= _GEN_4769;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_19 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_19 <= _GEN_4770;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_20 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_20 <= _GEN_4771;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_21 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_21 <= _GEN_4772;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_22 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_22 <= _GEN_4773;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_23 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_23 <= _GEN_4774;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_24 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_24 <= _GEN_4775;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_25 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_25 <= _GEN_4776;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_26 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_26 <= _GEN_4777;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_27 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_27 <= _GEN_4778;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_28 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_28 <= _GEN_4779;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_29 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_29 <= _GEN_4780;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_30 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_30 <= _GEN_4781;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_31 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_31 <= _GEN_4782;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_32 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_32 <= _GEN_4783;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_33 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_33 <= _GEN_4784;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_34 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_34 <= _GEN_4785;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_35 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_35 <= _GEN_4786;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_36 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_36 <= _GEN_4787;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_37 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_37 <= _GEN_4788;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_38 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_38 <= _GEN_4789;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_39 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_39 <= _GEN_4790;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_40 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_40 <= _GEN_4791;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_41 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_41 <= _GEN_4792;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_42 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_42 <= _GEN_4793;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_43 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_43 <= _GEN_4794;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_44 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_44 <= _GEN_4795;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_45 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_45 <= _GEN_4796;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_46 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_46 <= _GEN_4797;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_47 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_47 <= _GEN_4798;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_48 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_48 <= _GEN_4799;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_49 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_49 <= _GEN_4800;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_50 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_50 <= _GEN_4801;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_51 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_51 <= _GEN_4802;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_52 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_52 <= _GEN_4803;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_53 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_53 <= _GEN_4804;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_54 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_54 <= _GEN_4805;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_55 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_55 <= _GEN_4806;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_56 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_56 <= _GEN_4807;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_57 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_57 <= _GEN_4808;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_58 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_58 <= _GEN_4809;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_59 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_59 <= _GEN_4810;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_60 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_60 <= _GEN_4811;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_61 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_61 <= _GEN_4812;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_62 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_62 <= _GEN_4813;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_63 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_63 <= _GEN_4814;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_64 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_64 <= _GEN_4815;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_65 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_65 <= _GEN_4816;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_66 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_66 <= _GEN_4817;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_67 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_67 <= _GEN_4818;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_68 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_68 <= _GEN_4819;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_69 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_69 <= _GEN_4820;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_70 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_70 <= _GEN_4821;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_71 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_71 <= _GEN_4822;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_72 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_72 <= _GEN_4823;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_73 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_73 <= _GEN_4824;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_74 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_74 <= _GEN_4825;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_75 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_75 <= _GEN_4826;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_76 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_76 <= _GEN_4827;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_77 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_77 <= _GEN_4828;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_78 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_78 <= _GEN_4829;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_79 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_79 <= _GEN_4830;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_80 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_80 <= _GEN_4831;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_81 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_81 <= _GEN_4832;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_82 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_82 <= _GEN_4833;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_83 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_83 <= _GEN_4834;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_84 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_84 <= _GEN_4835;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_85 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_85 <= _GEN_4836;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_86 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_86 <= _GEN_4837;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_87 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_87 <= _GEN_4838;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_88 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_88 <= _GEN_4839;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_89 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_89 <= _GEN_4840;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_90 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_90 <= _GEN_4841;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_91 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_91 <= _GEN_4842;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_92 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_92 <= _GEN_4843;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_93 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_93 <= _GEN_4844;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_94 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_94 <= _GEN_4845;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_95 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_95 <= _GEN_4846;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_96 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_96 <= _GEN_4847;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_97 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_97 <= _GEN_4848;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_98 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_98 <= _GEN_4849;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_99 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_99 <= _GEN_4850;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_100 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_100 <= _GEN_4851;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_101 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_101 <= _GEN_4852;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_102 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_102 <= _GEN_4853;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_103 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_103 <= _GEN_4854;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_104 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_104 <= _GEN_4855;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_105 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_105 <= _GEN_4856;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_106 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_106 <= _GEN_4857;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_107 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_107 <= _GEN_4858;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_108 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_108 <= _GEN_4859;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_109 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_109 <= _GEN_4860;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_110 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_110 <= _GEN_4861;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_111 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_111 <= _GEN_4862;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_112 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_112 <= _GEN_4863;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_113 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_113 <= _GEN_4864;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_114 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_114 <= _GEN_4865;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_115 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_115 <= _GEN_4866;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_116 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_116 <= _GEN_4867;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_117 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_117 <= _GEN_4868;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_118 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_118 <= _GEN_4869;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_119 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_119 <= _GEN_4870;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_120 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_120 <= _GEN_4871;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_121 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_121 <= _GEN_4872;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_122 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_122 <= _GEN_4873;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_123 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_123 <= _GEN_4874;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_124 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_124 <= _GEN_4875;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_125 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_125 <= _GEN_4876;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_126 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_126 <= _GEN_4877;
        end
      end
    end
    if (reset) begin // @[cache.scala 18:24]
      ram_1_127 <= 64'h0; // @[cache.scala 18:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          ram_1_127 <= _GEN_4878;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_0 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_0 <= _GEN_4494;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_1 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_1 <= _GEN_4495;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_2 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_2 <= _GEN_4496;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_3 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_3 <= _GEN_4497;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_4 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_4 <= _GEN_4498;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_5 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_5 <= _GEN_4499;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_6 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_6 <= _GEN_4500;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_7 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_7 <= _GEN_4501;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_8 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_8 <= _GEN_4502;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_9 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_9 <= _GEN_4503;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_10 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_10 <= _GEN_4504;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_11 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_11 <= _GEN_4505;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_12 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_12 <= _GEN_4506;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_13 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_13 <= _GEN_4507;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_14 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_14 <= _GEN_4508;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_15 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_15 <= _GEN_4509;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_16 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_16 <= _GEN_4510;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_17 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_17 <= _GEN_4511;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_18 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_18 <= _GEN_4512;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_19 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_19 <= _GEN_4513;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_20 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_20 <= _GEN_4514;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_21 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_21 <= _GEN_4515;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_22 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_22 <= _GEN_4516;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_23 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_23 <= _GEN_4517;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_24 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_24 <= _GEN_4518;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_25 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_25 <= _GEN_4519;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_26 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_26 <= _GEN_4520;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_27 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_27 <= _GEN_4521;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_28 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_28 <= _GEN_4522;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_29 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_29 <= _GEN_4523;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_30 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_30 <= _GEN_4524;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_31 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_31 <= _GEN_4525;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_32 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_32 <= _GEN_4526;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_33 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_33 <= _GEN_4527;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_34 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_34 <= _GEN_4528;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_35 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_35 <= _GEN_4529;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_36 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_36 <= _GEN_4530;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_37 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_37 <= _GEN_4531;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_38 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_38 <= _GEN_4532;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_39 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_39 <= _GEN_4533;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_40 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_40 <= _GEN_4534;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_41 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_41 <= _GEN_4535;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_42 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_42 <= _GEN_4536;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_43 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_43 <= _GEN_4537;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_44 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_44 <= _GEN_4538;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_45 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_45 <= _GEN_4539;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_46 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_46 <= _GEN_4540;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_47 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_47 <= _GEN_4541;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_48 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_48 <= _GEN_4542;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_49 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_49 <= _GEN_4543;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_50 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_50 <= _GEN_4544;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_51 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_51 <= _GEN_4545;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_52 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_52 <= _GEN_4546;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_53 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_53 <= _GEN_4547;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_54 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_54 <= _GEN_4548;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_55 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_55 <= _GEN_4549;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_56 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_56 <= _GEN_4550;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_57 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_57 <= _GEN_4551;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_58 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_58 <= _GEN_4552;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_59 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_59 <= _GEN_4553;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_60 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_60 <= _GEN_4554;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_61 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_61 <= _GEN_4555;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_62 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_62 <= _GEN_4556;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_63 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_63 <= _GEN_4557;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_64 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_64 <= _GEN_4558;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_65 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_65 <= _GEN_4559;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_66 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_66 <= _GEN_4560;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_67 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_67 <= _GEN_4561;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_68 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_68 <= _GEN_4562;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_69 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_69 <= _GEN_4563;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_70 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_70 <= _GEN_4564;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_71 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_71 <= _GEN_4565;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_72 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_72 <= _GEN_4566;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_73 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_73 <= _GEN_4567;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_74 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_74 <= _GEN_4568;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_75 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_75 <= _GEN_4569;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_76 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_76 <= _GEN_4570;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_77 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_77 <= _GEN_4571;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_78 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_78 <= _GEN_4572;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_79 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_79 <= _GEN_4573;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_80 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_80 <= _GEN_4574;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_81 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_81 <= _GEN_4575;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_82 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_82 <= _GEN_4576;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_83 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_83 <= _GEN_4577;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_84 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_84 <= _GEN_4578;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_85 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_85 <= _GEN_4579;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_86 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_86 <= _GEN_4580;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_87 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_87 <= _GEN_4581;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_88 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_88 <= _GEN_4582;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_89 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_89 <= _GEN_4583;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_90 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_90 <= _GEN_4584;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_91 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_91 <= _GEN_4585;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_92 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_92 <= _GEN_4586;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_93 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_93 <= _GEN_4587;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_94 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_94 <= _GEN_4588;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_95 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_95 <= _GEN_4589;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_96 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_96 <= _GEN_4590;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_97 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_97 <= _GEN_4591;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_98 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_98 <= _GEN_4592;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_99 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_99 <= _GEN_4593;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_100 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_100 <= _GEN_4594;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_101 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_101 <= _GEN_4595;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_102 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_102 <= _GEN_4596;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_103 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_103 <= _GEN_4597;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_104 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_104 <= _GEN_4598;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_105 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_105 <= _GEN_4599;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_106 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_106 <= _GEN_4600;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_107 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_107 <= _GEN_4601;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_108 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_108 <= _GEN_4602;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_109 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_109 <= _GEN_4603;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_110 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_110 <= _GEN_4604;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_111 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_111 <= _GEN_4605;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_112 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_112 <= _GEN_4606;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_113 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_113 <= _GEN_4607;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_114 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_114 <= _GEN_4608;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_115 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_115 <= _GEN_4609;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_116 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_116 <= _GEN_4610;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_117 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_117 <= _GEN_4611;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_118 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_118 <= _GEN_4612;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_119 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_119 <= _GEN_4613;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_120 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_120 <= _GEN_4614;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_121 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_121 <= _GEN_4615;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_122 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_122 <= _GEN_4616;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_123 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_123 <= _GEN_4617;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_124 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_124 <= _GEN_4618;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_125 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_125 <= _GEN_4619;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_126 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_126 <= _GEN_4620;
        end
      end
    end
    if (reset) begin // @[cache.scala 19:24]
      tag_0_127 <= 32'h0; // @[cache.scala 19:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_0_127 <= _GEN_4621;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_0 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_0 <= _GEN_4879;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_1 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_1 <= _GEN_4880;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_2 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_2 <= _GEN_4881;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_3 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_3 <= _GEN_4882;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_4 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_4 <= _GEN_4883;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_5 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_5 <= _GEN_4884;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_6 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_6 <= _GEN_4885;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_7 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_7 <= _GEN_4886;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_8 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_8 <= _GEN_4887;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_9 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_9 <= _GEN_4888;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_10 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_10 <= _GEN_4889;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_11 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_11 <= _GEN_4890;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_12 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_12 <= _GEN_4891;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_13 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_13 <= _GEN_4892;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_14 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_14 <= _GEN_4893;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_15 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_15 <= _GEN_4894;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_16 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_16 <= _GEN_4895;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_17 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_17 <= _GEN_4896;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_18 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_18 <= _GEN_4897;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_19 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_19 <= _GEN_4898;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_20 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_20 <= _GEN_4899;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_21 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_21 <= _GEN_4900;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_22 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_22 <= _GEN_4901;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_23 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_23 <= _GEN_4902;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_24 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_24 <= _GEN_4903;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_25 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_25 <= _GEN_4904;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_26 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_26 <= _GEN_4905;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_27 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_27 <= _GEN_4906;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_28 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_28 <= _GEN_4907;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_29 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_29 <= _GEN_4908;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_30 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_30 <= _GEN_4909;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_31 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_31 <= _GEN_4910;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_32 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_32 <= _GEN_4911;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_33 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_33 <= _GEN_4912;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_34 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_34 <= _GEN_4913;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_35 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_35 <= _GEN_4914;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_36 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_36 <= _GEN_4915;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_37 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_37 <= _GEN_4916;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_38 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_38 <= _GEN_4917;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_39 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_39 <= _GEN_4918;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_40 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_40 <= _GEN_4919;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_41 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_41 <= _GEN_4920;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_42 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_42 <= _GEN_4921;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_43 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_43 <= _GEN_4922;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_44 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_44 <= _GEN_4923;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_45 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_45 <= _GEN_4924;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_46 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_46 <= _GEN_4925;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_47 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_47 <= _GEN_4926;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_48 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_48 <= _GEN_4927;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_49 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_49 <= _GEN_4928;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_50 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_50 <= _GEN_4929;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_51 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_51 <= _GEN_4930;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_52 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_52 <= _GEN_4931;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_53 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_53 <= _GEN_4932;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_54 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_54 <= _GEN_4933;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_55 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_55 <= _GEN_4934;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_56 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_56 <= _GEN_4935;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_57 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_57 <= _GEN_4936;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_58 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_58 <= _GEN_4937;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_59 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_59 <= _GEN_4938;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_60 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_60 <= _GEN_4939;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_61 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_61 <= _GEN_4940;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_62 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_62 <= _GEN_4941;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_63 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_63 <= _GEN_4942;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_64 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_64 <= _GEN_4943;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_65 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_65 <= _GEN_4944;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_66 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_66 <= _GEN_4945;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_67 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_67 <= _GEN_4946;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_68 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_68 <= _GEN_4947;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_69 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_69 <= _GEN_4948;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_70 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_70 <= _GEN_4949;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_71 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_71 <= _GEN_4950;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_72 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_72 <= _GEN_4951;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_73 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_73 <= _GEN_4952;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_74 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_74 <= _GEN_4953;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_75 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_75 <= _GEN_4954;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_76 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_76 <= _GEN_4955;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_77 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_77 <= _GEN_4956;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_78 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_78 <= _GEN_4957;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_79 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_79 <= _GEN_4958;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_80 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_80 <= _GEN_4959;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_81 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_81 <= _GEN_4960;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_82 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_82 <= _GEN_4961;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_83 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_83 <= _GEN_4962;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_84 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_84 <= _GEN_4963;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_85 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_85 <= _GEN_4964;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_86 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_86 <= _GEN_4965;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_87 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_87 <= _GEN_4966;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_88 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_88 <= _GEN_4967;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_89 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_89 <= _GEN_4968;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_90 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_90 <= _GEN_4969;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_91 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_91 <= _GEN_4970;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_92 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_92 <= _GEN_4971;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_93 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_93 <= _GEN_4972;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_94 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_94 <= _GEN_4973;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_95 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_95 <= _GEN_4974;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_96 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_96 <= _GEN_4975;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_97 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_97 <= _GEN_4976;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_98 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_98 <= _GEN_4977;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_99 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_99 <= _GEN_4978;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_100 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_100 <= _GEN_4979;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_101 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_101 <= _GEN_4980;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_102 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_102 <= _GEN_4981;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_103 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_103 <= _GEN_4982;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_104 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_104 <= _GEN_4983;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_105 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_105 <= _GEN_4984;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_106 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_106 <= _GEN_4985;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_107 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_107 <= _GEN_4986;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_108 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_108 <= _GEN_4987;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_109 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_109 <= _GEN_4988;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_110 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_110 <= _GEN_4989;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_111 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_111 <= _GEN_4990;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_112 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_112 <= _GEN_4991;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_113 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_113 <= _GEN_4992;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_114 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_114 <= _GEN_4993;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_115 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_115 <= _GEN_4994;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_116 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_116 <= _GEN_4995;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_117 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_117 <= _GEN_4996;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_118 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_118 <= _GEN_4997;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_119 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_119 <= _GEN_4998;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_120 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_120 <= _GEN_4999;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_121 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_121 <= _GEN_5000;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_122 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_122 <= _GEN_5001;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_123 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_123 <= _GEN_5002;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_124 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_124 <= _GEN_5003;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_125 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_125 <= _GEN_5004;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_126 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_126 <= _GEN_5005;
        end
      end
    end
    if (reset) begin // @[cache.scala 20:24]
      tag_1_127 <= 32'h0; // @[cache.scala 20:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          tag_1_127 <= _GEN_5006;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_0 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_0 <= _GEN_4622;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_1 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_1 <= _GEN_4623;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_2 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_2 <= _GEN_4624;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_3 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_3 <= _GEN_4625;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_4 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_4 <= _GEN_4626;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_5 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_5 <= _GEN_4627;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_6 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_6 <= _GEN_4628;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_7 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_7 <= _GEN_4629;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_8 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_8 <= _GEN_4630;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_9 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_9 <= _GEN_4631;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_10 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_10 <= _GEN_4632;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_11 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_11 <= _GEN_4633;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_12 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_12 <= _GEN_4634;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_13 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_13 <= _GEN_4635;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_14 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_14 <= _GEN_4636;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_15 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_15 <= _GEN_4637;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_16 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_16 <= _GEN_4638;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_17 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_17 <= _GEN_4639;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_18 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_18 <= _GEN_4640;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_19 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_19 <= _GEN_4641;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_20 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_20 <= _GEN_4642;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_21 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_21 <= _GEN_4643;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_22 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_22 <= _GEN_4644;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_23 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_23 <= _GEN_4645;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_24 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_24 <= _GEN_4646;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_25 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_25 <= _GEN_4647;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_26 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_26 <= _GEN_4648;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_27 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_27 <= _GEN_4649;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_28 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_28 <= _GEN_4650;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_29 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_29 <= _GEN_4651;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_30 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_30 <= _GEN_4652;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_31 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_31 <= _GEN_4653;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_32 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_32 <= _GEN_4654;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_33 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_33 <= _GEN_4655;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_34 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_34 <= _GEN_4656;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_35 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_35 <= _GEN_4657;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_36 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_36 <= _GEN_4658;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_37 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_37 <= _GEN_4659;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_38 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_38 <= _GEN_4660;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_39 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_39 <= _GEN_4661;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_40 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_40 <= _GEN_4662;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_41 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_41 <= _GEN_4663;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_42 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_42 <= _GEN_4664;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_43 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_43 <= _GEN_4665;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_44 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_44 <= _GEN_4666;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_45 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_45 <= _GEN_4667;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_46 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_46 <= _GEN_4668;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_47 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_47 <= _GEN_4669;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_48 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_48 <= _GEN_4670;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_49 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_49 <= _GEN_4671;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_50 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_50 <= _GEN_4672;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_51 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_51 <= _GEN_4673;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_52 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_52 <= _GEN_4674;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_53 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_53 <= _GEN_4675;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_54 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_54 <= _GEN_4676;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_55 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_55 <= _GEN_4677;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_56 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_56 <= _GEN_4678;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_57 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_57 <= _GEN_4679;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_58 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_58 <= _GEN_4680;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_59 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_59 <= _GEN_4681;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_60 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_60 <= _GEN_4682;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_61 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_61 <= _GEN_4683;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_62 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_62 <= _GEN_4684;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_63 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_63 <= _GEN_4685;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_64 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_64 <= _GEN_4686;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_65 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_65 <= _GEN_4687;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_66 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_66 <= _GEN_4688;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_67 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_67 <= _GEN_4689;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_68 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_68 <= _GEN_4690;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_69 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_69 <= _GEN_4691;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_70 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_70 <= _GEN_4692;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_71 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_71 <= _GEN_4693;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_72 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_72 <= _GEN_4694;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_73 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_73 <= _GEN_4695;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_74 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_74 <= _GEN_4696;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_75 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_75 <= _GEN_4697;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_76 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_76 <= _GEN_4698;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_77 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_77 <= _GEN_4699;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_78 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_78 <= _GEN_4700;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_79 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_79 <= _GEN_4701;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_80 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_80 <= _GEN_4702;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_81 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_81 <= _GEN_4703;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_82 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_82 <= _GEN_4704;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_83 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_83 <= _GEN_4705;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_84 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_84 <= _GEN_4706;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_85 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_85 <= _GEN_4707;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_86 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_86 <= _GEN_4708;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_87 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_87 <= _GEN_4709;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_88 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_88 <= _GEN_4710;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_89 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_89 <= _GEN_4711;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_90 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_90 <= _GEN_4712;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_91 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_91 <= _GEN_4713;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_92 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_92 <= _GEN_4714;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_93 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_93 <= _GEN_4715;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_94 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_94 <= _GEN_4716;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_95 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_95 <= _GEN_4717;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_96 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_96 <= _GEN_4718;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_97 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_97 <= _GEN_4719;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_98 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_98 <= _GEN_4720;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_99 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_99 <= _GEN_4721;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_100 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_100 <= _GEN_4722;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_101 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_101 <= _GEN_4723;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_102 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_102 <= _GEN_4724;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_103 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_103 <= _GEN_4725;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_104 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_104 <= _GEN_4726;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_105 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_105 <= _GEN_4727;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_106 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_106 <= _GEN_4728;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_107 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_107 <= _GEN_4729;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_108 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_108 <= _GEN_4730;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_109 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_109 <= _GEN_4731;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_110 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_110 <= _GEN_4732;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_111 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_111 <= _GEN_4733;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_112 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_112 <= _GEN_4734;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_113 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_113 <= _GEN_4735;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_114 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_114 <= _GEN_4736;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_115 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_115 <= _GEN_4737;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_116 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_116 <= _GEN_4738;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_117 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_117 <= _GEN_4739;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_118 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_118 <= _GEN_4740;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_119 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_119 <= _GEN_4741;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_120 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_120 <= _GEN_4742;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_121 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_121 <= _GEN_4743;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_122 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_122 <= _GEN_4744;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_123 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_123 <= _GEN_4745;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_124 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_124 <= _GEN_4746;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_125 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_125 <= _GEN_4747;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_126 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_126 <= _GEN_4748;
        end
      end
    end
    if (reset) begin // @[cache.scala 21:26]
      valid_0_127 <= 1'h0; // @[cache.scala 21:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_0_127 <= _GEN_4749;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_0 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_0 <= _GEN_5007;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_1 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_1 <= _GEN_5008;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_2 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_2 <= _GEN_5009;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_3 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_3 <= _GEN_5010;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_4 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_4 <= _GEN_5011;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_5 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_5 <= _GEN_5012;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_6 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_6 <= _GEN_5013;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_7 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_7 <= _GEN_5014;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_8 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_8 <= _GEN_5015;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_9 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_9 <= _GEN_5016;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_10 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_10 <= _GEN_5017;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_11 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_11 <= _GEN_5018;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_12 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_12 <= _GEN_5019;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_13 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_13 <= _GEN_5020;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_14 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_14 <= _GEN_5021;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_15 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_15 <= _GEN_5022;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_16 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_16 <= _GEN_5023;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_17 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_17 <= _GEN_5024;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_18 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_18 <= _GEN_5025;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_19 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_19 <= _GEN_5026;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_20 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_20 <= _GEN_5027;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_21 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_21 <= _GEN_5028;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_22 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_22 <= _GEN_5029;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_23 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_23 <= _GEN_5030;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_24 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_24 <= _GEN_5031;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_25 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_25 <= _GEN_5032;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_26 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_26 <= _GEN_5033;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_27 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_27 <= _GEN_5034;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_28 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_28 <= _GEN_5035;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_29 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_29 <= _GEN_5036;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_30 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_30 <= _GEN_5037;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_31 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_31 <= _GEN_5038;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_32 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_32 <= _GEN_5039;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_33 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_33 <= _GEN_5040;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_34 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_34 <= _GEN_5041;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_35 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_35 <= _GEN_5042;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_36 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_36 <= _GEN_5043;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_37 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_37 <= _GEN_5044;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_38 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_38 <= _GEN_5045;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_39 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_39 <= _GEN_5046;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_40 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_40 <= _GEN_5047;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_41 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_41 <= _GEN_5048;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_42 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_42 <= _GEN_5049;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_43 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_43 <= _GEN_5050;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_44 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_44 <= _GEN_5051;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_45 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_45 <= _GEN_5052;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_46 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_46 <= _GEN_5053;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_47 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_47 <= _GEN_5054;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_48 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_48 <= _GEN_5055;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_49 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_49 <= _GEN_5056;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_50 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_50 <= _GEN_5057;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_51 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_51 <= _GEN_5058;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_52 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_52 <= _GEN_5059;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_53 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_53 <= _GEN_5060;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_54 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_54 <= _GEN_5061;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_55 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_55 <= _GEN_5062;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_56 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_56 <= _GEN_5063;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_57 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_57 <= _GEN_5064;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_58 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_58 <= _GEN_5065;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_59 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_59 <= _GEN_5066;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_60 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_60 <= _GEN_5067;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_61 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_61 <= _GEN_5068;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_62 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_62 <= _GEN_5069;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_63 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_63 <= _GEN_5070;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_64 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_64 <= _GEN_5071;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_65 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_65 <= _GEN_5072;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_66 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_66 <= _GEN_5073;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_67 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_67 <= _GEN_5074;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_68 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_68 <= _GEN_5075;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_69 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_69 <= _GEN_5076;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_70 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_70 <= _GEN_5077;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_71 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_71 <= _GEN_5078;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_72 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_72 <= _GEN_5079;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_73 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_73 <= _GEN_5080;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_74 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_74 <= _GEN_5081;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_75 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_75 <= _GEN_5082;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_76 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_76 <= _GEN_5083;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_77 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_77 <= _GEN_5084;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_78 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_78 <= _GEN_5085;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_79 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_79 <= _GEN_5086;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_80 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_80 <= _GEN_5087;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_81 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_81 <= _GEN_5088;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_82 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_82 <= _GEN_5089;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_83 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_83 <= _GEN_5090;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_84 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_84 <= _GEN_5091;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_85 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_85 <= _GEN_5092;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_86 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_86 <= _GEN_5093;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_87 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_87 <= _GEN_5094;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_88 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_88 <= _GEN_5095;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_89 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_89 <= _GEN_5096;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_90 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_90 <= _GEN_5097;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_91 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_91 <= _GEN_5098;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_92 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_92 <= _GEN_5099;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_93 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_93 <= _GEN_5100;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_94 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_94 <= _GEN_5101;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_95 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_95 <= _GEN_5102;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_96 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_96 <= _GEN_5103;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_97 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_97 <= _GEN_5104;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_98 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_98 <= _GEN_5105;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_99 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_99 <= _GEN_5106;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_100 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_100 <= _GEN_5107;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_101 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_101 <= _GEN_5108;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_102 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_102 <= _GEN_5109;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_103 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_103 <= _GEN_5110;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_104 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_104 <= _GEN_5111;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_105 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_105 <= _GEN_5112;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_106 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_106 <= _GEN_5113;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_107 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_107 <= _GEN_5114;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_108 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_108 <= _GEN_5115;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_109 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_109 <= _GEN_5116;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_110 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_110 <= _GEN_5117;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_111 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_111 <= _GEN_5118;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_112 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_112 <= _GEN_5119;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_113 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_113 <= _GEN_5120;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_114 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_114 <= _GEN_5121;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_115 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_115 <= _GEN_5122;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_116 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_116 <= _GEN_5123;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_117 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_117 <= _GEN_5124;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_118 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_118 <= _GEN_5125;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_119 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_119 <= _GEN_5126;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_120 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_120 <= _GEN_5127;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_121 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_121 <= _GEN_5128;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_122 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_122 <= _GEN_5129;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_123 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_123 <= _GEN_5130;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_124 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_124 <= _GEN_5131;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_125 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_125 <= _GEN_5132;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_126 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_126 <= _GEN_5133;
        end
      end
    end
    if (reset) begin // @[cache.scala 22:26]
      valid_1_127 <= 1'h0; // @[cache.scala 22:26]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          valid_1_127 <= _GEN_5134;
        end
      end
    end
    if (reset) begin // @[cache.scala 23:27]
      way0_hit <= 1'h0; // @[cache.scala 23:27]
    end else begin
      way0_hit <= _GEN_256;
    end
    if (reset) begin // @[cache.scala 24:27]
      way1_hit <= 1'h0; // @[cache.scala 24:27]
    end else begin
      way1_hit <= _GEN_513;
    end
    if (reset) begin // @[cache.scala 26:28]
      unuse_way <= 2'h0; // @[cache.scala 26:28]
    end else if (~_GEN_255) begin // @[cache.scala 41:31]
      unuse_way <= 2'h1; // @[cache.scala 42:19]
    end else if (~_GEN_512) begin // @[cache.scala 43:37]
      unuse_way <= 2'h2; // @[cache.scala 44:19]
    end else begin
      unuse_way <= 2'h0; // @[cache.scala 46:19]
    end
    if (reset) begin // @[cache.scala 27:31]
      receive_data <= 64'h0; // @[cache.scala 27:31]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (2'h2 == state) begin // @[cache.scala 51:18]
          receive_data <= _GEN_521;
        end
      end
    end
    if (reset) begin // @[cache.scala 28:24]
      quene <= 1'h0; // @[cache.scala 28:24]
    end else if (!(2'h0 == state)) begin // @[cache.scala 51:18]
      if (!(2'h1 == state)) begin // @[cache.scala 51:18]
        if (!(2'h2 == state)) begin // @[cache.scala 51:18]
          quene <= _GEN_4750;
        end
      end
    end
    if (reset) begin // @[cache.scala 49:24]
      state <= 2'h0; // @[cache.scala 49:24]
    end else if (2'h0 == state) begin // @[cache.scala 51:18]
      if (io_from_ifu_arvalid) begin // @[cache.scala 53:38]
        state <= 2'h1; // @[cache.scala 54:23]
      end
    end else if (2'h1 == state) begin // @[cache.scala 51:18]
      if (way0_hit) begin // @[cache.scala 59:27]
        state <= _GEN_517;
      end else begin
        state <= _GEN_518;
      end
    end else if (2'h2 == state) begin // @[cache.scala 51:18]
      state <= _GEN_520;
    end else begin
      state <= _GEN_4365;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"enter cache\n"); // @[cache.scala 14:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"cache state:%d\n",state); // @[cache.scala 50:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ram_0_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ram_0_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ram_0_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ram_0_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ram_0_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ram_0_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ram_0_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ram_0_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  ram_0_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  ram_0_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  ram_0_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  ram_0_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  ram_0_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  ram_0_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  ram_0_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  ram_0_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  ram_0_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  ram_0_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  ram_0_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  ram_0_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  ram_0_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  ram_0_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  ram_0_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  ram_0_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  ram_0_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  ram_0_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  ram_0_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  ram_0_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  ram_0_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  ram_0_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  ram_0_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  ram_0_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  ram_0_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  ram_0_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  ram_0_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  ram_0_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ram_0_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  ram_0_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  ram_0_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  ram_0_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  ram_0_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  ram_0_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  ram_0_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  ram_0_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  ram_0_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  ram_0_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  ram_0_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  ram_0_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  ram_0_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  ram_0_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  ram_0_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  ram_0_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  ram_0_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  ram_0_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  ram_0_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  ram_0_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  ram_0_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  ram_0_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  ram_0_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  ram_0_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  ram_0_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  ram_0_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  ram_0_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  ram_0_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  ram_0_64 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  ram_0_65 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  ram_0_66 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  ram_0_67 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  ram_0_68 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  ram_0_69 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  ram_0_70 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  ram_0_71 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  ram_0_72 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  ram_0_73 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  ram_0_74 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  ram_0_75 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  ram_0_76 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  ram_0_77 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  ram_0_78 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  ram_0_79 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  ram_0_80 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  ram_0_81 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  ram_0_82 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  ram_0_83 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  ram_0_84 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  ram_0_85 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  ram_0_86 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  ram_0_87 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  ram_0_88 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  ram_0_89 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  ram_0_90 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  ram_0_91 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  ram_0_92 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  ram_0_93 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  ram_0_94 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  ram_0_95 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  ram_0_96 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  ram_0_97 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  ram_0_98 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  ram_0_99 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  ram_0_100 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  ram_0_101 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  ram_0_102 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  ram_0_103 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  ram_0_104 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  ram_0_105 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  ram_0_106 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  ram_0_107 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  ram_0_108 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  ram_0_109 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  ram_0_110 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  ram_0_111 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  ram_0_112 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  ram_0_113 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  ram_0_114 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  ram_0_115 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  ram_0_116 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  ram_0_117 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  ram_0_118 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  ram_0_119 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  ram_0_120 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  ram_0_121 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  ram_0_122 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  ram_0_123 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  ram_0_124 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  ram_0_125 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  ram_0_126 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  ram_0_127 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  ram_1_0 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  ram_1_1 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  ram_1_2 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  ram_1_3 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  ram_1_4 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  ram_1_5 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  ram_1_6 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  ram_1_7 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  ram_1_8 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  ram_1_9 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  ram_1_10 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  ram_1_11 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  ram_1_12 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  ram_1_13 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  ram_1_14 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  ram_1_15 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  ram_1_16 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  ram_1_17 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  ram_1_18 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  ram_1_19 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  ram_1_20 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  ram_1_21 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  ram_1_22 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  ram_1_23 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  ram_1_24 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  ram_1_25 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  ram_1_26 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  ram_1_27 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  ram_1_28 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  ram_1_29 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  ram_1_30 = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  ram_1_31 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  ram_1_32 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  ram_1_33 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  ram_1_34 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  ram_1_35 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  ram_1_36 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  ram_1_37 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  ram_1_38 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  ram_1_39 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  ram_1_40 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  ram_1_41 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  ram_1_42 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  ram_1_43 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  ram_1_44 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  ram_1_45 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  ram_1_46 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  ram_1_47 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  ram_1_48 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  ram_1_49 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  ram_1_50 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  ram_1_51 = _RAND_179[63:0];
  _RAND_180 = {2{`RANDOM}};
  ram_1_52 = _RAND_180[63:0];
  _RAND_181 = {2{`RANDOM}};
  ram_1_53 = _RAND_181[63:0];
  _RAND_182 = {2{`RANDOM}};
  ram_1_54 = _RAND_182[63:0];
  _RAND_183 = {2{`RANDOM}};
  ram_1_55 = _RAND_183[63:0];
  _RAND_184 = {2{`RANDOM}};
  ram_1_56 = _RAND_184[63:0];
  _RAND_185 = {2{`RANDOM}};
  ram_1_57 = _RAND_185[63:0];
  _RAND_186 = {2{`RANDOM}};
  ram_1_58 = _RAND_186[63:0];
  _RAND_187 = {2{`RANDOM}};
  ram_1_59 = _RAND_187[63:0];
  _RAND_188 = {2{`RANDOM}};
  ram_1_60 = _RAND_188[63:0];
  _RAND_189 = {2{`RANDOM}};
  ram_1_61 = _RAND_189[63:0];
  _RAND_190 = {2{`RANDOM}};
  ram_1_62 = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  ram_1_63 = _RAND_191[63:0];
  _RAND_192 = {2{`RANDOM}};
  ram_1_64 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  ram_1_65 = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  ram_1_66 = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  ram_1_67 = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  ram_1_68 = _RAND_196[63:0];
  _RAND_197 = {2{`RANDOM}};
  ram_1_69 = _RAND_197[63:0];
  _RAND_198 = {2{`RANDOM}};
  ram_1_70 = _RAND_198[63:0];
  _RAND_199 = {2{`RANDOM}};
  ram_1_71 = _RAND_199[63:0];
  _RAND_200 = {2{`RANDOM}};
  ram_1_72 = _RAND_200[63:0];
  _RAND_201 = {2{`RANDOM}};
  ram_1_73 = _RAND_201[63:0];
  _RAND_202 = {2{`RANDOM}};
  ram_1_74 = _RAND_202[63:0];
  _RAND_203 = {2{`RANDOM}};
  ram_1_75 = _RAND_203[63:0];
  _RAND_204 = {2{`RANDOM}};
  ram_1_76 = _RAND_204[63:0];
  _RAND_205 = {2{`RANDOM}};
  ram_1_77 = _RAND_205[63:0];
  _RAND_206 = {2{`RANDOM}};
  ram_1_78 = _RAND_206[63:0];
  _RAND_207 = {2{`RANDOM}};
  ram_1_79 = _RAND_207[63:0];
  _RAND_208 = {2{`RANDOM}};
  ram_1_80 = _RAND_208[63:0];
  _RAND_209 = {2{`RANDOM}};
  ram_1_81 = _RAND_209[63:0];
  _RAND_210 = {2{`RANDOM}};
  ram_1_82 = _RAND_210[63:0];
  _RAND_211 = {2{`RANDOM}};
  ram_1_83 = _RAND_211[63:0];
  _RAND_212 = {2{`RANDOM}};
  ram_1_84 = _RAND_212[63:0];
  _RAND_213 = {2{`RANDOM}};
  ram_1_85 = _RAND_213[63:0];
  _RAND_214 = {2{`RANDOM}};
  ram_1_86 = _RAND_214[63:0];
  _RAND_215 = {2{`RANDOM}};
  ram_1_87 = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  ram_1_88 = _RAND_216[63:0];
  _RAND_217 = {2{`RANDOM}};
  ram_1_89 = _RAND_217[63:0];
  _RAND_218 = {2{`RANDOM}};
  ram_1_90 = _RAND_218[63:0];
  _RAND_219 = {2{`RANDOM}};
  ram_1_91 = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  ram_1_92 = _RAND_220[63:0];
  _RAND_221 = {2{`RANDOM}};
  ram_1_93 = _RAND_221[63:0];
  _RAND_222 = {2{`RANDOM}};
  ram_1_94 = _RAND_222[63:0];
  _RAND_223 = {2{`RANDOM}};
  ram_1_95 = _RAND_223[63:0];
  _RAND_224 = {2{`RANDOM}};
  ram_1_96 = _RAND_224[63:0];
  _RAND_225 = {2{`RANDOM}};
  ram_1_97 = _RAND_225[63:0];
  _RAND_226 = {2{`RANDOM}};
  ram_1_98 = _RAND_226[63:0];
  _RAND_227 = {2{`RANDOM}};
  ram_1_99 = _RAND_227[63:0];
  _RAND_228 = {2{`RANDOM}};
  ram_1_100 = _RAND_228[63:0];
  _RAND_229 = {2{`RANDOM}};
  ram_1_101 = _RAND_229[63:0];
  _RAND_230 = {2{`RANDOM}};
  ram_1_102 = _RAND_230[63:0];
  _RAND_231 = {2{`RANDOM}};
  ram_1_103 = _RAND_231[63:0];
  _RAND_232 = {2{`RANDOM}};
  ram_1_104 = _RAND_232[63:0];
  _RAND_233 = {2{`RANDOM}};
  ram_1_105 = _RAND_233[63:0];
  _RAND_234 = {2{`RANDOM}};
  ram_1_106 = _RAND_234[63:0];
  _RAND_235 = {2{`RANDOM}};
  ram_1_107 = _RAND_235[63:0];
  _RAND_236 = {2{`RANDOM}};
  ram_1_108 = _RAND_236[63:0];
  _RAND_237 = {2{`RANDOM}};
  ram_1_109 = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  ram_1_110 = _RAND_238[63:0];
  _RAND_239 = {2{`RANDOM}};
  ram_1_111 = _RAND_239[63:0];
  _RAND_240 = {2{`RANDOM}};
  ram_1_112 = _RAND_240[63:0];
  _RAND_241 = {2{`RANDOM}};
  ram_1_113 = _RAND_241[63:0];
  _RAND_242 = {2{`RANDOM}};
  ram_1_114 = _RAND_242[63:0];
  _RAND_243 = {2{`RANDOM}};
  ram_1_115 = _RAND_243[63:0];
  _RAND_244 = {2{`RANDOM}};
  ram_1_116 = _RAND_244[63:0];
  _RAND_245 = {2{`RANDOM}};
  ram_1_117 = _RAND_245[63:0];
  _RAND_246 = {2{`RANDOM}};
  ram_1_118 = _RAND_246[63:0];
  _RAND_247 = {2{`RANDOM}};
  ram_1_119 = _RAND_247[63:0];
  _RAND_248 = {2{`RANDOM}};
  ram_1_120 = _RAND_248[63:0];
  _RAND_249 = {2{`RANDOM}};
  ram_1_121 = _RAND_249[63:0];
  _RAND_250 = {2{`RANDOM}};
  ram_1_122 = _RAND_250[63:0];
  _RAND_251 = {2{`RANDOM}};
  ram_1_123 = _RAND_251[63:0];
  _RAND_252 = {2{`RANDOM}};
  ram_1_124 = _RAND_252[63:0];
  _RAND_253 = {2{`RANDOM}};
  ram_1_125 = _RAND_253[63:0];
  _RAND_254 = {2{`RANDOM}};
  ram_1_126 = _RAND_254[63:0];
  _RAND_255 = {2{`RANDOM}};
  ram_1_127 = _RAND_255[63:0];
  _RAND_256 = {1{`RANDOM}};
  tag_0_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  tag_0_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  tag_0_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  tag_0_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  tag_0_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  tag_0_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  tag_0_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  tag_0_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  tag_0_8 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  tag_0_9 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  tag_0_10 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  tag_0_11 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  tag_0_12 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  tag_0_13 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  tag_0_14 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  tag_0_15 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  tag_0_16 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  tag_0_17 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  tag_0_18 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  tag_0_19 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  tag_0_20 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  tag_0_21 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  tag_0_22 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  tag_0_23 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  tag_0_24 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  tag_0_25 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  tag_0_26 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  tag_0_27 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  tag_0_28 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  tag_0_29 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  tag_0_30 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  tag_0_31 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  tag_0_32 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  tag_0_33 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  tag_0_34 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  tag_0_35 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  tag_0_36 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  tag_0_37 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  tag_0_38 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  tag_0_39 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  tag_0_40 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  tag_0_41 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  tag_0_42 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  tag_0_43 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  tag_0_44 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  tag_0_45 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  tag_0_46 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  tag_0_47 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  tag_0_48 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  tag_0_49 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  tag_0_50 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  tag_0_51 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  tag_0_52 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  tag_0_53 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  tag_0_54 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  tag_0_55 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  tag_0_56 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  tag_0_57 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  tag_0_58 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  tag_0_59 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  tag_0_60 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  tag_0_61 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  tag_0_62 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  tag_0_63 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  tag_0_64 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  tag_0_65 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  tag_0_66 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  tag_0_67 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  tag_0_68 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  tag_0_69 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  tag_0_70 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  tag_0_71 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  tag_0_72 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  tag_0_73 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  tag_0_74 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  tag_0_75 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  tag_0_76 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  tag_0_77 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  tag_0_78 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  tag_0_79 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  tag_0_80 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  tag_0_81 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  tag_0_82 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  tag_0_83 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  tag_0_84 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  tag_0_85 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  tag_0_86 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  tag_0_87 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  tag_0_88 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  tag_0_89 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  tag_0_90 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  tag_0_91 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  tag_0_92 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  tag_0_93 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  tag_0_94 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  tag_0_95 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  tag_0_96 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  tag_0_97 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  tag_0_98 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  tag_0_99 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  tag_0_100 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  tag_0_101 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  tag_0_102 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  tag_0_103 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  tag_0_104 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  tag_0_105 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  tag_0_106 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  tag_0_107 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  tag_0_108 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  tag_0_109 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  tag_0_110 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  tag_0_111 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  tag_0_112 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  tag_0_113 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  tag_0_114 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  tag_0_115 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  tag_0_116 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  tag_0_117 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  tag_0_118 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  tag_0_119 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  tag_0_120 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  tag_0_121 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  tag_0_122 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  tag_0_123 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  tag_0_124 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  tag_0_125 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  tag_0_126 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  tag_0_127 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  tag_1_0 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  tag_1_1 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  tag_1_2 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  tag_1_3 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  tag_1_4 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  tag_1_5 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  tag_1_6 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  tag_1_7 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  tag_1_8 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  tag_1_9 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  tag_1_10 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  tag_1_11 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  tag_1_12 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  tag_1_13 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  tag_1_14 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  tag_1_15 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  tag_1_16 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  tag_1_17 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  tag_1_18 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  tag_1_19 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  tag_1_20 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  tag_1_21 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  tag_1_22 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  tag_1_23 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  tag_1_24 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  tag_1_25 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  tag_1_26 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  tag_1_27 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  tag_1_28 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  tag_1_29 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  tag_1_30 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  tag_1_31 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  tag_1_32 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  tag_1_33 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  tag_1_34 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  tag_1_35 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  tag_1_36 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  tag_1_37 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  tag_1_38 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  tag_1_39 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  tag_1_40 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  tag_1_41 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  tag_1_42 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  tag_1_43 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  tag_1_44 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  tag_1_45 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  tag_1_46 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  tag_1_47 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  tag_1_48 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  tag_1_49 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  tag_1_50 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  tag_1_51 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  tag_1_52 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  tag_1_53 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  tag_1_54 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  tag_1_55 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  tag_1_56 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  tag_1_57 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  tag_1_58 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  tag_1_59 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  tag_1_60 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  tag_1_61 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  tag_1_62 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  tag_1_63 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  tag_1_64 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  tag_1_65 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  tag_1_66 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  tag_1_67 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  tag_1_68 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  tag_1_69 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  tag_1_70 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  tag_1_71 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  tag_1_72 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  tag_1_73 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  tag_1_74 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  tag_1_75 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  tag_1_76 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  tag_1_77 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  tag_1_78 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  tag_1_79 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  tag_1_80 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  tag_1_81 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  tag_1_82 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  tag_1_83 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  tag_1_84 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  tag_1_85 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  tag_1_86 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  tag_1_87 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  tag_1_88 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  tag_1_89 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  tag_1_90 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  tag_1_91 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  tag_1_92 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  tag_1_93 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  tag_1_94 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  tag_1_95 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  tag_1_96 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  tag_1_97 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  tag_1_98 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  tag_1_99 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  tag_1_100 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  tag_1_101 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  tag_1_102 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  tag_1_103 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  tag_1_104 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  tag_1_105 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  tag_1_106 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  tag_1_107 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  tag_1_108 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  tag_1_109 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  tag_1_110 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  tag_1_111 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  tag_1_112 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  tag_1_113 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  tag_1_114 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  tag_1_115 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  tag_1_116 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  tag_1_117 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  tag_1_118 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  tag_1_119 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  tag_1_120 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  tag_1_121 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  tag_1_122 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  tag_1_123 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  tag_1_124 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  tag_1_125 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  tag_1_126 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  tag_1_127 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  valid_0_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_0_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_0_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_0_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_0_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_0_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_0_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_0_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_0_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_0_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_0_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_0_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_0_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_0_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_0_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_0_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  valid_0_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  valid_0_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  valid_0_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  valid_0_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  valid_0_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  valid_0_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  valid_0_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  valid_0_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  valid_0_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  valid_0_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  valid_0_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  valid_0_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  valid_0_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  valid_0_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  valid_0_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  valid_0_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  valid_0_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  valid_0_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  valid_0_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  valid_0_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  valid_0_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  valid_0_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  valid_0_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  valid_0_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  valid_0_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  valid_0_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  valid_0_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  valid_0_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  valid_0_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  valid_0_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  valid_0_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  valid_0_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  valid_0_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  valid_0_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  valid_0_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  valid_0_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  valid_0_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  valid_0_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  valid_0_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  valid_0_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  valid_0_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  valid_0_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  valid_0_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  valid_0_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  valid_0_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  valid_0_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  valid_0_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  valid_0_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  valid_0_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_0_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_0_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_0_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_0_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_0_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_0_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_0_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_0_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_0_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_0_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_0_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_0_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_0_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_0_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_0_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_0_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_0_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_0_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_0_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_0_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_0_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_0_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_0_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_0_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_0_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_0_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_0_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_0_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_0_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_0_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_0_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_0_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_0_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_0_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_0_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_0_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_0_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_0_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_0_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_0_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_0_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_0_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_0_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_0_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_0_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_0_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_0_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_0_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_0_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_0_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_0_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_0_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_0_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_0_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_0_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_0_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_0_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_0_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_0_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_0_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_0_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_0_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_0_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  valid_1_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  valid_1_1 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  valid_1_2 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  valid_1_3 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  valid_1_4 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  valid_1_5 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  valid_1_6 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  valid_1_7 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  valid_1_8 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  valid_1_9 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  valid_1_10 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  valid_1_11 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  valid_1_12 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  valid_1_13 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  valid_1_14 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  valid_1_15 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  valid_1_16 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  valid_1_17 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  valid_1_18 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  valid_1_19 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  valid_1_20 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  valid_1_21 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  valid_1_22 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  valid_1_23 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  valid_1_24 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  valid_1_25 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  valid_1_26 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  valid_1_27 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  valid_1_28 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  valid_1_29 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  valid_1_30 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  valid_1_31 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  valid_1_32 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  valid_1_33 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  valid_1_34 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  valid_1_35 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  valid_1_36 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  valid_1_37 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  valid_1_38 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  valid_1_39 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  valid_1_40 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  valid_1_41 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  valid_1_42 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  valid_1_43 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  valid_1_44 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  valid_1_45 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  valid_1_46 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  valid_1_47 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  valid_1_48 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  valid_1_49 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  valid_1_50 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  valid_1_51 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  valid_1_52 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  valid_1_53 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  valid_1_54 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  valid_1_55 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  valid_1_56 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  valid_1_57 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  valid_1_58 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  valid_1_59 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  valid_1_60 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  valid_1_61 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  valid_1_62 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  valid_1_63 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  valid_1_64 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  valid_1_65 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  valid_1_66 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  valid_1_67 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  valid_1_68 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  valid_1_69 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  valid_1_70 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  valid_1_71 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  valid_1_72 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  valid_1_73 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  valid_1_74 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  valid_1_75 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  valid_1_76 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  valid_1_77 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  valid_1_78 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  valid_1_79 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  valid_1_80 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  valid_1_81 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  valid_1_82 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  valid_1_83 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  valid_1_84 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  valid_1_85 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  valid_1_86 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  valid_1_87 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  valid_1_88 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  valid_1_89 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  valid_1_90 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  valid_1_91 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  valid_1_92 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  valid_1_93 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  valid_1_94 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  valid_1_95 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  valid_1_96 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  valid_1_97 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  valid_1_98 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  valid_1_99 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  valid_1_100 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  valid_1_101 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  valid_1_102 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  valid_1_103 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  valid_1_104 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  valid_1_105 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  valid_1_106 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  valid_1_107 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  valid_1_108 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  valid_1_109 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  valid_1_110 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  valid_1_111 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  valid_1_112 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  valid_1_113 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  valid_1_114 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  valid_1_115 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  valid_1_116 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  valid_1_117 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  valid_1_118 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  valid_1_119 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  valid_1_120 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  valid_1_121 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  valid_1_122 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  valid_1_123 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  valid_1_124 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  valid_1_125 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  valid_1_126 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  valid_1_127 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  way0_hit = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  way1_hit = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  unuse_way = _RAND_770[1:0];
  _RAND_771 = {2{`RANDOM}};
  receive_data = _RAND_771[63:0];
  _RAND_772 = {1{`RANDOM}};
  quene = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  state = _RAND_773[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDU(
  input  [31:0] io_inst,
  output [31:0] io_inst_now,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  output [4:0]  io_rd,
  output [63:0] io_imm,
  output        io_ctrl_sign_reg_write,
  output        io_ctrl_sign_csr_write,
  output        io_ctrl_sign_src2_is_imm,
  output        io_ctrl_sign_src1_is_pc,
  output        io_ctrl_sign_Writemem_en,
  output        io_ctrl_sign_Readmem_en,
  output [7:0]  io_ctrl_sign_Wmask
);
  wire [4:0] rd = io_inst[11:7]; // @[IDU.scala 150:15]
  wire [31:0] _inst_type_T = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_1 = 32'h13 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_2 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_3 = 32'h17 == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_5 = 32'h37 == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_7 = 32'h6f == _inst_type_T_2; // @[Lookup.scala 31:38]
  wire  _inst_type_T_9 = 32'h67 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_11 = 32'h3023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_13 = 32'h3013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_15 = 32'h2003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_16 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_17 = 32'h3b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_19 = 32'h40000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_21 = 32'h1063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_23 = 32'h63 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_25 = 32'h3003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_27 = 32'h1b == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_29 = 32'h33 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_30 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_31 = 32'h40005013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_33 = 32'h4003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_35 = 32'h1023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_37 = 32'h23 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_39 = 32'h6033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_41 = 32'h4013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_43 = 32'h7033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_45 = 32'h7013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_47 = 32'h4000003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_49 = 32'h103b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_51 = 32'h1013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_53 = 32'h5013 == _inst_type_T_30; // @[Lookup.scala 31:38]
  wire  _inst_type_T_55 = 32'h101b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_57 = 32'h4000501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_59 = 32'h501b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_61 = 32'h4000503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_63 = 32'h503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_65 = 32'h3033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_67 = 32'h2033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_69 = 32'h5063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_71 = 32'h4063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_73 = 32'h6063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_75 = 32'h2023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_77 = 32'h1003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_79 = 32'h5003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_81 = 32'h2000033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_83 = 32'h200003b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_85 = 32'h200403b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_87 = 32'h200603b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_89 = 32'h4033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_91 = 32'h6013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_93 = 32'h2005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_95 = 32'h2004033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_97 = 32'h200503b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_99 = 32'h200703b == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_101 = 32'h2007033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_103 = 32'h2006033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_105 = 32'h1033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_107 = 32'h5033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_109 = 32'h40005033 == _inst_type_T_16; // @[Lookup.scala 31:38]
  wire  _inst_type_T_111 = 32'h2013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_113 = 32'h6003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_115 = 32'h3 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_117 = 32'h7063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_119 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _inst_type_T_121 = 32'h1073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_123 = 32'h2073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_125 = 32'h3073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [6:0] _inst_type_T_126 = _inst_type_T_125 ? 7'h40 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_127 = _inst_type_T_123 ? 7'h40 : _inst_type_T_126; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_128 = _inst_type_T_121 ? 7'h40 : _inst_type_T_127; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_129 = _inst_type_T_119 ? 7'h40 : _inst_type_T_128; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_130 = _inst_type_T_117 ? 7'h45 : _inst_type_T_129; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_131 = _inst_type_T_115 ? 7'h40 : _inst_type_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_132 = _inst_type_T_113 ? 7'h40 : _inst_type_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_133 = _inst_type_T_111 ? 7'h40 : _inst_type_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_134 = _inst_type_T_109 ? 7'h41 : _inst_type_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_135 = _inst_type_T_107 ? 7'h41 : _inst_type_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_136 = _inst_type_T_105 ? 7'h41 : _inst_type_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_137 = _inst_type_T_103 ? 7'h41 : _inst_type_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_138 = _inst_type_T_101 ? 7'h41 : _inst_type_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_139 = _inst_type_T_99 ? 7'h41 : _inst_type_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_140 = _inst_type_T_97 ? 7'h41 : _inst_type_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_141 = _inst_type_T_95 ? 7'h41 : _inst_type_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_142 = _inst_type_T_93 ? 7'h41 : _inst_type_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_143 = _inst_type_T_91 ? 7'h40 : _inst_type_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_144 = _inst_type_T_89 ? 7'h41 : _inst_type_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_145 = _inst_type_T_87 ? 7'h41 : _inst_type_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_146 = _inst_type_T_85 ? 7'h41 : _inst_type_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_147 = _inst_type_T_83 ? 7'h41 : _inst_type_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_148 = _inst_type_T_81 ? 7'h41 : _inst_type_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_149 = _inst_type_T_79 ? 7'h40 : _inst_type_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_150 = _inst_type_T_77 ? 7'h40 : _inst_type_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_151 = _inst_type_T_75 ? 7'h44 : _inst_type_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_152 = _inst_type_T_73 ? 7'h45 : _inst_type_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_153 = _inst_type_T_71 ? 7'h45 : _inst_type_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_154 = _inst_type_T_69 ? 7'h45 : _inst_type_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_155 = _inst_type_T_67 ? 7'h41 : _inst_type_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_156 = _inst_type_T_65 ? 7'h41 : _inst_type_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_157 = _inst_type_T_63 ? 7'h41 : _inst_type_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_158 = _inst_type_T_61 ? 7'h41 : _inst_type_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_159 = _inst_type_T_59 ? 7'h40 : _inst_type_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_160 = _inst_type_T_57 ? 7'h40 : _inst_type_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_161 = _inst_type_T_55 ? 7'h40 : _inst_type_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_162 = _inst_type_T_53 ? 7'h40 : _inst_type_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_163 = _inst_type_T_51 ? 7'h40 : _inst_type_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_164 = _inst_type_T_49 ? 7'h41 : _inst_type_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_165 = _inst_type_T_47 ? 7'h41 : _inst_type_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_166 = _inst_type_T_45 ? 7'h40 : _inst_type_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_167 = _inst_type_T_43 ? 7'h41 : _inst_type_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_168 = _inst_type_T_41 ? 7'h40 : _inst_type_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_169 = _inst_type_T_39 ? 7'h41 : _inst_type_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_170 = _inst_type_T_37 ? 7'h44 : _inst_type_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_171 = _inst_type_T_35 ? 7'h44 : _inst_type_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_172 = _inst_type_T_33 ? 7'h40 : _inst_type_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_173 = _inst_type_T_31 ? 7'h40 : _inst_type_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_174 = _inst_type_T_29 ? 7'h41 : _inst_type_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_175 = _inst_type_T_27 ? 7'h40 : _inst_type_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_176 = _inst_type_T_25 ? 7'h40 : _inst_type_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_177 = _inst_type_T_23 ? 7'h45 : _inst_type_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_178 = _inst_type_T_21 ? 7'h45 : _inst_type_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_179 = _inst_type_T_19 ? 7'h41 : _inst_type_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_180 = _inst_type_T_17 ? 7'h41 : _inst_type_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_181 = _inst_type_T_15 ? 7'h40 : _inst_type_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_182 = _inst_type_T_13 ? 7'h40 : _inst_type_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_183 = _inst_type_T_11 ? 7'h44 : _inst_type_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_184 = _inst_type_T_9 ? 7'h40 : _inst_type_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_185 = _inst_type_T_7 ? 7'h43 : _inst_type_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_186 = _inst_type_T_5 ? 7'h42 : _inst_type_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_187 = _inst_type_T_3 ? 7'h42 : _inst_type_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_type_T_188 = _inst_type_T_1 ? 7'h40 : _inst_type_T_187; // @[Lookup.scala 34:39]
  wire [11:0] imm_imm = io_inst[31:20]; // @[IDU.scala 24:23]
  wire [51:0] _imm_T_2 = imm_imm[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_3 = {_imm_T_2,imm_imm}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_1 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21]}; // @[Cat.scala 31:58]
  wire [42:0] _imm_T_6 = imm_imm_1[19] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_7 = {_imm_T_6,io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 31:58]
  wire [19:0] imm_imm_2 = io_inst[31:12]; // @[IDU.scala 28:23]
  wire [31:0] _imm_T_10 = imm_imm_2[19] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_12 = {_imm_T_10,imm_imm_2,12'h0}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_3 = {io_inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [51:0] _imm_T_15 = imm_imm_3[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_16 = {_imm_T_15,io_inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [11:0] imm_imm_4 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8]}; // @[Cat.scala 31:58]
  wire [50:0] _imm_T_19 = imm_imm_4[11] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _imm_T_20 = {_imm_T_19,io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] inst_type = {{25'd0}, _inst_type_T_188}; // @[IDU.scala 133:25 152:15]
  wire [63:0] _imm_T_22 = 32'h40 == inst_type ? _imm_T_3 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_24 = 32'h43 == inst_type ? _imm_T_7 : _imm_T_22; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_26 = 32'h42 == inst_type ? _imm_T_12 : _imm_T_24; // @[Mux.scala 81:58]
  wire [63:0] _imm_T_28 = 32'h44 == inst_type ? _imm_T_16 : _imm_T_26; // @[Mux.scala 81:58]
  wire  _inst_now_T_3 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  wire  _inst_now_T_123 = 32'h30200073 == io_inst; // @[Lookup.scala 31:38]
  wire [6:0] _inst_now_T_130 = _inst_type_T_125 ? 7'h47 : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_131 = _inst_type_T_123 ? 7'h46 : _inst_now_T_130; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_132 = _inst_type_T_121 ? 7'h3f : _inst_now_T_131; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_133 = _inst_now_T_123 ? 7'h3e : _inst_now_T_132; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_134 = _inst_type_T_119 ? 7'h3d : _inst_now_T_133; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_135 = _inst_type_T_117 ? 7'h3c : _inst_now_T_134; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_136 = _inst_type_T_115 ? 7'h3b : _inst_now_T_135; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_137 = _inst_type_T_113 ? 7'h3a : _inst_now_T_136; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_138 = _inst_type_T_111 ? 7'h36 : _inst_now_T_137; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_139 = _inst_type_T_109 ? 7'h39 : _inst_now_T_138; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_140 = _inst_type_T_107 ? 7'h38 : _inst_now_T_139; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_141 = _inst_type_T_105 ? 7'h37 : _inst_now_T_140; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_142 = _inst_type_T_103 ? 7'h34 : _inst_now_T_141; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_143 = _inst_type_T_101 ? 7'h33 : _inst_now_T_142; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_144 = _inst_type_T_99 ? 7'h32 : _inst_now_T_143; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_145 = _inst_type_T_97 ? 7'h35 : _inst_now_T_144; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_146 = _inst_type_T_95 ? 7'h31 : _inst_now_T_145; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_147 = _inst_type_T_93 ? 7'h30 : _inst_now_T_146; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_148 = _inst_type_T_91 ? 7'h2f : _inst_now_T_147; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_149 = _inst_type_T_89 ? 7'h2e : _inst_now_T_148; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_150 = _inst_type_T_87 ? 7'h14 : _inst_now_T_149; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_151 = _inst_type_T_85 ? 7'h13 : _inst_now_T_150; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_152 = _inst_type_T_83 ? 7'h12 : _inst_now_T_151; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_153 = _inst_type_T_81 ? 7'h11 : _inst_now_T_152; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_154 = _inst_type_T_79 ? 7'h25 : _inst_now_T_153; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_155 = _inst_type_T_77 ? 7'h24 : _inst_now_T_154; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_156 = _inst_type_T_75 ? 7'h27 : _inst_now_T_155; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_157 = _inst_type_T_73 ? 7'h2d : _inst_now_T_156; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_158 = _inst_type_T_71 ? 7'h2c : _inst_now_T_157; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_159 = _inst_type_T_69 ? 7'h2b : _inst_now_T_158; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_160 = _inst_type_T_67 ? 7'h1f : _inst_now_T_159; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_161 = _inst_type_T_65 ? 7'h1e : _inst_now_T_160; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_162 = _inst_type_T_63 ? 7'h1d : _inst_now_T_161; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_163 = _inst_type_T_61 ? 7'h1c : _inst_now_T_162; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_164 = _inst_type_T_59 ? 7'h1b : _inst_now_T_163; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_165 = _inst_type_T_57 ? 7'h1a : _inst_now_T_164; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_166 = _inst_type_T_55 ? 7'h19 : _inst_now_T_165; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_167 = _inst_type_T_53 ? 7'h18 : _inst_now_T_166; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_168 = _inst_type_T_51 ? 7'h17 : _inst_now_T_167; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_169 = _inst_type_T_49 ? 7'h16 : _inst_now_T_168; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_170 = _inst_type_T_47 ? 7'hd : _inst_now_T_169; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_171 = _inst_type_T_45 ? 7'h9 : _inst_now_T_170; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_172 = _inst_type_T_43 ? 7'h8 : _inst_now_T_171; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_173 = _inst_type_T_41 ? 7'ha : _inst_now_T_172; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_174 = _inst_type_T_39 ? 7'hb : _inst_now_T_173; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_175 = _inst_type_T_37 ? 7'h28 : _inst_now_T_174; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_176 = _inst_type_T_35 ? 7'h26 : _inst_now_T_175; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_177 = _inst_type_T_33 ? 7'h23 : _inst_now_T_176; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_178 = _inst_type_T_31 ? 7'h15 : _inst_now_T_177; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_179 = _inst_type_T_29 ? 7'hf : _inst_now_T_178; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_180 = _inst_type_T_27 ? 7'h10 : _inst_now_T_179; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_181 = _inst_type_T_25 ? 7'h22 : _inst_now_T_180; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_182 = _inst_type_T_23 ? 7'h29 : _inst_now_T_181; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_183 = _inst_type_T_21 ? 7'h2a : _inst_now_T_182; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_184 = _inst_type_T_19 ? 7'he : _inst_now_T_183; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_185 = _inst_type_T_17 ? 7'hc : _inst_now_T_184; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_186 = _inst_type_T_15 ? 7'h21 : _inst_now_T_185; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_187 = _inst_type_T_13 ? 7'h20 : _inst_now_T_186; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_188 = _inst_type_T_11 ? 7'h7 : _inst_now_T_187; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_189 = _inst_type_T_9 ? 7'h6 : _inst_now_T_188; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_190 = _inst_type_T_7 ? 7'h5 : _inst_now_T_189; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_191 = _inst_type_T_5 ? 7'h4 : _inst_now_T_190; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_192 = _inst_type_T_3 ? 7'h3 : _inst_now_T_191; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_193 = _inst_now_T_3 ? 7'h2 : _inst_now_T_192; // @[Lookup.scala 34:39]
  wire [6:0] _inst_now_T_194 = _inst_type_T_1 ? 7'h1 : _inst_now_T_193; // @[Lookup.scala 34:39]
  wire  _reg_write_T_26 = _inst_now_T_123 ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _reg_write_T_27 = _inst_type_T_119 ? 1'h0 : _reg_write_T_26; // @[Lookup.scala 34:39]
  wire  _reg_write_T_28 = _inst_type_T_117 ? 1'h0 : _reg_write_T_27; // @[Lookup.scala 34:39]
  wire  _reg_write_T_29 = _inst_type_T_73 ? 1'h0 : _reg_write_T_28; // @[Lookup.scala 34:39]
  wire  _reg_write_T_30 = _inst_type_T_71 ? 1'h0 : _reg_write_T_29; // @[Lookup.scala 34:39]
  wire  _reg_write_T_31 = _inst_type_T_69 ? 1'h0 : _reg_write_T_30; // @[Lookup.scala 34:39]
  wire  _reg_write_T_32 = _inst_type_T_23 ? 1'h0 : _reg_write_T_31; // @[Lookup.scala 34:39]
  wire  _reg_write_T_33 = _inst_type_T_21 ? 1'h0 : _reg_write_T_32; // @[Lookup.scala 34:39]
  wire  _reg_write_T_34 = _inst_type_T_75 ? 1'h0 : _reg_write_T_33; // @[Lookup.scala 34:39]
  wire  _reg_write_T_35 = _inst_type_T_37 ? 1'h0 : _reg_write_T_34; // @[Lookup.scala 34:39]
  wire  _reg_write_T_36 = _inst_type_T_35 ? 1'h0 : _reg_write_T_35; // @[Lookup.scala 34:39]
  wire  _reg_write_T_37 = _inst_type_T_11 ? 1'h0 : _reg_write_T_36; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_8 = _inst_type_T_75 ? 4'hf : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_9 = _inst_type_T_37 ? 4'h1 : _Wmask_T_8; // @[Lookup.scala 34:39]
  wire [3:0] _Wmask_T_10 = _inst_type_T_35 ? 4'h3 : _Wmask_T_9; // @[Lookup.scala 34:39]
  assign io_inst_now = {{25'd0}, _inst_now_T_194}; // @[IDU.scala 132:24 226:14]
  assign io_rs1 = io_inst[19:15]; // @[IDU.scala 149:16]
  assign io_rs2 = io_inst[24:20]; // @[IDU.scala 148:16]
  assign io_rd = io_inst[11:7]; // @[IDU.scala 150:15]
  assign io_imm = 32'h45 == inst_type ? _imm_T_20 : _imm_T_28; // @[Mux.scala 81:58]
  assign io_ctrl_sign_reg_write = _inst_now_T_3 ? 1'h0 : _reg_write_T_37; // @[Lookup.scala 34:39]
  assign io_ctrl_sign_csr_write = _inst_type_T_121 | (_inst_type_T_123 | _inst_type_T_125); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_src2_is_imm = 32'h45 == inst_type | (32'h43 == inst_type | (32'h44 == inst_type | (32'h42 ==
    inst_type | 32'h40 == inst_type))); // @[Mux.scala 81:58]
  assign io_ctrl_sign_src1_is_pc = _inst_type_T_7 | (_inst_type_T_3 | (_inst_type_T_21 | (_inst_type_T_23 | (
    _inst_type_T_69 | (_inst_type_T_71 | (_inst_type_T_73 | _inst_type_T_117)))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Writemem_en = 32'h44 == inst_type; // @[Mux.scala 81:61]
  assign io_ctrl_sign_Readmem_en = _inst_type_T_25 | (_inst_type_T_15 | (_inst_type_T_113 | (_inst_type_T_77 | (
    _inst_type_T_79 | (_inst_type_T_115 | _inst_type_T_33))))); // @[Lookup.scala 34:39]
  assign io_ctrl_sign_Wmask = _inst_type_T_11 ? 8'hff : {{4'd0}, _Wmask_T_10}; // @[Lookup.scala 34:39]
endmodule
module EXU_AXI(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  output [63:0] io_pc_next,
  input  [31:0] io_inst_now,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd,
  input  [63:0] io_imm,
  input         io_ctrl_sign_reg_write,
  input         io_ctrl_sign_csr_write,
  input         io_ctrl_sign_src2_is_imm,
  input         io_ctrl_sign_src1_is_pc,
  input         io_ctrl_sign_Writemem_en,
  input         io_ctrl_sign_Readmem_en,
  input  [7:0]  io_ctrl_sign_Wmask,
  output [63:0] io_res2rd,
  input         io_inst_valid,
  output        io_inst_store,
  output        io_inst_load,
  output [31:0] io_Mem_addr,
  input  [63:0] io_Mem_rdata,
  output [63:0] io_Mem_wdata,
  output [7:0]  io_Mem_wstrb,
  input         io_rdata_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] Regfile [0:31]; // @[EXU_AXI.scala 37:22]
  wire  Regfile_src1_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_src1_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_src1_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_src2_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_src2_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_src2_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_value_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_value_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_value_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_4_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_MPORT_4_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_MPORT_4_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_1_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_1_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_1_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_2_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_2_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_2_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_3_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_3_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_3_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_4_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_4_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_4_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_5_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_5_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_5_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_6_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_6_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_6_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_7_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_7_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_7_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_8_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_8_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_8_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_9_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_9_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_9_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_10_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_10_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_10_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_j_pc_MPORT_11_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_j_pc_MPORT_11_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_j_pc_MPORT_11_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_0_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_0_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_0_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_1_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_1_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_1_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_2_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_2_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_2_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_3_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_3_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_3_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_4_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_4_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_4_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_5_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_5_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_5_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_6_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_6_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_6_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_7_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_7_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_7_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_8_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_8_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_8_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_9_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_9_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_9_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_10_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_10_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_10_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_11_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_11_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_11_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_12_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_12_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_12_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_13_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_13_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_13_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_14_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_14_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_14_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_15_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_15_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_15_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_16_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_16_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_16_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_17_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_17_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_17_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_18_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_18_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_18_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_19_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_19_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_19_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_20_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_20_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_20_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_21_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_21_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_21_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_22_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_22_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_22_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_23_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_23_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_23_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_24_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_24_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_24_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_25_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_25_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_25_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_26_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_26_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_26_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_27_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_27_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_27_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_28_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_28_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_28_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_29_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_29_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_29_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_30_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_30_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_30_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_reg_trace_io_input_reg_31_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_reg_trace_io_input_reg_31_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_reg_trace_io_input_reg_31_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_1_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_1_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_1_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_2_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_2_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_2_data; // @[EXU_AXI.scala 37:22]
  wire  Regfile_mem_wdata_MPORT_3_en; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_mem_wdata_MPORT_3_addr; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_mem_wdata_MPORT_3_data; // @[EXU_AXI.scala 37:22]
  wire [63:0] Regfile_MPORT_data; // @[EXU_AXI.scala 37:22]
  wire [4:0] Regfile_MPORT_addr; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_mask; // @[EXU_AXI.scala 37:22]
  wire  Regfile_MPORT_en; // @[EXU_AXI.scala 37:22]
  reg [63:0] CSR_Reg [0:3]; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_io_res2rd_MPORT_2_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_io_res2rd_MPORT_2_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_io_res2rd_MPORT_2_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_csr_wdata_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_csr_wdata_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_csr_wdata_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_csr_wdata_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_csr_wdata_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_csr_wdata_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_2_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_2_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_2_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_5_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_5_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_5_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_7_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_7_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_7_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_j_pc_MPORT_12_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_j_pc_MPORT_12_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_j_pc_MPORT_12_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_j_pc_MPORT_13_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_j_pc_MPORT_13_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_j_pc_MPORT_13_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_0_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_1_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_reg_trace_io_csr_reg_2_MPORT_en; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_1_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_1_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_1_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_1_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_3_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_3_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_3_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_3_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] CSR_Reg_MPORT_6_data; // @[EXU_AXI.scala 38:22]
  wire [1:0] CSR_Reg_MPORT_6_addr; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_6_mask; // @[EXU_AXI.scala 38:22]
  wire  CSR_Reg_MPORT_6_en; // @[EXU_AXI.scala 38:22]
  wire [63:0] reg_trace_input_reg_0; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_1; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_2; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_3; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_4; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_5; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_6; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_7; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_8; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_9; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_10; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_11; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_12; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_13; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_14; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_15; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_16; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_17; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_18; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_19; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_20; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_21; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_22; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_23; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_24; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_25; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_26; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_27; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_28; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_29; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_30; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_input_reg_31; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_0; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_1; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_2; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_csr_reg_3; // @[EXU_AXI.scala 163:27]
  wire [63:0] reg_trace_pc; // @[EXU_AXI.scala 163:27]
  wire [11:0] csr_addr = io_imm[11:0]; // @[EXU_AXI.scala 39:26]
  wire [1:0] _csr_index_T_5 = 12'h300 == csr_addr ? 2'h2 : {{1'd0}, 12'h341 == csr_addr}; // @[Mux.scala 81:58]
  wire  _csr_index_T_6 = 12'h342 == csr_addr; // @[Mux.scala 81:61]
  wire [63:0] _src1_value_T_1 = io_rs1 == 5'h0 ? 64'h0 : Regfile_src1_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] src1_value = io_ctrl_sign_src1_is_pc ? io_pc : _src1_value_T_1; // @[EXU_AXI.scala 49:25]
  wire [63:0] _src2_value_T_1 = io_rs2 == 5'h0 ? 64'h0 : Regfile_src2_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] src2_value = io_ctrl_sign_src2_is_imm ? io_imm : _src2_value_T_1; // @[EXU_AXI.scala 50:25]
  wire [63:0] add_res = src1_value + src2_value; // @[EXU_AXI.scala 51:30]
  wire [63:0] sub_res = src1_value - src2_value; // @[EXU_AXI.scala 52:30]
  wire [63:0] _sra_res_T = io_ctrl_sign_src1_is_pc ? io_pc : _src1_value_T_1; // @[EXU_AXI.scala 53:37]
  wire [63:0] sra_res = $signed(_sra_res_T) >>> src2_value[5:0]; // @[EXU_AXI.scala 53:60]
  wire [63:0] srl_res = src1_value >> src2_value[5:0]; // @[EXU_AXI.scala 54:30]
  wire [126:0] _GEN_1 = {{63'd0}, src1_value}; // @[EXU_AXI.scala 55:30]
  wire [126:0] sll_res = _GEN_1 << src2_value[5:0]; // @[EXU_AXI.scala 55:30]
  wire [31:0] _sraw_res_T_1 = src1_value[31:0]; // @[EXU_AXI.scala 56:43]
  wire [31:0] sraw_res = $signed(_sraw_res_T_1) >>> src2_value[4:0]; // @[EXU_AXI.scala 56:46]
  wire [31:0] srlw_res = src1_value[31:0] >> src2_value[4:0]; // @[EXU_AXI.scala 57:37]
  wire [62:0] _GEN_2 = {{31'd0}, src1_value[31:0]}; // @[EXU_AXI.scala 58:37]
  wire [62:0] sllw_res = _GEN_2 << src2_value[4:0]; // @[EXU_AXI.scala 58:37]
  wire [63:0] or_res = src1_value | src2_value; // @[EXU_AXI.scala 59:29]
  wire [63:0] xor_res = src1_value ^ src2_value; // @[EXU_AXI.scala 60:30]
  wire [63:0] and_res = src1_value & src2_value; // @[EXU_AXI.scala 61:30]
  wire [127:0] _mlu_res_T = src1_value * src2_value; // @[EXU_AXI.scala 62:31]
  wire [63:0] mlu_res = _mlu_res_T[63:0]; // @[EXU_AXI.scala 62:44]
  wire [63:0] _mluw_res_T_2 = src1_value[31:0] * src2_value[31:0]; // @[EXU_AXI.scala 63:38]
  wire [31:0] mluw_res = _mluw_res_T_2[31:0]; // @[EXU_AXI.scala 63:57]
  wire [31:0] _divw_res_T_3 = src2_value[31:0]; // @[EXU_AXI.scala 64:64]
  wire [32:0] _divw_res_T_4 = $signed(_sraw_res_T_1) / $signed(_divw_res_T_3); // @[EXU_AXI.scala 64:45]
  wire [31:0] divw_res = _divw_res_T_4[31:0]; // @[EXU_AXI.scala 64:71]
  wire [31:0] divuw_res = src1_value[31:0] / src2_value[31:0]; // @[EXU_AXI.scala 65:39]
  wire [31:0] remw_res = $signed(_sraw_res_T_1) % $signed(_divw_res_T_3); // @[EXU_AXI.scala 66:71]
  wire [31:0] remuw_res = src1_value[31:0] % src2_value[31:0]; // @[EXU_AXI.scala 67:39]
  wire [63:0] _div_res_T_1 = io_ctrl_sign_src2_is_imm ? io_imm : _src2_value_T_1; // @[EXU_AXI.scala 68:51]
  wire [64:0] div_res = $signed(_sra_res_T) / $signed(_div_res_T_1); // @[EXU_AXI.scala 68:59]
  wire [63:0] divu_res = src1_value / src2_value; // @[EXU_AXI.scala 69:31]
  wire [63:0] rem_res = $signed(_sra_res_T) % $signed(_div_res_T_1); // @[EXU_AXI.scala 70:59]
  wire [63:0] remu_res = src1_value % src2_value; // @[EXU_AXI.scala 71:31]
  wire [63:0] _io_res2rd_T_1 = io_pc + 64'h4; // @[EXU_AXI.scala 76:24]
  wire  _io_res2rd_T_4 = src1_value < src2_value; // @[EXU_AXI.scala 78:34]
  wire  _io_res2rd_T_10 = $signed(_sra_res_T) < $signed(_div_res_T_1); // @[EXU_AXI.scala 80:42]
  wire [31:0] _io_res2rd_T_18 = io_Mem_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_20 = {_io_res2rd_T_18,io_Mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_23 = {56'h0,io_Mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_26 = {32'h0,io_Mem_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [47:0] _io_res2rd_T_29 = io_Mem_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_31 = {_io_res2rd_T_29,io_Mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [55:0] _io_res2rd_T_34 = io_Mem_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_36 = {_io_res2rd_T_34,io_Mem_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_39 = {48'h0,io_Mem_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_42 = add_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_44 = {_io_res2rd_T_42,add_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_52 = sub_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_54 = {_io_res2rd_T_52,sub_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_57 = sllw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_59 = {_io_res2rd_T_57,sllw_res[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_67 = sraw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _io_res2rd_T_68 = $signed(_sraw_res_T_1) >>> src2_value[4:0]; // @[EXU_AXI.scala 105:56]
  wire [63:0] _io_res2rd_T_69 = {_io_res2rd_T_67,_io_res2rd_T_68}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_72 = srlw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_74 = {_io_res2rd_T_72,srlw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_87 = mluw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_88 = {_io_res2rd_T_87,mluw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_91 = divw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_92 = {_io_res2rd_T_91,divw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_95 = divuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_96 = {_io_res2rd_T_95,divuw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_99 = remw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_100 = {_io_res2rd_T_99,remw_res}; // @[Cat.scala 31:58]
  wire [31:0] _io_res2rd_T_103 = remuw_res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_res2rd_T_104 = {_io_res2rd_T_103,remuw_res}; // @[Cat.scala 31:58]
  wire [63:0] _io_res2rd_T_106 = 32'h1 == io_inst_now ? add_res : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_108 = 32'h3 == io_inst_now ? add_res : _io_res2rd_T_106; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_110 = 32'h4 == io_inst_now ? io_imm : _io_res2rd_T_108; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_112 = 32'h5 == io_inst_now ? _io_res2rd_T_1 : _io_res2rd_T_110; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_114 = 32'h6 == io_inst_now ? _io_res2rd_T_1 : _io_res2rd_T_112; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_116 = 32'h20 == io_inst_now ? {{63'd0}, _io_res2rd_T_4} : _io_res2rd_T_114; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_118 = 32'h1e == io_inst_now ? {{63'd0}, _io_res2rd_T_4} : _io_res2rd_T_116; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_120 = 32'h36 == io_inst_now ? {{63'd0}, _io_res2rd_T_10} : _io_res2rd_T_118; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_122 = 32'h1f == io_inst_now ? {{63'd0}, _io_res2rd_T_10} : _io_res2rd_T_120; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_124 = 32'h21 == io_inst_now ? _io_res2rd_T_20 : _io_res2rd_T_122; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_126 = 32'h22 == io_inst_now ? io_Mem_rdata : _io_res2rd_T_124; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_128 = 32'h23 == io_inst_now ? _io_res2rd_T_23 : _io_res2rd_T_126; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_130 = 32'h3a == io_inst_now ? _io_res2rd_T_26 : _io_res2rd_T_128; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_132 = 32'h24 == io_inst_now ? _io_res2rd_T_31 : _io_res2rd_T_130; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_134 = 32'h3b == io_inst_now ? _io_res2rd_T_36 : _io_res2rd_T_132; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_136 = 32'h25 == io_inst_now ? _io_res2rd_T_39 : _io_res2rd_T_134; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_138 = 32'hc == io_inst_now ? _io_res2rd_T_44 : _io_res2rd_T_136; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_140 = 32'he == io_inst_now ? sub_res : _io_res2rd_T_138; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_142 = 32'h10 == io_inst_now ? _io_res2rd_T_44 : _io_res2rd_T_140; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_144 = 32'hf == io_inst_now ? add_res : _io_res2rd_T_142; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_146 = 32'h15 == io_inst_now ? sra_res : _io_res2rd_T_144; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_148 = 32'hb == io_inst_now ? or_res : _io_res2rd_T_146; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_150 = 32'h2f == io_inst_now ? or_res : _io_res2rd_T_148; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_152 = 32'h2e == io_inst_now ? xor_res : _io_res2rd_T_150; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_154 = 32'ha == io_inst_now ? xor_res : _io_res2rd_T_152; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_156 = 32'h8 == io_inst_now ? and_res : _io_res2rd_T_154; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_158 = 32'h9 == io_inst_now ? and_res : _io_res2rd_T_156; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_160 = 32'hd == io_inst_now ? _io_res2rd_T_54 : _io_res2rd_T_158; // @[Mux.scala 81:58]
  wire [63:0] _io_res2rd_T_162 = 32'h16 == io_inst_now ? _io_res2rd_T_59 : _io_res2rd_T_160; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_164 = 32'h17 == io_inst_now ? sll_res : {{63'd0}, _io_res2rd_T_162}; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_166 = 32'h18 == io_inst_now ? {{63'd0}, srl_res} : _io_res2rd_T_164; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_168 = 32'h19 == io_inst_now ? {{63'd0}, _io_res2rd_T_59} : _io_res2rd_T_166; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_170 = 32'h1a == io_inst_now ? {{63'd0}, _io_res2rd_T_69} : _io_res2rd_T_168; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_172 = 32'h1b == io_inst_now ? {{63'd0}, _io_res2rd_T_74} : _io_res2rd_T_170; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_174 = 32'h1c == io_inst_now ? {{63'd0}, _io_res2rd_T_69} : _io_res2rd_T_172; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_176 = 32'h1d == io_inst_now ? {{63'd0}, _io_res2rd_T_74} : _io_res2rd_T_174; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_178 = 32'h11 == io_inst_now ? {{63'd0}, mlu_res} : _io_res2rd_T_176; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_180 = 32'h12 == io_inst_now ? {{63'd0}, _io_res2rd_T_88} : _io_res2rd_T_178; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_182 = 32'h13 == io_inst_now ? {{63'd0}, _io_res2rd_T_92} : _io_res2rd_T_180; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_184 = 32'h30 == io_inst_now ? {{63'd0}, divu_res} : _io_res2rd_T_182; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_186 = 32'h31 == io_inst_now ? {{62'd0}, div_res} : _io_res2rd_T_184; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_188 = 32'h35 == io_inst_now ? {{63'd0}, _io_res2rd_T_96} : _io_res2rd_T_186; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_190 = 32'h14 == io_inst_now ? {{63'd0}, _io_res2rd_T_100} : _io_res2rd_T_188; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_192 = 32'h32 == io_inst_now ? {{63'd0}, _io_res2rd_T_104} : _io_res2rd_T_190; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_194 = 32'h33 == io_inst_now ? {{63'd0}, remu_res} : _io_res2rd_T_192; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_196 = 32'h34 == io_inst_now ? {{63'd0}, rem_res} : _io_res2rd_T_194; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_198 = 32'h37 == io_inst_now ? sll_res : _io_res2rd_T_196; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_200 = 32'h39 == io_inst_now ? {{63'd0}, sra_res} : _io_res2rd_T_198; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_202 = 32'h38 == io_inst_now ? {{63'd0}, srl_res} : _io_res2rd_T_200; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_204 = 32'h3f == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_data} : _io_res2rd_T_202; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_206 = 32'h46 == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_1_data} : _io_res2rd_T_204; // @[Mux.scala 81:58]
  wire [126:0] _io_res2rd_T_208 = 32'h47 == io_inst_now ? {{63'd0}, CSR_Reg_io_res2rd_MPORT_2_data} : _io_res2rd_T_206; // @[Mux.scala 81:58]
  wire [63:0] reg_value = io_rd == 5'h0 ? 64'h0 : Regfile_reg_value_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire  _T_6 = io_ctrl_sign_reg_write & io_rd != 5'h0 & (io_inst_valid & ~io_ctrl_sign_Readmem_en |
    io_ctrl_sign_Readmem_en & io_rdata_valid); // @[EXU_AXI.scala 129:63]
  wire [63:0] _csr_wdata_T = src1_value | CSR_Reg_csr_wdata_MPORT_data; // @[EXU_AXI.scala 134:32]
  wire [63:0] _csr_wdata_T_1 = ~CSR_Reg_csr_wdata_MPORT_1_data; // @[EXU_AXI.scala 135:35]
  wire [63:0] _csr_wdata_T_2 = src1_value & _csr_wdata_T_1; // @[EXU_AXI.scala 135:32]
  wire [63:0] _csr_wdata_T_4 = 32'h3f == io_inst_now ? src1_value : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _csr_wdata_T_6 = 32'h46 == io_inst_now ? _csr_wdata_T : _csr_wdata_T_4; // @[Mux.scala 81:58]
  wire [63:0] csr_wdata = 32'h47 == io_inst_now ? _csr_wdata_T_2 : _csr_wdata_T_6; // @[Mux.scala 81:58]
  wire  _T_9 = io_inst_now == 32'h3d & io_inst_valid; // @[EXU_AXI.scala 138:48]
  wire  _T_14 = io_ctrl_sign_csr_write & io_inst_valid; // @[EXU_AXI.scala 141:53]
  wire [63:0] _j_pc_T = add_res & 64'hfffffffffffffffe; // @[EXU_AXI.scala 148:28]
  wire [63:0] _j_pc_T_3 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_data; // @[EXU_AXI.scala 149:39]
  wire [63:0] _j_pc_T_6 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_1_data; // @[EXU_AXI.scala 149:67]
  wire [63:0] _j_pc_T_8 = $signed(_j_pc_T_3) != $signed(_j_pc_T_6) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 149:21]
  wire [63:0] _j_pc_T_11 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_2_data; // @[EXU_AXI.scala 150:39]
  wire [63:0] _j_pc_T_14 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_3_data; // @[EXU_AXI.scala 150:67]
  wire [63:0] _j_pc_T_16 = $signed(_j_pc_T_11) == $signed(_j_pc_T_14) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 150:21]
  wire [63:0] _j_pc_T_19 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_4_data; // @[EXU_AXI.scala 151:39]
  wire [63:0] _j_pc_T_22 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_5_data; // @[EXU_AXI.scala 151:66]
  wire [63:0] _j_pc_T_24 = $signed(_j_pc_T_19) >= $signed(_j_pc_T_22) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 151:21]
  wire [63:0] _j_pc_T_27 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_6_data; // @[EXU_AXI.scala 152:39]
  wire [63:0] _j_pc_T_30 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_7_data; // @[EXU_AXI.scala 152:65]
  wire [63:0] _j_pc_T_32 = $signed(_j_pc_T_27) < $signed(_j_pc_T_30) ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 152:21]
  wire [63:0] _j_pc_T_34 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_8_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_36 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_9_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_38 = _j_pc_T_34 < _j_pc_T_36 ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 153:22]
  wire [63:0] _j_pc_T_40 = io_rs1 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_10_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_42 = io_rs2 == 5'h0 ? 64'h0 : Regfile_j_pc_MPORT_11_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _j_pc_T_44 = _j_pc_T_40 >= _j_pc_T_42 ? add_res : _io_res2rd_T_1; // @[EXU_AXI.scala 154:22]
  wire [63:0] _j_pc_T_46 = CSR_Reg_j_pc_MPORT_13_data + 64'h4; // @[EXU_AXI.scala 156:33]
  wire [63:0] _j_pc_T_48 = 32'h5 == io_inst_now ? add_res : _io_res2rd_T_1; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_50 = 32'h6 == io_inst_now ? _j_pc_T : _j_pc_T_48; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_52 = 32'h2a == io_inst_now ? _j_pc_T_8 : _j_pc_T_50; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_54 = 32'h29 == io_inst_now ? _j_pc_T_16 : _j_pc_T_52; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_56 = 32'h2b == io_inst_now ? _j_pc_T_24 : _j_pc_T_54; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_58 = 32'h2c == io_inst_now ? _j_pc_T_32 : _j_pc_T_56; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_60 = 32'h2d == io_inst_now ? _j_pc_T_38 : _j_pc_T_58; // @[Mux.scala 81:58]
  wire [63:0] _j_pc_T_62 = 32'h3c == io_inst_now ? _j_pc_T_44 : _j_pc_T_60; // @[Mux.scala 81:58]
  reg [63:0] pc_next; // @[EXU_AXI.scala 158:26]
  wire [63:0] _mem_wdata_T_1 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_3 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_1_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_6 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_2_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_9 = io_rs2 == 5'h0 ? 64'h0 : Regfile_mem_wdata_MPORT_3_data; // @[EXU_AXI.scala 47:12]
  wire [63:0] _mem_wdata_T_12 = 32'h7 == io_inst_now ? _mem_wdata_T_1 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _mem_wdata_T_14 = 32'h26 == io_inst_now ? {{48'd0}, _mem_wdata_T_3[15:0]} : _mem_wdata_T_12; // @[Mux.scala 81:58]
  wire [63:0] _mem_wdata_T_16 = 32'h28 == io_inst_now ? {{56'd0}, _mem_wdata_T_6[7:0]} : _mem_wdata_T_14; // @[Mux.scala 81:58]
  traceregs reg_trace ( // @[EXU_AXI.scala 163:27]
    .input_reg_0(reg_trace_input_reg_0),
    .input_reg_1(reg_trace_input_reg_1),
    .input_reg_2(reg_trace_input_reg_2),
    .input_reg_3(reg_trace_input_reg_3),
    .input_reg_4(reg_trace_input_reg_4),
    .input_reg_5(reg_trace_input_reg_5),
    .input_reg_6(reg_trace_input_reg_6),
    .input_reg_7(reg_trace_input_reg_7),
    .input_reg_8(reg_trace_input_reg_8),
    .input_reg_9(reg_trace_input_reg_9),
    .input_reg_10(reg_trace_input_reg_10),
    .input_reg_11(reg_trace_input_reg_11),
    .input_reg_12(reg_trace_input_reg_12),
    .input_reg_13(reg_trace_input_reg_13),
    .input_reg_14(reg_trace_input_reg_14),
    .input_reg_15(reg_trace_input_reg_15),
    .input_reg_16(reg_trace_input_reg_16),
    .input_reg_17(reg_trace_input_reg_17),
    .input_reg_18(reg_trace_input_reg_18),
    .input_reg_19(reg_trace_input_reg_19),
    .input_reg_20(reg_trace_input_reg_20),
    .input_reg_21(reg_trace_input_reg_21),
    .input_reg_22(reg_trace_input_reg_22),
    .input_reg_23(reg_trace_input_reg_23),
    .input_reg_24(reg_trace_input_reg_24),
    .input_reg_25(reg_trace_input_reg_25),
    .input_reg_26(reg_trace_input_reg_26),
    .input_reg_27(reg_trace_input_reg_27),
    .input_reg_28(reg_trace_input_reg_28),
    .input_reg_29(reg_trace_input_reg_29),
    .input_reg_30(reg_trace_input_reg_30),
    .input_reg_31(reg_trace_input_reg_31),
    .csr_reg_0(reg_trace_csr_reg_0),
    .csr_reg_1(reg_trace_csr_reg_1),
    .csr_reg_2(reg_trace_csr_reg_2),
    .csr_reg_3(reg_trace_csr_reg_3),
    .pc(reg_trace_pc)
  );
  assign Regfile_src1_value_MPORT_en = 1'h1;
  assign Regfile_src1_value_MPORT_addr = io_rs1;
  assign Regfile_src1_value_MPORT_data = Regfile[Regfile_src1_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_src2_value_MPORT_en = 1'h1;
  assign Regfile_src2_value_MPORT_addr = io_rs2;
  assign Regfile_src2_value_MPORT_data = Regfile[Regfile_src2_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_value_MPORT_en = 1'h1;
  assign Regfile_reg_value_MPORT_addr = io_rd;
  assign Regfile_reg_value_MPORT_data = Regfile[Regfile_reg_value_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_MPORT_4_en = 1'h1;
  assign Regfile_MPORT_4_addr = 5'h11;
  assign Regfile_MPORT_4_data = Regfile[Regfile_MPORT_4_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_en = 1'h1;
  assign Regfile_j_pc_MPORT_addr = io_rs1;
  assign Regfile_j_pc_MPORT_data = Regfile[Regfile_j_pc_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_1_en = 1'h1;
  assign Regfile_j_pc_MPORT_1_addr = io_rs2;
  assign Regfile_j_pc_MPORT_1_data = Regfile[Regfile_j_pc_MPORT_1_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_2_en = 1'h1;
  assign Regfile_j_pc_MPORT_2_addr = io_rs1;
  assign Regfile_j_pc_MPORT_2_data = Regfile[Regfile_j_pc_MPORT_2_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_3_en = 1'h1;
  assign Regfile_j_pc_MPORT_3_addr = io_rs2;
  assign Regfile_j_pc_MPORT_3_data = Regfile[Regfile_j_pc_MPORT_3_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_4_en = 1'h1;
  assign Regfile_j_pc_MPORT_4_addr = io_rs1;
  assign Regfile_j_pc_MPORT_4_data = Regfile[Regfile_j_pc_MPORT_4_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_5_en = 1'h1;
  assign Regfile_j_pc_MPORT_5_addr = io_rs2;
  assign Regfile_j_pc_MPORT_5_data = Regfile[Regfile_j_pc_MPORT_5_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_6_en = 1'h1;
  assign Regfile_j_pc_MPORT_6_addr = io_rs1;
  assign Regfile_j_pc_MPORT_6_data = Regfile[Regfile_j_pc_MPORT_6_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_7_en = 1'h1;
  assign Regfile_j_pc_MPORT_7_addr = io_rs2;
  assign Regfile_j_pc_MPORT_7_data = Regfile[Regfile_j_pc_MPORT_7_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_8_en = 1'h1;
  assign Regfile_j_pc_MPORT_8_addr = io_rs1;
  assign Regfile_j_pc_MPORT_8_data = Regfile[Regfile_j_pc_MPORT_8_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_9_en = 1'h1;
  assign Regfile_j_pc_MPORT_9_addr = io_rs2;
  assign Regfile_j_pc_MPORT_9_data = Regfile[Regfile_j_pc_MPORT_9_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_10_en = 1'h1;
  assign Regfile_j_pc_MPORT_10_addr = io_rs1;
  assign Regfile_j_pc_MPORT_10_data = Regfile[Regfile_j_pc_MPORT_10_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_j_pc_MPORT_11_en = 1'h1;
  assign Regfile_j_pc_MPORT_11_addr = io_rs2;
  assign Regfile_j_pc_MPORT_11_data = Regfile[Regfile_j_pc_MPORT_11_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_0_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_0_MPORT_addr = 5'h0;
  assign Regfile_reg_trace_io_input_reg_0_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_0_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_1_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_1_MPORT_addr = 5'h1;
  assign Regfile_reg_trace_io_input_reg_1_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_1_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_2_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_2_MPORT_addr = 5'h2;
  assign Regfile_reg_trace_io_input_reg_2_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_2_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_3_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_3_MPORT_addr = 5'h3;
  assign Regfile_reg_trace_io_input_reg_3_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_3_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_4_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_4_MPORT_addr = 5'h4;
  assign Regfile_reg_trace_io_input_reg_4_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_4_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_5_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_5_MPORT_addr = 5'h5;
  assign Regfile_reg_trace_io_input_reg_5_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_5_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_6_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_6_MPORT_addr = 5'h6;
  assign Regfile_reg_trace_io_input_reg_6_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_6_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_7_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_7_MPORT_addr = 5'h7;
  assign Regfile_reg_trace_io_input_reg_7_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_7_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_8_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_8_MPORT_addr = 5'h8;
  assign Regfile_reg_trace_io_input_reg_8_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_8_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_9_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_9_MPORT_addr = 5'h9;
  assign Regfile_reg_trace_io_input_reg_9_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_9_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_10_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_10_MPORT_addr = 5'ha;
  assign Regfile_reg_trace_io_input_reg_10_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_10_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_11_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_11_MPORT_addr = 5'hb;
  assign Regfile_reg_trace_io_input_reg_11_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_11_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_12_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_12_MPORT_addr = 5'hc;
  assign Regfile_reg_trace_io_input_reg_12_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_12_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_13_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_13_MPORT_addr = 5'hd;
  assign Regfile_reg_trace_io_input_reg_13_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_13_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_14_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_14_MPORT_addr = 5'he;
  assign Regfile_reg_trace_io_input_reg_14_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_14_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_15_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_15_MPORT_addr = 5'hf;
  assign Regfile_reg_trace_io_input_reg_15_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_15_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_16_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_16_MPORT_addr = 5'h10;
  assign Regfile_reg_trace_io_input_reg_16_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_16_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_17_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_17_MPORT_addr = 5'h11;
  assign Regfile_reg_trace_io_input_reg_17_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_17_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_18_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_18_MPORT_addr = 5'h12;
  assign Regfile_reg_trace_io_input_reg_18_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_18_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_19_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_19_MPORT_addr = 5'h13;
  assign Regfile_reg_trace_io_input_reg_19_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_19_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_20_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_20_MPORT_addr = 5'h14;
  assign Regfile_reg_trace_io_input_reg_20_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_20_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_21_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_21_MPORT_addr = 5'h15;
  assign Regfile_reg_trace_io_input_reg_21_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_21_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_22_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_22_MPORT_addr = 5'h16;
  assign Regfile_reg_trace_io_input_reg_22_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_22_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_23_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_23_MPORT_addr = 5'h17;
  assign Regfile_reg_trace_io_input_reg_23_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_23_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_24_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_24_MPORT_addr = 5'h18;
  assign Regfile_reg_trace_io_input_reg_24_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_24_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_25_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_25_MPORT_addr = 5'h19;
  assign Regfile_reg_trace_io_input_reg_25_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_25_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_26_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_26_MPORT_addr = 5'h1a;
  assign Regfile_reg_trace_io_input_reg_26_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_26_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_27_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_27_MPORT_addr = 5'h1b;
  assign Regfile_reg_trace_io_input_reg_27_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_27_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_28_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_28_MPORT_addr = 5'h1c;
  assign Regfile_reg_trace_io_input_reg_28_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_28_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_29_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_29_MPORT_addr = 5'h1d;
  assign Regfile_reg_trace_io_input_reg_29_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_29_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_30_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_30_MPORT_addr = 5'h1e;
  assign Regfile_reg_trace_io_input_reg_30_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_30_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_reg_trace_io_input_reg_31_MPORT_en = 1'h1;
  assign Regfile_reg_trace_io_input_reg_31_MPORT_addr = 5'h1f;
  assign Regfile_reg_trace_io_input_reg_31_MPORT_data = Regfile[Regfile_reg_trace_io_input_reg_31_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_data = Regfile[Regfile_mem_wdata_MPORT_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_1_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_1_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_1_data = Regfile[Regfile_mem_wdata_MPORT_1_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_2_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_2_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_2_data = Regfile[Regfile_mem_wdata_MPORT_2_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_mem_wdata_MPORT_3_en = 1'h1;
  assign Regfile_mem_wdata_MPORT_3_addr = io_rs2;
  assign Regfile_mem_wdata_MPORT_3_data = Regfile[Regfile_mem_wdata_MPORT_3_addr]; // @[EXU_AXI.scala 37:22]
  assign Regfile_MPORT_data = _T_6 ? io_res2rd : reg_value;
  assign Regfile_MPORT_addr = io_rd;
  assign Regfile_MPORT_mask = 1'h1;
  assign Regfile_MPORT_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_io_res2rd_MPORT_1_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_1_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_1_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_1_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_io_res2rd_MPORT_2_en = 1'h1;
  assign CSR_Reg_io_res2rd_MPORT_2_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_io_res2rd_MPORT_2_data = CSR_Reg[CSR_Reg_io_res2rd_MPORT_2_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_csr_wdata_MPORT_en = 1'h1;
  assign CSR_Reg_csr_wdata_MPORT_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_csr_wdata_MPORT_data = CSR_Reg[CSR_Reg_csr_wdata_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_csr_wdata_MPORT_1_en = 1'h1;
  assign CSR_Reg_csr_wdata_MPORT_1_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_csr_wdata_MPORT_1_data = CSR_Reg[CSR_Reg_csr_wdata_MPORT_1_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_2_en = 1'h1;
  assign CSR_Reg_MPORT_2_addr = 2'h1;
  assign CSR_Reg_MPORT_2_data = CSR_Reg[CSR_Reg_MPORT_2_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_5_en = 1'h1;
  assign CSR_Reg_MPORT_5_addr = 2'h3;
  assign CSR_Reg_MPORT_5_data = CSR_Reg[CSR_Reg_MPORT_5_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_7_en = 1'h1;
  assign CSR_Reg_MPORT_7_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_MPORT_7_data = CSR_Reg[CSR_Reg_MPORT_7_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_j_pc_MPORT_12_en = 1'h1;
  assign CSR_Reg_j_pc_MPORT_12_addr = 2'h0;
  assign CSR_Reg_j_pc_MPORT_12_data = CSR_Reg[CSR_Reg_j_pc_MPORT_12_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_j_pc_MPORT_13_en = 1'h1;
  assign CSR_Reg_j_pc_MPORT_13_addr = 2'h1;
  assign CSR_Reg_j_pc_MPORT_13_data = CSR_Reg[CSR_Reg_j_pc_MPORT_13_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr = 2'h0;
  assign CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_0_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr = 2'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_1_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_en = 1'h1;
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr = 2'h2;
  assign CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data = CSR_Reg[CSR_Reg_reg_trace_io_csr_reg_2_MPORT_addr]; // @[EXU_AXI.scala 38:22]
  assign CSR_Reg_MPORT_1_data = _T_9 ? io_pc : CSR_Reg_MPORT_2_data;
  assign CSR_Reg_MPORT_1_addr = 2'h1;
  assign CSR_Reg_MPORT_1_mask = 1'h1;
  assign CSR_Reg_MPORT_1_en = 1'h1;
  assign CSR_Reg_MPORT_3_data = _T_9 ? Regfile_MPORT_4_data : CSR_Reg_MPORT_5_data;
  assign CSR_Reg_MPORT_3_addr = 2'h3;
  assign CSR_Reg_MPORT_3_mask = 1'h1;
  assign CSR_Reg_MPORT_3_en = 1'h1;
  assign CSR_Reg_MPORT_6_data = _T_14 ? csr_wdata : CSR_Reg_MPORT_7_data;
  assign CSR_Reg_MPORT_6_addr = _csr_index_T_6 ? 2'h3 : _csr_index_T_5;
  assign CSR_Reg_MPORT_6_mask = 1'h1;
  assign CSR_Reg_MPORT_6_en = 1'h1;
  assign io_pc_next = pc_next; // @[EXU_AXI.scala 162:16]
  assign io_res2rd = _io_res2rd_T_208[63:0]; // @[EXU_AXI.scala 72:15]
  assign io_inst_store = io_ctrl_sign_Writemem_en; // @[EXU_AXI.scala 188:19]
  assign io_inst_load = io_ctrl_sign_Readmem_en; // @[EXU_AXI.scala 189:18]
  assign io_Mem_addr = add_res[31:0]; // @[EXU_AXI.scala 190:17]
  assign io_Mem_wdata = 32'h27 == io_inst_now ? {{32'd0}, _mem_wdata_T_9[31:0]} : _mem_wdata_T_16; // @[Mux.scala 81:58]
  assign io_Mem_wstrb = io_ctrl_sign_Wmask; // @[EXU_AXI.scala 192:18]
  assign reg_trace_input_reg_0 = Regfile_reg_trace_io_input_reg_0_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_1 = Regfile_reg_trace_io_input_reg_1_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_2 = Regfile_reg_trace_io_input_reg_2_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_3 = Regfile_reg_trace_io_input_reg_3_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_4 = Regfile_reg_trace_io_input_reg_4_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_5 = Regfile_reg_trace_io_input_reg_5_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_6 = Regfile_reg_trace_io_input_reg_6_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_7 = Regfile_reg_trace_io_input_reg_7_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_8 = Regfile_reg_trace_io_input_reg_8_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_9 = Regfile_reg_trace_io_input_reg_9_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_10 = Regfile_reg_trace_io_input_reg_10_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_11 = Regfile_reg_trace_io_input_reg_11_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_12 = Regfile_reg_trace_io_input_reg_12_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_13 = Regfile_reg_trace_io_input_reg_13_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_14 = Regfile_reg_trace_io_input_reg_14_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_15 = Regfile_reg_trace_io_input_reg_15_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_16 = Regfile_reg_trace_io_input_reg_16_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_17 = Regfile_reg_trace_io_input_reg_17_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_18 = Regfile_reg_trace_io_input_reg_18_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_19 = Regfile_reg_trace_io_input_reg_19_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_20 = Regfile_reg_trace_io_input_reg_20_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_21 = Regfile_reg_trace_io_input_reg_21_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_22 = Regfile_reg_trace_io_input_reg_22_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_23 = Regfile_reg_trace_io_input_reg_23_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_24 = Regfile_reg_trace_io_input_reg_24_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_25 = Regfile_reg_trace_io_input_reg_25_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_26 = Regfile_reg_trace_io_input_reg_26_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_27 = Regfile_reg_trace_io_input_reg_27_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_28 = Regfile_reg_trace_io_input_reg_28_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_29 = Regfile_reg_trace_io_input_reg_29_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_30 = Regfile_reg_trace_io_input_reg_30_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_input_reg_31 = Regfile_reg_trace_io_input_reg_31_MPORT_data; // @[EXU_AXI.scala 165:57]
  assign reg_trace_csr_reg_0 = CSR_Reg_reg_trace_io_csr_reg_0_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_1 = CSR_Reg_reg_trace_io_csr_reg_1_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_2 = CSR_Reg_reg_trace_io_csr_reg_2_MPORT_data; // @[EXU_AXI.scala 168:54]
  assign reg_trace_csr_reg_3 = 64'h0; // @[EXU_AXI.scala 167:{36,36}]
  assign reg_trace_pc = io_pc; // @[EXU_AXI.scala 166:21]
  always @(posedge clock) begin
    if (Regfile_MPORT_en & Regfile_MPORT_mask) begin
      Regfile[Regfile_MPORT_addr] <= Regfile_MPORT_data; // @[EXU_AXI.scala 37:22]
    end
    if (CSR_Reg_MPORT_1_en & CSR_Reg_MPORT_1_mask) begin
      CSR_Reg[CSR_Reg_MPORT_1_addr] <= CSR_Reg_MPORT_1_data; // @[EXU_AXI.scala 38:22]
    end
    if (CSR_Reg_MPORT_3_en & CSR_Reg_MPORT_3_mask) begin
      CSR_Reg[CSR_Reg_MPORT_3_addr] <= CSR_Reg_MPORT_3_data; // @[EXU_AXI.scala 38:22]
    end
    if (CSR_Reg_MPORT_6_en & CSR_Reg_MPORT_6_mask) begin
      CSR_Reg[CSR_Reg_MPORT_6_addr] <= CSR_Reg_MPORT_6_data; // @[EXU_AXI.scala 38:22]
    end
    if (reset) begin // @[EXU_AXI.scala 158:26]
      pc_next <= 64'h0; // @[EXU_AXI.scala 158:26]
    end else if (io_inst_valid) begin // @[EXU_AXI.scala 159:24]
      if (32'h3e == io_inst_now) begin // @[Mux.scala 81:58]
        pc_next <= _j_pc_T_46;
      end else if (32'h3d == io_inst_now) begin // @[Mux.scala 81:58]
        pc_next <= CSR_Reg_j_pc_MPORT_12_data;
      end else begin
        pc_next <= _j_pc_T_62;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    Regfile[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    CSR_Reg[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  pc_next = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input         clock,
  input         reset,
  output [31:0] io_inst,
  output [63:0] io_pc,
  output [63:0] io_pc_next,
  output [63:0] io_outval,
  output        io_step
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  axi_clock; // @[top.scala 18:21]
  wire  axi_reset; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_araddr; // @[top.scala 18:21]
  wire  axi_io_axi_in_arvalid; // @[top.scala 18:21]
  wire  axi_io_axi_in_rready; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_awaddr; // @[top.scala 18:21]
  wire  axi_io_axi_in_awvalid; // @[top.scala 18:21]
  wire [31:0] axi_io_axi_in_wdata; // @[top.scala 18:21]
  wire [7:0] axi_io_axi_in_wstrb; // @[top.scala 18:21]
  wire  axi_io_axi_in_wvalid; // @[top.scala 18:21]
  wire  axi_io_axi_in_bready; // @[top.scala 18:21]
  wire  axi_io_axi_out_arready; // @[top.scala 18:21]
  wire [63:0] axi_io_axi_out_rdata; // @[top.scala 18:21]
  wire  axi_io_axi_out_rvalid; // @[top.scala 18:21]
  wire  axi_io_axi_out_awready; // @[top.scala 18:21]
  wire  axi_io_axi_out_wready; // @[top.scala 18:21]
  wire  axi_io_axi_out_bvalid; // @[top.scala 18:21]
  wire  lsu_step_clock; // @[top.scala 19:26]
  wire  lsu_step_reset; // @[top.scala 19:26]
  wire  lsu_step_io_inst_store; // @[top.scala 19:26]
  wire  lsu_step_io_inst_load; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_mem_addr; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_mem_wdata; // @[top.scala 19:26]
  wire [7:0] lsu_step_io_mem_wstrb; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_mem_rdata; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_arready; // @[top.scala 19:26]
  wire [63:0] lsu_step_io_axi_in_rdata; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_rvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_awready; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_wready; // @[top.scala 19:26]
  wire  lsu_step_io_axi_in_bvalid; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_araddr; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_arvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_rready; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_awaddr; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_awvalid; // @[top.scala 19:26]
  wire [31:0] lsu_step_io_axi_out_wdata; // @[top.scala 19:26]
  wire [7:0] lsu_step_io_axi_out_wstrb; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_wvalid; // @[top.scala 19:26]
  wire  lsu_step_io_axi_out_bready; // @[top.scala 19:26]
  wire  arbiter_clock; // @[top.scala 20:25]
  wire  arbiter_reset; // @[top.scala 20:25]
  wire [31:0] arbiter_io_ifu_axi_in_araddr; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_in_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_in_rready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_ifu_axi_out_rdata; // @[top.scala 20:25]
  wire  arbiter_io_ifu_axi_out_rvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_araddr; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_rready; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_awaddr; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_awvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_lsu_axi_in_wdata; // @[top.scala 20:25]
  wire [7:0] arbiter_io_lsu_axi_in_wstrb; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_wvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_in_bready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_arready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_lsu_axi_out_rdata; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_rvalid; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_awready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_wready; // @[top.scala 20:25]
  wire  arbiter_io_lsu_axi_out_bvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_arready; // @[top.scala 20:25]
  wire [63:0] arbiter_io_axi_in_rdata; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_rvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_awready; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_wready; // @[top.scala 20:25]
  wire  arbiter_io_axi_in_bvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_araddr; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_arvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_rready; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_awaddr; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_awvalid; // @[top.scala 20:25]
  wire [31:0] arbiter_io_axi_out_wdata; // @[top.scala 20:25]
  wire [7:0] arbiter_io_axi_out_wstrb; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_wvalid; // @[top.scala 20:25]
  wire  arbiter_io_axi_out_bready; // @[top.scala 20:25]
  wire  ifu_step_clock; // @[top.scala 21:26]
  wire  ifu_step_reset; // @[top.scala 21:26]
  wire [63:0] ifu_step_io_pc; // @[top.scala 21:26]
  wire  ifu_step_io_pc_valid; // @[top.scala 21:26]
  wire  ifu_step_io_inst_valid; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_inst; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_inst_reg; // @[top.scala 21:26]
  wire [63:0] ifu_step_io_axi_in_rdata; // @[top.scala 21:26]
  wire  ifu_step_io_axi_in_rvalid; // @[top.scala 21:26]
  wire [31:0] ifu_step_io_axi_out_araddr; // @[top.scala 21:26]
  wire  ifu_step_io_axi_out_arvalid; // @[top.scala 21:26]
  wire  ifu_step_io_axi_out_rready; // @[top.scala 21:26]
  wire  cache_clock; // @[top.scala 22:23]
  wire  cache_reset; // @[top.scala 22:23]
  wire [31:0] cache_io_from_ifu_araddr; // @[top.scala 22:23]
  wire  cache_io_from_ifu_arvalid; // @[top.scala 22:23]
  wire  cache_io_from_ifu_rready; // @[top.scala 22:23]
  wire [63:0] cache_io_to_ifu_rdata; // @[top.scala 22:23]
  wire  cache_io_to_ifu_rvalid; // @[top.scala 22:23]
  wire [31:0] cache_io_to_axi_araddr; // @[top.scala 22:23]
  wire  cache_io_to_axi_arvalid; // @[top.scala 22:23]
  wire  cache_io_to_axi_rready; // @[top.scala 22:23]
  wire [63:0] cache_io_from_axi_rdata; // @[top.scala 22:23]
  wire  cache_io_from_axi_rvalid; // @[top.scala 22:23]
  wire [31:0] idu_step_io_inst; // @[top.scala 39:26]
  wire [31:0] idu_step_io_inst_now; // @[top.scala 39:26]
  wire [4:0] idu_step_io_rs1; // @[top.scala 39:26]
  wire [4:0] idu_step_io_rs2; // @[top.scala 39:26]
  wire [4:0] idu_step_io_rd; // @[top.scala 39:26]
  wire [63:0] idu_step_io_imm; // @[top.scala 39:26]
  wire  idu_step_io_ctrl_sign_reg_write; // @[top.scala 39:26]
  wire  idu_step_io_ctrl_sign_csr_write; // @[top.scala 39:26]
  wire  idu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 39:26]
  wire  idu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 39:26]
  wire  idu_step_io_ctrl_sign_Writemem_en; // @[top.scala 39:26]
  wire  idu_step_io_ctrl_sign_Readmem_en; // @[top.scala 39:26]
  wire [7:0] idu_step_io_ctrl_sign_Wmask; // @[top.scala 39:26]
  wire  exu_step_clock; // @[top.scala 44:26]
  wire  exu_step_reset; // @[top.scala 44:26]
  wire [63:0] exu_step_io_pc; // @[top.scala 44:26]
  wire [63:0] exu_step_io_pc_next; // @[top.scala 44:26]
  wire [31:0] exu_step_io_inst_now; // @[top.scala 44:26]
  wire [4:0] exu_step_io_rs1; // @[top.scala 44:26]
  wire [4:0] exu_step_io_rs2; // @[top.scala 44:26]
  wire [4:0] exu_step_io_rd; // @[top.scala 44:26]
  wire [63:0] exu_step_io_imm; // @[top.scala 44:26]
  wire  exu_step_io_ctrl_sign_reg_write; // @[top.scala 44:26]
  wire  exu_step_io_ctrl_sign_csr_write; // @[top.scala 44:26]
  wire  exu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 44:26]
  wire  exu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 44:26]
  wire  exu_step_io_ctrl_sign_Writemem_en; // @[top.scala 44:26]
  wire  exu_step_io_ctrl_sign_Readmem_en; // @[top.scala 44:26]
  wire [7:0] exu_step_io_ctrl_sign_Wmask; // @[top.scala 44:26]
  wire [63:0] exu_step_io_res2rd; // @[top.scala 44:26]
  wire  exu_step_io_inst_valid; // @[top.scala 44:26]
  wire  exu_step_io_inst_store; // @[top.scala 44:26]
  wire  exu_step_io_inst_load; // @[top.scala 44:26]
  wire [31:0] exu_step_io_Mem_addr; // @[top.scala 44:26]
  wire [63:0] exu_step_io_Mem_rdata; // @[top.scala 44:26]
  wire [63:0] exu_step_io_Mem_wdata; // @[top.scala 44:26]
  wire [7:0] exu_step_io_Mem_wstrb; // @[top.scala 44:26]
  wire  exu_step_io_rdata_valid; // @[top.scala 44:26]
  wire [31:0] dpi_flag; // @[top.scala 66:21]
  wire [31:0] dpi_ecall_flag; // @[top.scala 66:21]
  reg [63:0] pc_now; // @[top.scala 15:25]
  reg  execute_end; // @[top.scala 17:30]
  reg  pc_valid; // @[top.scala 80:27]
  reg  diff_step; // @[top.scala 83:28]
  AXI axi ( // @[top.scala 18:21]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_axi_in_araddr(axi_io_axi_in_araddr),
    .io_axi_in_arvalid(axi_io_axi_in_arvalid),
    .io_axi_in_rready(axi_io_axi_in_rready),
    .io_axi_in_awaddr(axi_io_axi_in_awaddr),
    .io_axi_in_awvalid(axi_io_axi_in_awvalid),
    .io_axi_in_wdata(axi_io_axi_in_wdata),
    .io_axi_in_wstrb(axi_io_axi_in_wstrb),
    .io_axi_in_wvalid(axi_io_axi_in_wvalid),
    .io_axi_in_bready(axi_io_axi_in_bready),
    .io_axi_out_arready(axi_io_axi_out_arready),
    .io_axi_out_rdata(axi_io_axi_out_rdata),
    .io_axi_out_rvalid(axi_io_axi_out_rvalid),
    .io_axi_out_awready(axi_io_axi_out_awready),
    .io_axi_out_wready(axi_io_axi_out_wready),
    .io_axi_out_bvalid(axi_io_axi_out_bvalid)
  );
  LSU lsu_step ( // @[top.scala 19:26]
    .clock(lsu_step_clock),
    .reset(lsu_step_reset),
    .io_inst_store(lsu_step_io_inst_store),
    .io_inst_load(lsu_step_io_inst_load),
    .io_mem_addr(lsu_step_io_mem_addr),
    .io_mem_wdata(lsu_step_io_mem_wdata),
    .io_mem_wstrb(lsu_step_io_mem_wstrb),
    .io_mem_rdata(lsu_step_io_mem_rdata),
    .io_axi_in_arready(lsu_step_io_axi_in_arready),
    .io_axi_in_rdata(lsu_step_io_axi_in_rdata),
    .io_axi_in_rvalid(lsu_step_io_axi_in_rvalid),
    .io_axi_in_awready(lsu_step_io_axi_in_awready),
    .io_axi_in_wready(lsu_step_io_axi_in_wready),
    .io_axi_in_bvalid(lsu_step_io_axi_in_bvalid),
    .io_axi_out_araddr(lsu_step_io_axi_out_araddr),
    .io_axi_out_arvalid(lsu_step_io_axi_out_arvalid),
    .io_axi_out_rready(lsu_step_io_axi_out_rready),
    .io_axi_out_awaddr(lsu_step_io_axi_out_awaddr),
    .io_axi_out_awvalid(lsu_step_io_axi_out_awvalid),
    .io_axi_out_wdata(lsu_step_io_axi_out_wdata),
    .io_axi_out_wstrb(lsu_step_io_axi_out_wstrb),
    .io_axi_out_wvalid(lsu_step_io_axi_out_wvalid),
    .io_axi_out_bready(lsu_step_io_axi_out_bready)
  );
  AXI_ARBITER arbiter ( // @[top.scala 20:25]
    .clock(arbiter_clock),
    .reset(arbiter_reset),
    .io_ifu_axi_in_araddr(arbiter_io_ifu_axi_in_araddr),
    .io_ifu_axi_in_arvalid(arbiter_io_ifu_axi_in_arvalid),
    .io_ifu_axi_in_rready(arbiter_io_ifu_axi_in_rready),
    .io_ifu_axi_out_rdata(arbiter_io_ifu_axi_out_rdata),
    .io_ifu_axi_out_rvalid(arbiter_io_ifu_axi_out_rvalid),
    .io_lsu_axi_in_araddr(arbiter_io_lsu_axi_in_araddr),
    .io_lsu_axi_in_arvalid(arbiter_io_lsu_axi_in_arvalid),
    .io_lsu_axi_in_rready(arbiter_io_lsu_axi_in_rready),
    .io_lsu_axi_in_awaddr(arbiter_io_lsu_axi_in_awaddr),
    .io_lsu_axi_in_awvalid(arbiter_io_lsu_axi_in_awvalid),
    .io_lsu_axi_in_wdata(arbiter_io_lsu_axi_in_wdata),
    .io_lsu_axi_in_wstrb(arbiter_io_lsu_axi_in_wstrb),
    .io_lsu_axi_in_wvalid(arbiter_io_lsu_axi_in_wvalid),
    .io_lsu_axi_in_bready(arbiter_io_lsu_axi_in_bready),
    .io_lsu_axi_out_arready(arbiter_io_lsu_axi_out_arready),
    .io_lsu_axi_out_rdata(arbiter_io_lsu_axi_out_rdata),
    .io_lsu_axi_out_rvalid(arbiter_io_lsu_axi_out_rvalid),
    .io_lsu_axi_out_awready(arbiter_io_lsu_axi_out_awready),
    .io_lsu_axi_out_wready(arbiter_io_lsu_axi_out_wready),
    .io_lsu_axi_out_bvalid(arbiter_io_lsu_axi_out_bvalid),
    .io_axi_in_arready(arbiter_io_axi_in_arready),
    .io_axi_in_rdata(arbiter_io_axi_in_rdata),
    .io_axi_in_rvalid(arbiter_io_axi_in_rvalid),
    .io_axi_in_awready(arbiter_io_axi_in_awready),
    .io_axi_in_wready(arbiter_io_axi_in_wready),
    .io_axi_in_bvalid(arbiter_io_axi_in_bvalid),
    .io_axi_out_araddr(arbiter_io_axi_out_araddr),
    .io_axi_out_arvalid(arbiter_io_axi_out_arvalid),
    .io_axi_out_rready(arbiter_io_axi_out_rready),
    .io_axi_out_awaddr(arbiter_io_axi_out_awaddr),
    .io_axi_out_awvalid(arbiter_io_axi_out_awvalid),
    .io_axi_out_wdata(arbiter_io_axi_out_wdata),
    .io_axi_out_wstrb(arbiter_io_axi_out_wstrb),
    .io_axi_out_wvalid(arbiter_io_axi_out_wvalid),
    .io_axi_out_bready(arbiter_io_axi_out_bready)
  );
  IFU_AXI ifu_step ( // @[top.scala 21:26]
    .clock(ifu_step_clock),
    .reset(ifu_step_reset),
    .io_pc(ifu_step_io_pc),
    .io_pc_valid(ifu_step_io_pc_valid),
    .io_inst_valid(ifu_step_io_inst_valid),
    .io_inst(ifu_step_io_inst),
    .io_inst_reg(ifu_step_io_inst_reg),
    .io_axi_in_rdata(ifu_step_io_axi_in_rdata),
    .io_axi_in_rvalid(ifu_step_io_axi_in_rvalid),
    .io_axi_out_araddr(ifu_step_io_axi_out_araddr),
    .io_axi_out_arvalid(ifu_step_io_axi_out_arvalid),
    .io_axi_out_rready(ifu_step_io_axi_out_rready)
  );
  I_CACHE cache ( // @[top.scala 22:23]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_from_ifu_araddr(cache_io_from_ifu_araddr),
    .io_from_ifu_arvalid(cache_io_from_ifu_arvalid),
    .io_from_ifu_rready(cache_io_from_ifu_rready),
    .io_to_ifu_rdata(cache_io_to_ifu_rdata),
    .io_to_ifu_rvalid(cache_io_to_ifu_rvalid),
    .io_to_axi_araddr(cache_io_to_axi_araddr),
    .io_to_axi_arvalid(cache_io_to_axi_arvalid),
    .io_to_axi_rready(cache_io_to_axi_rready),
    .io_from_axi_rdata(cache_io_from_axi_rdata),
    .io_from_axi_rvalid(cache_io_from_axi_rvalid)
  );
  IDU idu_step ( // @[top.scala 39:26]
    .io_inst(idu_step_io_inst),
    .io_inst_now(idu_step_io_inst_now),
    .io_rs1(idu_step_io_rs1),
    .io_rs2(idu_step_io_rs2),
    .io_rd(idu_step_io_rd),
    .io_imm(idu_step_io_imm),
    .io_ctrl_sign_reg_write(idu_step_io_ctrl_sign_reg_write),
    .io_ctrl_sign_csr_write(idu_step_io_ctrl_sign_csr_write),
    .io_ctrl_sign_src2_is_imm(idu_step_io_ctrl_sign_src2_is_imm),
    .io_ctrl_sign_src1_is_pc(idu_step_io_ctrl_sign_src1_is_pc),
    .io_ctrl_sign_Writemem_en(idu_step_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(idu_step_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(idu_step_io_ctrl_sign_Wmask)
  );
  EXU_AXI exu_step ( // @[top.scala 44:26]
    .clock(exu_step_clock),
    .reset(exu_step_reset),
    .io_pc(exu_step_io_pc),
    .io_pc_next(exu_step_io_pc_next),
    .io_inst_now(exu_step_io_inst_now),
    .io_rs1(exu_step_io_rs1),
    .io_rs2(exu_step_io_rs2),
    .io_rd(exu_step_io_rd),
    .io_imm(exu_step_io_imm),
    .io_ctrl_sign_reg_write(exu_step_io_ctrl_sign_reg_write),
    .io_ctrl_sign_csr_write(exu_step_io_ctrl_sign_csr_write),
    .io_ctrl_sign_src2_is_imm(exu_step_io_ctrl_sign_src2_is_imm),
    .io_ctrl_sign_src1_is_pc(exu_step_io_ctrl_sign_src1_is_pc),
    .io_ctrl_sign_Writemem_en(exu_step_io_ctrl_sign_Writemem_en),
    .io_ctrl_sign_Readmem_en(exu_step_io_ctrl_sign_Readmem_en),
    .io_ctrl_sign_Wmask(exu_step_io_ctrl_sign_Wmask),
    .io_res2rd(exu_step_io_res2rd),
    .io_inst_valid(exu_step_io_inst_valid),
    .io_inst_store(exu_step_io_inst_store),
    .io_inst_load(exu_step_io_inst_load),
    .io_Mem_addr(exu_step_io_Mem_addr),
    .io_Mem_rdata(exu_step_io_Mem_rdata),
    .io_Mem_wdata(exu_step_io_Mem_wdata),
    .io_Mem_wstrb(exu_step_io_Mem_wstrb),
    .io_rdata_valid(exu_step_io_rdata_valid)
  );
  DPI dpi ( // @[top.scala 66:21]
    .flag(dpi_flag),
    .ecall_flag(dpi_ecall_flag)
  );
  assign io_inst = ifu_step_io_inst; // @[top.scala 24:13]
  assign io_pc = pc_now; // @[top.scala 16:11]
  assign io_pc_next = exu_step_io_pc_next; // @[top.scala 87:16]
  assign io_outval = exu_step_io_res2rd; // @[top.scala 62:15]
  assign io_step = diff_step; // @[top.scala 85:13]
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_axi_in_araddr = arbiter_io_axi_out_araddr; // @[top.scala 36:19]
  assign axi_io_axi_in_arvalid = arbiter_io_axi_out_arvalid; // @[top.scala 36:19]
  assign axi_io_axi_in_rready = arbiter_io_axi_out_rready; // @[top.scala 36:19]
  assign axi_io_axi_in_awaddr = arbiter_io_axi_out_awaddr; // @[top.scala 36:19]
  assign axi_io_axi_in_awvalid = arbiter_io_axi_out_awvalid; // @[top.scala 36:19]
  assign axi_io_axi_in_wdata = arbiter_io_axi_out_wdata; // @[top.scala 36:19]
  assign axi_io_axi_in_wstrb = arbiter_io_axi_out_wstrb; // @[top.scala 36:19]
  assign axi_io_axi_in_wvalid = arbiter_io_axi_out_wvalid; // @[top.scala 36:19]
  assign axi_io_axi_in_bready = arbiter_io_axi_out_bready; // @[top.scala 36:19]
  assign lsu_step_clock = clock;
  assign lsu_step_reset = reset;
  assign lsu_step_io_inst_store = exu_step_io_inst_store; // @[top.scala 54:28]
  assign lsu_step_io_inst_load = exu_step_io_inst_load; // @[top.scala 53:27]
  assign lsu_step_io_mem_addr = exu_step_io_Mem_addr; // @[top.scala 55:26]
  assign lsu_step_io_mem_wdata = exu_step_io_Mem_wdata; // @[top.scala 56:27]
  assign lsu_step_io_mem_wstrb = exu_step_io_Mem_wstrb; // @[top.scala 57:27]
  assign lsu_step_io_axi_in_arready = arbiter_io_lsu_axi_out_arready; // @[top.scala 34:24]
  assign lsu_step_io_axi_in_rdata = arbiter_io_lsu_axi_out_rdata; // @[top.scala 34:24]
  assign lsu_step_io_axi_in_rvalid = arbiter_io_lsu_axi_out_rvalid; // @[top.scala 34:24]
  assign lsu_step_io_axi_in_awready = arbiter_io_lsu_axi_out_awready; // @[top.scala 34:24]
  assign lsu_step_io_axi_in_wready = arbiter_io_lsu_axi_out_wready; // @[top.scala 34:24]
  assign lsu_step_io_axi_in_bvalid = arbiter_io_lsu_axi_out_bvalid; // @[top.scala 34:24]
  assign arbiter_clock = clock;
  assign arbiter_reset = reset;
  assign arbiter_io_ifu_axi_in_araddr = cache_io_to_axi_araddr; // @[top.scala 25:27]
  assign arbiter_io_ifu_axi_in_arvalid = cache_io_to_axi_arvalid; // @[top.scala 25:27]
  assign arbiter_io_ifu_axi_in_rready = cache_io_to_axi_rready; // @[top.scala 25:27]
  assign arbiter_io_lsu_axi_in_araddr = lsu_step_io_axi_out_araddr; // @[top.scala 33:27]
  assign arbiter_io_lsu_axi_in_arvalid = lsu_step_io_axi_out_arvalid; // @[top.scala 33:27]
  assign arbiter_io_lsu_axi_in_rready = lsu_step_io_axi_out_rready; // @[top.scala 33:27]
  assign arbiter_io_lsu_axi_in_awaddr = lsu_step_io_axi_out_awaddr; // @[top.scala 33:27]
  assign arbiter_io_lsu_axi_in_awvalid = lsu_step_io_axi_out_awvalid; // @[top.scala 33:27]
  assign arbiter_io_lsu_axi_in_wdata = lsu_step_io_axi_out_wdata; // @[top.scala 33:27]
  assign arbiter_io_lsu_axi_in_wstrb = lsu_step_io_axi_out_wstrb; // @[top.scala 33:27]
  assign arbiter_io_lsu_axi_in_wvalid = lsu_step_io_axi_out_wvalid; // @[top.scala 33:27]
  assign arbiter_io_lsu_axi_in_bready = lsu_step_io_axi_out_bready; // @[top.scala 33:27]
  assign arbiter_io_axi_in_arready = axi_io_axi_out_arready; // @[top.scala 35:23]
  assign arbiter_io_axi_in_rdata = axi_io_axi_out_rdata; // @[top.scala 35:23]
  assign arbiter_io_axi_in_rvalid = axi_io_axi_out_rvalid; // @[top.scala 35:23]
  assign arbiter_io_axi_in_awready = axi_io_axi_out_awready; // @[top.scala 35:23]
  assign arbiter_io_axi_in_wready = axi_io_axi_out_wready; // @[top.scala 35:23]
  assign arbiter_io_axi_in_bvalid = axi_io_axi_out_bvalid; // @[top.scala 35:23]
  assign ifu_step_clock = clock;
  assign ifu_step_reset = reset;
  assign ifu_step_io_pc = pc_now; // @[top.scala 23:20]
  assign ifu_step_io_pc_valid = pc_valid; // @[top.scala 82:26]
  assign ifu_step_io_axi_in_rdata = cache_io_to_ifu_rdata; // @[top.scala 27:24]
  assign ifu_step_io_axi_in_rvalid = cache_io_to_ifu_rvalid; // @[top.scala 27:24]
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_from_ifu_araddr = ifu_step_io_axi_out_araddr; // @[top.scala 28:23]
  assign cache_io_from_ifu_arvalid = ifu_step_io_axi_out_arvalid; // @[top.scala 28:23]
  assign cache_io_from_ifu_rready = ifu_step_io_axi_out_rready; // @[top.scala 28:23]
  assign cache_io_from_axi_rdata = arbiter_io_ifu_axi_out_rdata; // @[top.scala 26:23]
  assign cache_io_from_axi_rvalid = arbiter_io_ifu_axi_out_rvalid; // @[top.scala 26:23]
  assign idu_step_io_inst = ~ifu_step_io_inst_valid & ~pc_valid & ~execute_end ? ifu_step_io_inst_reg : ifu_step_io_inst
    ; // @[top.scala 89:28]
  assign exu_step_clock = clock;
  assign exu_step_reset = reset;
  assign exu_step_io_pc = pc_now; // @[top.scala 45:20]
  assign exu_step_io_inst_now = idu_step_io_inst_now; // @[top.scala 46:26]
  assign exu_step_io_rs1 = idu_step_io_rs1; // @[top.scala 48:21]
  assign exu_step_io_rs2 = idu_step_io_rs2; // @[top.scala 49:21]
  assign exu_step_io_rd = idu_step_io_rd; // @[top.scala 50:20]
  assign exu_step_io_imm = idu_step_io_imm; // @[top.scala 51:21]
  assign exu_step_io_ctrl_sign_reg_write = idu_step_io_ctrl_sign_reg_write; // @[top.scala 52:27]
  assign exu_step_io_ctrl_sign_csr_write = idu_step_io_ctrl_sign_csr_write; // @[top.scala 52:27]
  assign exu_step_io_ctrl_sign_src2_is_imm = idu_step_io_ctrl_sign_src2_is_imm; // @[top.scala 52:27]
  assign exu_step_io_ctrl_sign_src1_is_pc = idu_step_io_ctrl_sign_src1_is_pc; // @[top.scala 52:27]
  assign exu_step_io_ctrl_sign_Writemem_en = idu_step_io_ctrl_sign_Writemem_en; // @[top.scala 52:27]
  assign exu_step_io_ctrl_sign_Readmem_en = idu_step_io_ctrl_sign_Readmem_en; // @[top.scala 52:27]
  assign exu_step_io_ctrl_sign_Wmask = idu_step_io_ctrl_sign_Wmask; // @[top.scala 52:27]
  assign exu_step_io_inst_valid = ifu_step_io_inst_valid; // @[top.scala 61:28]
  assign exu_step_io_Mem_rdata = lsu_step_io_mem_rdata; // @[top.scala 58:27]
  assign exu_step_io_rdata_valid = lsu_step_io_axi_in_rvalid; // @[top.scala 59:29]
  assign dpi_flag = {{31'd0}, idu_step_io_inst_now == 32'h2}; // @[top.scala 67:17]
  assign dpi_ecall_flag = {{31'd0}, idu_step_io_inst_now == 32'h3d}; // @[top.scala 68:23]
  always @(posedge clock) begin
    if (reset) begin // @[top.scala 15:25]
      pc_now <= 64'h80000000; // @[top.scala 15:25]
    end else if (execute_end) begin // @[top.scala 86:18]
      pc_now <= exu_step_io_pc_next;
    end
    if (reset) begin // @[top.scala 17:30]
      execute_end <= 1'h0; // @[top.scala 17:30]
    end else if (exu_step_io_inst_store) begin // @[top.scala 78:23]
      execute_end <= lsu_step_io_axi_in_bvalid;
    end else if (exu_step_io_inst_load) begin // @[top.scala 78:76]
      execute_end <= lsu_step_io_axi_in_rvalid;
    end else begin
      execute_end <= ifu_step_io_inst_valid;
    end
    pc_valid <= reset | execute_end; // @[top.scala 80:{27,27} 81:14]
    if (reset) begin // @[top.scala 83:28]
      diff_step <= 1'h0; // @[top.scala 83:28]
    end else begin
      diff_step <= execute_end; // @[top.scala 84:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc_now = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  execute_end = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pc_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  diff_step = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
