module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [63:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_bvalid,
  output [31:0] io_to_axi_araddr,
  output [7:0]  io_to_axi_arlen,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output [7:0]  io_to_axi_awlen,
  output        io_to_axi_awvalid,
  output [63:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rlast,
  input         io_from_axi_rvalid,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [1023:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [1023:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
`endif // RANDOMIZE_REG_INIT
  reg [1023:0] cacheLine [0:63]; // @[d_cache.scala 24:24]
  wire  cacheLine_MPORT_1_en; // @[d_cache.scala 24:24]
  wire [5:0] cacheLine_MPORT_1_addr; // @[d_cache.scala 24:24]
  wire [1023:0] cacheLine_MPORT_1_data; // @[d_cache.scala 24:24]
  wire  cacheLine_write_back_data_MPORT_en; // @[d_cache.scala 24:24]
  wire [5:0] cacheLine_write_back_data_MPORT_addr; // @[d_cache.scala 24:24]
  wire [1023:0] cacheLine_write_back_data_MPORT_data; // @[d_cache.scala 24:24]
  wire  cacheLine_io_to_lsu_rdata_MPORT_en; // @[d_cache.scala 24:24]
  wire [5:0] cacheLine_io_to_lsu_rdata_MPORT_addr; // @[d_cache.scala 24:24]
  wire [1023:0] cacheLine_io_to_lsu_rdata_MPORT_data; // @[d_cache.scala 24:24]
  wire [1023:0] cacheLine_MPORT_data; // @[d_cache.scala 24:24]
  wire [5:0] cacheLine_MPORT_addr; // @[d_cache.scala 24:24]
  wire  cacheLine_MPORT_mask; // @[d_cache.scala 24:24]
  wire  cacheLine_MPORT_en; // @[d_cache.scala 24:24]
  wire [1023:0] cacheLine_MPORT_3_data; // @[d_cache.scala 24:24]
  wire [5:0] cacheLine_MPORT_3_addr; // @[d_cache.scala 24:24]
  wire  cacheLine_MPORT_3_mask; // @[d_cache.scala 24:24]
  wire  cacheLine_MPORT_3_en; // @[d_cache.scala 24:24]
  wire [1023:0] cacheLine_MPORT_6_data; // @[d_cache.scala 24:24]
  wire [5:0] cacheLine_MPORT_6_addr; // @[d_cache.scala 24:24]
  wire  cacheLine_MPORT_6_mask; // @[d_cache.scala 24:24]
  wire  cacheLine_MPORT_6_en; // @[d_cache.scala 24:24]
  reg  validMem [0:63]; // @[d_cache.scala 25:23]
  wire  validMem_valid_0_MPORT_en; // @[d_cache.scala 25:23]
  wire [5:0] validMem_valid_0_MPORT_addr; // @[d_cache.scala 25:23]
  wire  validMem_valid_0_MPORT_data; // @[d_cache.scala 25:23]
  wire  validMem_valid_1_MPORT_en; // @[d_cache.scala 25:23]
  wire [5:0] validMem_valid_1_MPORT_addr; // @[d_cache.scala 25:23]
  wire  validMem_valid_1_MPORT_data; // @[d_cache.scala 25:23]
  wire  validMem_valid_2_MPORT_en; // @[d_cache.scala 25:23]
  wire [5:0] validMem_valid_2_MPORT_addr; // @[d_cache.scala 25:23]
  wire  validMem_valid_2_MPORT_data; // @[d_cache.scala 25:23]
  wire  validMem_valid_3_MPORT_en; // @[d_cache.scala 25:23]
  wire [5:0] validMem_valid_3_MPORT_addr; // @[d_cache.scala 25:23]
  wire  validMem_valid_3_MPORT_data; // @[d_cache.scala 25:23]
  wire  validMem_MPORT_5_data; // @[d_cache.scala 25:23]
  wire [5:0] validMem_MPORT_5_addr; // @[d_cache.scala 25:23]
  wire  validMem_MPORT_5_mask; // @[d_cache.scala 25:23]
  wire  validMem_MPORT_5_en; // @[d_cache.scala 25:23]
  wire  validMem_MPORT_8_data; // @[d_cache.scala 25:23]
  wire [5:0] validMem_MPORT_8_addr; // @[d_cache.scala 25:23]
  wire  validMem_MPORT_8_mask; // @[d_cache.scala 25:23]
  wire  validMem_MPORT_8_en; // @[d_cache.scala 25:23]
  reg [31:0] tagMem [0:63]; // @[d_cache.scala 28:21]
  wire  tagMem_tagMatch_0_MPORT_en; // @[d_cache.scala 28:21]
  wire [5:0] tagMem_tagMatch_0_MPORT_addr; // @[d_cache.scala 28:21]
  wire [31:0] tagMem_tagMatch_0_MPORT_data; // @[d_cache.scala 28:21]
  wire  tagMem_tagMatch_1_MPORT_en; // @[d_cache.scala 28:21]
  wire [5:0] tagMem_tagMatch_1_MPORT_addr; // @[d_cache.scala 28:21]
  wire [31:0] tagMem_tagMatch_1_MPORT_data; // @[d_cache.scala 28:21]
  wire  tagMem_tagMatch_2_MPORT_en; // @[d_cache.scala 28:21]
  wire [5:0] tagMem_tagMatch_2_MPORT_addr; // @[d_cache.scala 28:21]
  wire [31:0] tagMem_tagMatch_2_MPORT_data; // @[d_cache.scala 28:21]
  wire  tagMem_tagMatch_3_MPORT_en; // @[d_cache.scala 28:21]
  wire [5:0] tagMem_tagMatch_3_MPORT_addr; // @[d_cache.scala 28:21]
  wire [31:0] tagMem_tagMatch_3_MPORT_data; // @[d_cache.scala 28:21]
  wire  tagMem_write_back_addr_MPORT_en; // @[d_cache.scala 28:21]
  wire [5:0] tagMem_write_back_addr_MPORT_addr; // @[d_cache.scala 28:21]
  wire [31:0] tagMem_write_back_addr_MPORT_data; // @[d_cache.scala 28:21]
  wire [31:0] tagMem_MPORT_4_data; // @[d_cache.scala 28:21]
  wire [5:0] tagMem_MPORT_4_addr; // @[d_cache.scala 28:21]
  wire  tagMem_MPORT_4_mask; // @[d_cache.scala 28:21]
  wire  tagMem_MPORT_4_en; // @[d_cache.scala 28:21]
  wire [31:0] tagMem_MPORT_7_data; // @[d_cache.scala 28:21]
  wire [5:0] tagMem_MPORT_7_addr; // @[d_cache.scala 28:21]
  wire  tagMem_MPORT_7_mask; // @[d_cache.scala 28:21]
  wire  tagMem_MPORT_7_en; // @[d_cache.scala 28:21]
  reg  dirtyMem [0:63]; // @[d_cache.scala 29:23]
  wire  dirtyMem_MPORT_9_en; // @[d_cache.scala 29:23]
  wire [5:0] dirtyMem_MPORT_9_addr; // @[d_cache.scala 29:23]
  wire  dirtyMem_MPORT_9_data; // @[d_cache.scala 29:23]
  wire  dirtyMem_MPORT_2_data; // @[d_cache.scala 29:23]
  wire [5:0] dirtyMem_MPORT_2_addr; // @[d_cache.scala 29:23]
  wire  dirtyMem_MPORT_2_mask; // @[d_cache.scala 29:23]
  wire  dirtyMem_MPORT_2_en; // @[d_cache.scala 29:23]
  wire  dirtyMem_MPORT_10_data; // @[d_cache.scala 29:23]
  wire [5:0] dirtyMem_MPORT_10_addr; // @[d_cache.scala 29:23]
  wire  dirtyMem_MPORT_10_mask; // @[d_cache.scala 29:23]
  wire  dirtyMem_MPORT_10_en; // @[d_cache.scala 29:23]
  wire [6:0] offset = io_from_lsu_araddr[6:0]; // @[d_cache.scala 20:36]
  wire [3:0] index = io_from_lsu_araddr[10:7]; // @[d_cache.scala 21:35]
  wire [20:0] tag = io_from_lsu_araddr[31:11]; // @[d_cache.scala 22:33]
  wire [7:0] _GEN_503 = {{4'd0}, index}; // @[d_cache.scala 41:48]
  wire [8:0] _valid_0_T_1 = {{1'd0}, _GEN_503}; // @[d_cache.scala 41:48]
  wire [7:0] _valid_1_T_2 = 8'h10 + _GEN_503; // @[d_cache.scala 41:48]
  wire [8:0] _GEN_507 = {{5'd0}, index}; // @[d_cache.scala 41:48]
  wire [8:0] _valid_2_T_2 = 9'h20 + _GEN_507; // @[d_cache.scala 41:48]
  wire [8:0] _valid_3_T_2 = 9'h30 + _GEN_507; // @[d_cache.scala 41:48]
  wire  valid_0 = validMem_valid_0_MPORT_data; // @[d_cache.scala 39:21 41:18]
  wire  valid_1 = validMem_valid_1_MPORT_data; // @[d_cache.scala 39:21 41:18]
  wire  valid_2 = validMem_valid_2_MPORT_data; // @[d_cache.scala 39:21 41:18]
  wire  valid_3 = validMem_valid_3_MPORT_data; // @[d_cache.scala 39:21 41:18]
  wire  allvalid = valid_0 & valid_1 & valid_2 & valid_3; // @[d_cache.scala 43:35]
  wire  _foundUnvalidIndex_T = ~valid_0; // @[d_cache.scala 45:10]
  wire  _foundUnvalidIndex_T_1 = ~valid_1; // @[d_cache.scala 46:10]
  wire  _foundUnvalidIndex_T_2 = ~valid_2; // @[d_cache.scala 47:10]
  wire  _foundUnvalidIndex_T_3 = ~valid_3; // @[d_cache.scala 48:10]
  wire [1:0] _foundUnvalidIndex_T_4 = _foundUnvalidIndex_T_3 ? 2'h3 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _foundUnvalidIndex_T_5 = _foundUnvalidIndex_T_2 ? 2'h2 : _foundUnvalidIndex_T_4; // @[Mux.scala 101:16]
  wire [1:0] _foundUnvalidIndex_T_6 = _foundUnvalidIndex_T_1 ? 2'h1 : _foundUnvalidIndex_T_5; // @[Mux.scala 101:16]
  wire [1:0] foundUnvalidIndex = _foundUnvalidIndex_T ? 2'h0 : _foundUnvalidIndex_T_6; // @[Mux.scala 101:16]
  wire [5:0] _GEN_512 = {foundUnvalidIndex, 4'h0}; // @[d_cache.scala 50:43]
  wire [8:0] _unvalidIndex_T = {{3'd0}, _GEN_512}; // @[d_cache.scala 50:43]
  wire [8:0] unvalidIndex = _unvalidIndex_T + _GEN_507; // @[d_cache.scala 50:51]
  wire [31:0] _GEN_519 = {{11'd0}, tag}; // @[d_cache.scala 55:71]
  wire  tagMatch_0 = valid_0 & tagMem_tagMatch_0_MPORT_data == _GEN_519; // @[d_cache.scala 55:33]
  wire  tagMatch_1 = valid_1 & tagMem_tagMatch_1_MPORT_data == _GEN_519; // @[d_cache.scala 55:33]
  wire  tagMatch_2 = valid_2 & tagMem_tagMatch_2_MPORT_data == _GEN_519; // @[d_cache.scala 55:33]
  wire  tagMatch_3 = valid_3 & tagMem_tagMatch_3_MPORT_data == _GEN_519; // @[d_cache.scala 55:33]
  wire  anyMatch = tagMatch_0 | tagMatch_1 | tagMatch_2 | tagMatch_3; // @[d_cache.scala 57:38]
  wire [1:0] _foundtagIndex_T = tagMatch_3 ? 2'h3 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _foundtagIndex_T_1 = tagMatch_2 ? 2'h2 : _foundtagIndex_T; // @[Mux.scala 101:16]
  wire [1:0] _foundtagIndex_T_2 = tagMatch_1 ? 2'h1 : _foundtagIndex_T_1; // @[Mux.scala 101:16]
  wire [1:0] foundtagIndex = tagMatch_0 ? 2'h0 : _foundtagIndex_T_2; // @[Mux.scala 101:16]
  wire [5:0] _GEN_537 = {foundtagIndex, 4'h0}; // @[d_cache.scala 64:35]
  wire [8:0] _tagIndex_T = {{3'd0}, _GEN_537}; // @[d_cache.scala 64:35]
  wire [8:0] tagIndex = _tagIndex_T + _GEN_507; // @[d_cache.scala 64:43]
  reg [1023:0] write_back_data; // @[d_cache.scala 70:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 71:34]
  reg [63:0] receive_data_0; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_1; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_2; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_3; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_4; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_5; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_6; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_7; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_8; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_9; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_10; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_11; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_12; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_13; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_14; // @[d_cache.scala 75:31]
  reg [63:0] receive_data_15; // @[d_cache.scala 75:31]
  reg [2:0] receive_num; // @[d_cache.scala 76:30]
  reg [7:0] quene_0; // @[d_cache.scala 77:24]
  reg [7:0] quene_1; // @[d_cache.scala 77:24]
  reg [7:0] quene_2; // @[d_cache.scala 77:24]
  reg [7:0] quene_3; // @[d_cache.scala 77:24]
  reg [7:0] quene_4; // @[d_cache.scala 77:24]
  reg [7:0] quene_5; // @[d_cache.scala 77:24]
  reg [7:0] quene_6; // @[d_cache.scala 77:24]
  reg [7:0] quene_7; // @[d_cache.scala 77:24]
  reg [7:0] quene_8; // @[d_cache.scala 77:24]
  reg [7:0] quene_9; // @[d_cache.scala 77:24]
  reg [7:0] quene_10; // @[d_cache.scala 77:24]
  reg [7:0] quene_11; // @[d_cache.scala 77:24]
  reg [7:0] quene_12; // @[d_cache.scala 77:24]
  reg [7:0] quene_13; // @[d_cache.scala 77:24]
  reg [7:0] quene_14; // @[d_cache.scala 77:24]
  reg [7:0] quene_15; // @[d_cache.scala 77:24]
  wire [7:0] _GEN_1 = 4'h1 == index ? quene_1 : quene_0; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_2 = 4'h2 == index ? quene_2 : _GEN_1; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_3 = 4'h3 == index ? quene_3 : _GEN_2; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_4 = 4'h4 == index ? quene_4 : _GEN_3; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_5 = 4'h5 == index ? quene_5 : _GEN_4; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_6 = 4'h6 == index ? quene_6 : _GEN_5; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_7 = 4'h7 == index ? quene_7 : _GEN_6; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_8 = 4'h8 == index ? quene_8 : _GEN_7; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_9 = 4'h9 == index ? quene_9 : _GEN_8; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_10 = 4'ha == index ? quene_10 : _GEN_9; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_11 = 4'hb == index ? quene_11 : _GEN_10; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_12 = 4'hc == index ? quene_12 : _GEN_11; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_13 = 4'hd == index ? quene_13 : _GEN_12; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_14 = 4'he == index ? quene_14 : _GEN_13; // @[d_cache.scala 79:{35,35}]
  wire [7:0] _GEN_15 = 4'hf == index ? quene_15 : _GEN_14; // @[d_cache.scala 79:{35,35}]
  wire [1:0] replace_way = _GEN_15[7:6]; // @[d_cache.scala 79:35]
  wire [5:0] _GEN_543 = {replace_way, 4'h0}; // @[d_cache.scala 80:34]
  wire [8:0] _replaceIndex_T = {{3'd0}, _GEN_543}; // @[d_cache.scala 80:34]
  wire [8:0] _replaceIndex_T_2 = _replaceIndex_T + _GEN_507; // @[d_cache.scala 80:42]
  wire [9:0] shift_bit = {offset, 3'h0}; // @[d_cache.scala 82:28]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 88:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 87:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 86:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 85:20]
  reg [2:0] state; // @[d_cache.scala 95:24]
  wire  _T = 3'h0 == state; // @[d_cache.scala 101:18]
  wire  _T_3 = (io_from_lsu_arvalid | io_from_lsu_awvalid) & io_from_lsu_araddr >= 32'ha0000000; // @[d_cache.scala 103:60]
  wire [2:0] _GEN_16 = io_from_lsu_awvalid ? 3'h2 : state; // @[d_cache.scala 107:44 108:23 95:24]
  wire [63:0] _T_7 = io_from_lsu_wdata & wmask; // @[d_cache.scala 127:60]
  wire [1086:0] _GEN_589 = {{1023'd0}, _T_7}; // @[d_cache.scala 127:69]
  wire [1086:0] _T_8 = _GEN_589 << shift_bit; // @[d_cache.scala 127:69]
  wire [1086:0] _GEN_592 = {{1023'd0}, wmask}; // @[d_cache.scala 127:116]
  wire [1086:0] _T_10 = _GEN_592 << shift_bit; // @[d_cache.scala 127:116]
  wire [1086:0] _T_11 = ~_T_10; // @[d_cache.scala 127:108]
  wire [1086:0] _GEN_550 = {{63'd0}, cacheLine_MPORT_1_data}; // @[d_cache.scala 127:106]
  wire [1086:0] _T_12 = _GEN_550 & _T_11; // @[d_cache.scala 127:106]
  wire [1086:0] _T_13 = _T_8 | _T_12; // @[d_cache.scala 127:83]
  wire [2:0] _GEN_23 = anyMatch ? 3'h0 : 3'h4; // @[d_cache.scala 122:27 131:23]
  wire [63:0] _GEN_31 = 3'h0 == receive_num ? io_from_axi_rdata : receive_data_0; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_32 = 3'h1 == receive_num ? io_from_axi_rdata : receive_data_1; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_33 = 3'h2 == receive_num ? io_from_axi_rdata : receive_data_2; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_34 = 3'h3 == receive_num ? io_from_axi_rdata : receive_data_3; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_35 = 3'h4 == receive_num ? io_from_axi_rdata : receive_data_4; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_36 = 3'h5 == receive_num ? io_from_axi_rdata : receive_data_5; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_37 = 3'h6 == receive_num ? io_from_axi_rdata : receive_data_6; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_38 = 3'h7 == receive_num ? io_from_axi_rdata : receive_data_7; // @[d_cache.scala 136:{43,43} 75:31]
  wire [3:0] _GEN_552 = {{1'd0}, receive_num}; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_39 = 4'h8 == _GEN_552 ? io_from_axi_rdata : receive_data_8; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_40 = 4'h9 == _GEN_552 ? io_from_axi_rdata : receive_data_9; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_41 = 4'ha == _GEN_552 ? io_from_axi_rdata : receive_data_10; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_42 = 4'hb == _GEN_552 ? io_from_axi_rdata : receive_data_11; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_43 = 4'hc == _GEN_552 ? io_from_axi_rdata : receive_data_12; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_44 = 4'hd == _GEN_552 ? io_from_axi_rdata : receive_data_13; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_45 = 4'he == _GEN_552 ? io_from_axi_rdata : receive_data_14; // @[d_cache.scala 136:{43,43} 75:31]
  wire [63:0] _GEN_46 = 4'hf == _GEN_552 ? io_from_axi_rdata : receive_data_15; // @[d_cache.scala 136:{43,43} 75:31]
  wire [2:0] _receive_num_T_1 = receive_num + 3'h1; // @[d_cache.scala 137:44]
  wire [2:0] _GEN_47 = io_from_axi_rlast ? 3'h5 : state; // @[d_cache.scala 138:40 139:27 95:24]
  wire [63:0] _GEN_48 = io_from_axi_rvalid ? _GEN_31 : receive_data_0; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_49 = io_from_axi_rvalid ? _GEN_32 : receive_data_1; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_50 = io_from_axi_rvalid ? _GEN_33 : receive_data_2; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_51 = io_from_axi_rvalid ? _GEN_34 : receive_data_3; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_52 = io_from_axi_rvalid ? _GEN_35 : receive_data_4; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_53 = io_from_axi_rvalid ? _GEN_36 : receive_data_5; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_54 = io_from_axi_rvalid ? _GEN_37 : receive_data_6; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_55 = io_from_axi_rvalid ? _GEN_38 : receive_data_7; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_56 = io_from_axi_rvalid ? _GEN_39 : receive_data_8; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_57 = io_from_axi_rvalid ? _GEN_40 : receive_data_9; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_58 = io_from_axi_rvalid ? _GEN_41 : receive_data_10; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_59 = io_from_axi_rvalid ? _GEN_42 : receive_data_11; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_60 = io_from_axi_rvalid ? _GEN_43 : receive_data_12; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_61 = io_from_axi_rvalid ? _GEN_44 : receive_data_13; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_62 = io_from_axi_rvalid ? _GEN_45 : receive_data_14; // @[d_cache.scala 135:37 75:31]
  wire [63:0] _GEN_63 = io_from_axi_rvalid ? _GEN_46 : receive_data_15; // @[d_cache.scala 135:37 75:31]
  wire [2:0] _GEN_64 = io_from_axi_rvalid ? _receive_num_T_1 : receive_num; // @[d_cache.scala 135:37 137:29 76:30]
  wire [2:0] _GEN_65 = io_from_axi_rvalid ? _GEN_47 : state; // @[d_cache.scala 135:37 95:24]
  wire [2:0] _GEN_66 = io_from_axi_bvalid ? 3'h0 : state; // @[d_cache.scala 144:59 145:23 95:24]
  wire  _T_19 = ~allvalid; // @[d_cache.scala 149:18]
  wire [511:0] lo = {receive_data_7,receive_data_6,receive_data_5,receive_data_4,receive_data_3,receive_data_2,
    receive_data_1,receive_data_0}; // @[Cat.scala 31:58]
  wire [511:0] hi = {receive_data_15,receive_data_14,receive_data_13,receive_data_12,receive_data_11,receive_data_10,
    receive_data_9,receive_data_8}; // @[Cat.scala 31:58]
  wire [9:0] _GEN_573 = {_GEN_15, 2'h0}; // @[d_cache.scala 157:46]
  wire [10:0] _quene_T = {{1'd0}, _GEN_573}; // @[d_cache.scala 157:46]
  wire [10:0] _GEN_575 = {{9'd0}, foundUnvalidIndex}; // @[d_cache.scala 157:53]
  wire [10:0] _quene_T_1 = _quene_T | _GEN_575; // @[d_cache.scala 157:53]
  wire [7:0] _GEN_67 = 4'h0 == index ? _quene_T_1[7:0] : quene_0; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_68 = 4'h1 == index ? _quene_T_1[7:0] : quene_1; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_69 = 4'h2 == index ? _quene_T_1[7:0] : quene_2; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_70 = 4'h3 == index ? _quene_T_1[7:0] : quene_3; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_71 = 4'h4 == index ? _quene_T_1[7:0] : quene_4; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_72 = 4'h5 == index ? _quene_T_1[7:0] : quene_5; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_73 = 4'h6 == index ? _quene_T_1[7:0] : quene_6; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_74 = 4'h7 == index ? _quene_T_1[7:0] : quene_7; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_75 = 4'h8 == index ? _quene_T_1[7:0] : quene_8; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_76 = 4'h9 == index ? _quene_T_1[7:0] : quene_9; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_77 = 4'ha == index ? _quene_T_1[7:0] : quene_10; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_78 = 4'hb == index ? _quene_T_1[7:0] : quene_11; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_79 = 4'hc == index ? _quene_T_1[7:0] : quene_12; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_80 = 4'hd == index ? _quene_T_1[7:0] : quene_13; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_81 = 4'he == index ? _quene_T_1[7:0] : quene_14; // @[d_cache.scala 157:{30,30} 77:24]
  wire [7:0] _GEN_82 = 4'hf == index ? _quene_T_1[7:0] : quene_15; // @[d_cache.scala 157:{30,30} 77:24]
  wire [31:0] replaceIndex = {{23'd0}, _replaceIndex_T_2}; // @[d_cache.scala 66:28 80:18]
  wire [10:0] _GEN_578 = {{9'd0}, replace_way}; // @[d_cache.scala 162:53]
  wire [10:0] _quene_T_3 = _quene_T | _GEN_578; // @[d_cache.scala 162:53]
  wire [7:0] _GEN_83 = 4'h0 == index ? _quene_T_3[7:0] : quene_0; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_84 = 4'h1 == index ? _quene_T_3[7:0] : quene_1; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_85 = 4'h2 == index ? _quene_T_3[7:0] : quene_2; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_86 = 4'h3 == index ? _quene_T_3[7:0] : quene_3; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_87 = 4'h4 == index ? _quene_T_3[7:0] : quene_4; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_88 = 4'h5 == index ? _quene_T_3[7:0] : quene_5; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_89 = 4'h6 == index ? _quene_T_3[7:0] : quene_6; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_90 = 4'h7 == index ? _quene_T_3[7:0] : quene_7; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_91 = 4'h8 == index ? _quene_T_3[7:0] : quene_8; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_92 = 4'h9 == index ? _quene_T_3[7:0] : quene_9; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_93 = 4'ha == index ? _quene_T_3[7:0] : quene_10; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_94 = 4'hb == index ? _quene_T_3[7:0] : quene_11; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_95 = 4'hc == index ? _quene_T_3[7:0] : quene_12; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_96 = 4'hd == index ? _quene_T_3[7:0] : quene_13; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_97 = 4'he == index ? _quene_T_3[7:0] : quene_14; // @[d_cache.scala 162:{30,30} 77:24]
  wire [7:0] _GEN_98 = 4'hf == index ? _quene_T_3[7:0] : quene_15; // @[d_cache.scala 162:{30,30} 77:24]
  wire  _T_29 = dirtyMem_MPORT_9_data; // @[d_cache.scala 163:44]
  wire [42:0] _write_back_addr_T_2 = {tagMem_write_back_addr_MPORT_data,index,7'h0}; // @[Cat.scala 31:58]
  wire [1023:0] _GEN_102 = dirtyMem_MPORT_9_data ? cacheLine_write_back_data_MPORT_data : write_back_data; // @[d_cache.scala 163:51 165:37 70:34]
  wire [42:0] _GEN_104 = dirtyMem_MPORT_9_data ? _write_back_addr_T_2 : {{11'd0}, write_back_addr}; // @[d_cache.scala 163:51 166:37 71:34]
  wire [2:0] _GEN_108 = dirtyMem_MPORT_9_data ? 3'h6 : 3'h1; // @[d_cache.scala 163:51 168:27 170:27]
  wire [2:0] _GEN_109 = ~allvalid ? 3'h1 : _GEN_108; // @[d_cache.scala 149:28 150:23]
  wire [7:0] _GEN_118 = ~allvalid ? _GEN_67 : _GEN_83; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_119 = ~allvalid ? _GEN_68 : _GEN_84; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_120 = ~allvalid ? _GEN_69 : _GEN_85; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_121 = ~allvalid ? _GEN_70 : _GEN_86; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_122 = ~allvalid ? _GEN_71 : _GEN_87; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_123 = ~allvalid ? _GEN_72 : _GEN_88; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_124 = ~allvalid ? _GEN_73 : _GEN_89; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_125 = ~allvalid ? _GEN_74 : _GEN_90; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_126 = ~allvalid ? _GEN_75 : _GEN_91; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_127 = ~allvalid ? _GEN_76 : _GEN_92; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_128 = ~allvalid ? _GEN_77 : _GEN_93; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_129 = ~allvalid ? _GEN_78 : _GEN_94; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_130 = ~allvalid ? _GEN_79 : _GEN_95; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_131 = ~allvalid ? _GEN_80 : _GEN_96; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_132 = ~allvalid ? _GEN_81 : _GEN_97; // @[d_cache.scala 149:28]
  wire [7:0] _GEN_133 = ~allvalid ? _GEN_82 : _GEN_98; // @[d_cache.scala 149:28]
  wire  _GEN_136 = ~allvalid ? 1'h0 : 1'h1; // @[d_cache.scala 149:28 24:24 159:26]
  wire  _GEN_145 = ~allvalid ? 1'h0 : _T_29; // @[d_cache.scala 149:28 24:24]
  wire [1023:0] _GEN_146 = ~allvalid ? write_back_data : _GEN_102; // @[d_cache.scala 149:28 70:34]
  wire [42:0] _GEN_148 = ~allvalid ? {{11'd0}, write_back_addr} : _GEN_104; // @[d_cache.scala 149:28 71:34]
  wire [1023:0] _write_back_data_T_1 = {{64'd0}, write_back_data[1023:64]}; // @[d_cache.scala 176:52]
  wire [1023:0] _GEN_152 = io_from_axi_wready ? _write_back_data_T_1 : write_back_data; // @[d_cache.scala 175:37 176:33 70:34]
  wire [2:0] _GEN_153 = io_from_axi_bvalid ? 3'h1 : state; // @[d_cache.scala 178:37 179:23 95:24]
  wire [1023:0] _GEN_154 = 3'h6 == state ? _GEN_152 : write_back_data; // @[d_cache.scala 101:18 70:34]
  wire [2:0] _GEN_155 = 3'h6 == state ? _GEN_153 : state; // @[d_cache.scala 101:18 95:24]
  wire [2:0] _GEN_156 = 3'h5 == state ? _GEN_109 : _GEN_155; // @[d_cache.scala 101:18]
  wire [7:0] _GEN_165 = 3'h5 == state ? _GEN_118 : quene_0; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_166 = 3'h5 == state ? _GEN_119 : quene_1; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_167 = 3'h5 == state ? _GEN_120 : quene_2; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_168 = 3'h5 == state ? _GEN_121 : quene_3; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_169 = 3'h5 == state ? _GEN_122 : quene_4; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_170 = 3'h5 == state ? _GEN_123 : quene_5; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_171 = 3'h5 == state ? _GEN_124 : quene_6; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_172 = 3'h5 == state ? _GEN_125 : quene_7; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_173 = 3'h5 == state ? _GEN_126 : quene_8; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_174 = 3'h5 == state ? _GEN_127 : quene_9; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_175 = 3'h5 == state ? _GEN_128 : quene_10; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_176 = 3'h5 == state ? _GEN_129 : quene_11; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_177 = 3'h5 == state ? _GEN_130 : quene_12; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_178 = 3'h5 == state ? _GEN_131 : quene_13; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_179 = 3'h5 == state ? _GEN_132 : quene_14; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_180 = 3'h5 == state ? _GEN_133 : quene_15; // @[d_cache.scala 101:18 77:24]
  wire [1023:0] _GEN_193 = 3'h5 == state ? _GEN_146 : _GEN_154; // @[d_cache.scala 101:18]
  wire [42:0] _GEN_195 = 3'h5 == state ? _GEN_148 : {{11'd0}, write_back_addr}; // @[d_cache.scala 101:18 71:34]
  wire [2:0] _GEN_199 = 3'h4 == state ? _GEN_66 : _GEN_156; // @[d_cache.scala 101:18]
  wire  _GEN_202 = 3'h4 == state ? 1'h0 : 3'h5 == state & _T_19; // @[d_cache.scala 101:18 24:24]
  wire [7:0] _GEN_208 = 3'h4 == state ? quene_0 : _GEN_165; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_209 = 3'h4 == state ? quene_1 : _GEN_166; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_210 = 3'h4 == state ? quene_2 : _GEN_167; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_211 = 3'h4 == state ? quene_3 : _GEN_168; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_212 = 3'h4 == state ? quene_4 : _GEN_169; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_213 = 3'h4 == state ? quene_5 : _GEN_170; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_214 = 3'h4 == state ? quene_6 : _GEN_171; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_215 = 3'h4 == state ? quene_7 : _GEN_172; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_216 = 3'h4 == state ? quene_8 : _GEN_173; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_217 = 3'h4 == state ? quene_9 : _GEN_174; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_218 = 3'h4 == state ? quene_10 : _GEN_175; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_219 = 3'h4 == state ? quene_11 : _GEN_176; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_220 = 3'h4 == state ? quene_12 : _GEN_177; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_221 = 3'h4 == state ? quene_13 : _GEN_178; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_222 = 3'h4 == state ? quene_14 : _GEN_179; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_223 = 3'h4 == state ? quene_15 : _GEN_180; // @[d_cache.scala 101:18 77:24]
  wire  _GEN_226 = 3'h4 == state ? 1'h0 : 3'h5 == state & _GEN_136; // @[d_cache.scala 101:18 24:24]
  wire  _GEN_235 = 3'h4 == state ? 1'h0 : 3'h5 == state & _GEN_145; // @[d_cache.scala 101:18 24:24]
  wire [1023:0] _GEN_236 = 3'h4 == state ? write_back_data : _GEN_193; // @[d_cache.scala 101:18 70:34]
  wire [42:0] _GEN_238 = 3'h4 == state ? {{11'd0}, write_back_addr} : _GEN_195; // @[d_cache.scala 101:18 71:34]
  wire [63:0] _GEN_242 = 3'h3 == state ? _GEN_48 : receive_data_0; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_243 = 3'h3 == state ? _GEN_49 : receive_data_1; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_244 = 3'h3 == state ? _GEN_50 : receive_data_2; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_245 = 3'h3 == state ? _GEN_51 : receive_data_3; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_246 = 3'h3 == state ? _GEN_52 : receive_data_4; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_247 = 3'h3 == state ? _GEN_53 : receive_data_5; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_248 = 3'h3 == state ? _GEN_54 : receive_data_6; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_249 = 3'h3 == state ? _GEN_55 : receive_data_7; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_250 = 3'h3 == state ? _GEN_56 : receive_data_8; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_251 = 3'h3 == state ? _GEN_57 : receive_data_9; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_252 = 3'h3 == state ? _GEN_58 : receive_data_10; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_253 = 3'h3 == state ? _GEN_59 : receive_data_11; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_254 = 3'h3 == state ? _GEN_60 : receive_data_12; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_255 = 3'h3 == state ? _GEN_61 : receive_data_13; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_256 = 3'h3 == state ? _GEN_62 : receive_data_14; // @[d_cache.scala 101:18 75:31]
  wire [63:0] _GEN_257 = 3'h3 == state ? _GEN_63 : receive_data_15; // @[d_cache.scala 101:18 75:31]
  wire [2:0] _GEN_258 = 3'h3 == state ? _GEN_64 : receive_num; // @[d_cache.scala 101:18 76:30]
  wire [2:0] _GEN_259 = 3'h3 == state ? _GEN_65 : _GEN_199; // @[d_cache.scala 101:18]
  wire  _GEN_262 = 3'h3 == state ? 1'h0 : _GEN_202; // @[d_cache.scala 101:18 24:24]
  wire [7:0] _GEN_268 = 3'h3 == state ? quene_0 : _GEN_208; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_269 = 3'h3 == state ? quene_1 : _GEN_209; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_270 = 3'h3 == state ? quene_2 : _GEN_210; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_271 = 3'h3 == state ? quene_3 : _GEN_211; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_272 = 3'h3 == state ? quene_4 : _GEN_212; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_273 = 3'h3 == state ? quene_5 : _GEN_213; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_274 = 3'h3 == state ? quene_6 : _GEN_214; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_275 = 3'h3 == state ? quene_7 : _GEN_215; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_276 = 3'h3 == state ? quene_8 : _GEN_216; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_277 = 3'h3 == state ? quene_9 : _GEN_217; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_278 = 3'h3 == state ? quene_10 : _GEN_218; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_279 = 3'h3 == state ? quene_11 : _GEN_219; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_280 = 3'h3 == state ? quene_12 : _GEN_220; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_281 = 3'h3 == state ? quene_13 : _GEN_221; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_282 = 3'h3 == state ? quene_14 : _GEN_222; // @[d_cache.scala 101:18 77:24]
  wire [7:0] _GEN_283 = 3'h3 == state ? quene_15 : _GEN_223; // @[d_cache.scala 101:18 77:24]
  wire  _GEN_286 = 3'h3 == state ? 1'h0 : _GEN_226; // @[d_cache.scala 101:18 24:24]
  wire  _GEN_295 = 3'h3 == state ? 1'h0 : _GEN_235; // @[d_cache.scala 101:18 24:24]
  wire [1023:0] _GEN_296 = 3'h3 == state ? write_back_data : _GEN_236; // @[d_cache.scala 101:18 70:34]
  wire [42:0] _GEN_298 = 3'h3 == state ? {{11'd0}, write_back_addr} : _GEN_238; // @[d_cache.scala 101:18 71:34]
  wire  _GEN_329 = 3'h2 == state ? 1'h0 : _GEN_262; // @[d_cache.scala 101:18 24:24]
  wire  _GEN_353 = 3'h2 == state ? 1'h0 : _GEN_286; // @[d_cache.scala 101:18 24:24]
  wire  _GEN_362 = 3'h2 == state ? 1'h0 : _GEN_295; // @[d_cache.scala 101:18 24:24]
  wire [42:0] _GEN_365 = 3'h2 == state ? {{11'd0}, write_back_addr} : _GEN_298; // @[d_cache.scala 101:18 71:34]
  wire  _GEN_373 = 3'h1 == state ? 1'h0 : 3'h2 == state & anyMatch; // @[d_cache.scala 101:18 24:24]
  wire  _GEN_396 = 3'h1 == state ? 1'h0 : _GEN_329; // @[d_cache.scala 101:18 24:24]
  wire  _GEN_420 = 3'h1 == state ? 1'h0 : _GEN_353; // @[d_cache.scala 101:18 24:24]
  wire  _GEN_429 = 3'h1 == state ? 1'h0 : _GEN_362; // @[d_cache.scala 101:18 24:24]
  wire [42:0] _GEN_432 = 3'h1 == state ? {{11'd0}, write_back_addr} : _GEN_365; // @[d_cache.scala 101:18 71:34]
  wire [42:0] _GEN_499 = 3'h0 == state ? {{11'd0}, write_back_addr} : _GEN_432; // @[d_cache.scala 101:18 71:34]
  wire [1023:0] _io_to_lsu_rdata_T_1 = cacheLine_io_to_lsu_rdata_MPORT_data >> shift_bit; // @[d_cache.scala 201:48]
  wire [63:0] _GEN_583 = {{32'd0}, io_from_lsu_araddr}; // @[d_cache.scala 242:49]
  wire [63:0] _io_to_axi_araddr_T = _GEN_583 & 64'hffffffffffffff80; // @[d_cache.scala 242:49]
  wire  _T_41 = state == 3'h0 & _T_3; // @[d_cache.scala 307:27]
  wire [63:0] _GEN_504 = state == 3'h0 & _T_3 ? io_from_axi_rdata : 64'h0; // @[d_cache.scala 307:117 308:23 311:29]
  wire  _GEN_506 = state == 3'h0 & _T_3 & io_from_axi_rvalid; // @[d_cache.scala 307:117 308:23 313:30]
  wire  _GEN_509 = state == 3'h0 & _T_3 & io_from_axi_bvalid; // @[d_cache.scala 307:117 308:23 316:30]
  wire  _GEN_514 = state == 3'h0 & _T_3 & io_from_lsu_arvalid; // @[d_cache.scala 307:117 309:23 318:31]
  wire [31:0] _GEN_516 = state == 3'h0 & _T_3 ? io_from_lsu_awaddr : 32'h0; // @[d_cache.scala 307:117 309:23 324:30]
  wire  _GEN_520 = state == 3'h0 & _T_3 & io_from_lsu_awvalid; // @[d_cache.scala 307:117 309:23 325:31]
  wire [63:0] _GEN_521 = state == 3'h0 & _T_3 ? io_from_lsu_wdata : 64'h0; // @[d_cache.scala 307:117 309:23 329:29]
  wire [7:0] _GEN_522 = state == 3'h0 & _T_3 ? io_from_lsu_wstrb : 8'h0; // @[d_cache.scala 307:117 309:23 330:29]
  wire  _GEN_524 = state == 3'h0 & _T_3 & io_from_lsu_wvalid; // @[d_cache.scala 307:117 309:23 332:30]
  wire [63:0] _GEN_526 = state == 3'h6 ? 64'h0 : _GEN_504; // @[d_cache.scala 282:35 283:25]
  wire  _GEN_528 = state == 3'h6 ? 1'h0 : _GEN_506; // @[d_cache.scala 282:35 285:26]
  wire  _GEN_531 = state == 3'h6 ? 1'h0 : _GEN_509; // @[d_cache.scala 282:35 288:26]
  wire  _GEN_533 = state == 3'h6 ? 1'h0 : _GEN_514; // @[d_cache.scala 282:35 290:27]
  wire [31:0] _GEN_534 = state == 3'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 282:35 291:26]
  wire  _GEN_538 = state == 3'h6 ? 1'h0 : 1'h1; // @[d_cache.scala 282:35 295:26]
  wire [31:0] _GEN_539 = state == 3'h6 ? write_back_addr : _GEN_516; // @[d_cache.scala 282:35 296:26]
  wire  _GEN_540 = state == 3'h6 | _GEN_520; // @[d_cache.scala 282:35 297:27]
  wire [7:0] _GEN_541 = state == 3'h6 ? 8'hf : 8'h0; // @[d_cache.scala 282:35 298:25]
  wire [63:0] _GEN_544 = state == 3'h6 ? write_back_data[63:0] : _GEN_521; // @[d_cache.scala 282:35 301:25]
  wire [7:0] _GEN_545 = state == 3'h6 ? 8'hff : _GEN_522; // @[d_cache.scala 282:35 302:25]
  wire  _GEN_547 = state == 3'h6 | _GEN_524; // @[d_cache.scala 282:35 304:26]
  wire  _GEN_548 = state == 3'h6 | _T_41; // @[d_cache.scala 282:35 305:26]
  wire [63:0] _GEN_549 = state == 3'h4 ? 64'h0 : _GEN_526; // @[d_cache.scala 257:31 258:25]
  wire  _GEN_551 = state == 3'h4 ? 1'h0 : _GEN_528; // @[d_cache.scala 257:31 260:26]
  wire  _GEN_554 = state == 3'h4 ? io_from_axi_bvalid : _GEN_531; // @[d_cache.scala 257:31 263:26]
  wire  _GEN_556 = state == 3'h4 ? 1'h0 : _GEN_533; // @[d_cache.scala 257:31 265:27]
  wire [31:0] _GEN_557 = state == 3'h4 ? 32'h0 : _GEN_534; // @[d_cache.scala 257:31 266:26]
  wire  _GEN_561 = state == 3'h4 | _GEN_538; // @[d_cache.scala 257:31 270:26]
  wire [31:0] _GEN_562 = state == 3'h4 ? io_from_lsu_awaddr : _GEN_539; // @[d_cache.scala 257:31 271:26]
  wire  _GEN_563 = state == 3'h4 ? io_from_lsu_awvalid : _GEN_540; // @[d_cache.scala 257:31 272:27]
  wire [7:0] _GEN_564 = state == 3'h4 ? 8'h0 : _GEN_541; // @[d_cache.scala 257:31 273:25]
  wire [63:0] _GEN_567 = state == 3'h4 ? io_from_lsu_wdata : _GEN_544; // @[d_cache.scala 257:31 276:25]
  wire [7:0] _GEN_568 = state == 3'h4 ? io_from_lsu_wstrb : _GEN_545; // @[d_cache.scala 257:31 277:25]
  wire  _GEN_570 = state == 3'h4 ? io_from_lsu_wvalid : _GEN_547; // @[d_cache.scala 257:31 279:26]
  wire  _GEN_571 = state == 3'h4 | _GEN_548; // @[d_cache.scala 257:31 280:26]
  wire [63:0] _GEN_572 = state == 3'h3 ? 64'h0 : _GEN_549; // @[d_cache.scala 233:31 234:25]
  wire  _GEN_574 = state == 3'h3 ? 1'h0 : _GEN_551; // @[d_cache.scala 233:31 236:26]
  wire  _GEN_577 = state == 3'h3 ? 1'h0 : _GEN_554; // @[d_cache.scala 233:31 239:26]
  wire  _GEN_579 = state == 3'h3 | _GEN_556; // @[d_cache.scala 233:31 241:27]
  wire [63:0] _GEN_580 = state == 3'h3 ? _io_to_axi_araddr_T : {{32'd0}, _GEN_557}; // @[d_cache.scala 233:31 242:26]
  wire [7:0] _GEN_581 = state == 3'h3 ? 8'hf : 8'h0; // @[d_cache.scala 233:31 243:25]
  wire  _GEN_584 = state == 3'h3 | _GEN_561; // @[d_cache.scala 233:31 246:26]
  wire [31:0] _GEN_585 = state == 3'h3 ? 32'h0 : _GEN_562; // @[d_cache.scala 233:31 247:26]
  wire  _GEN_586 = state == 3'h3 ? 1'h0 : _GEN_563; // @[d_cache.scala 233:31 248:27]
  wire [7:0] _GEN_587 = state == 3'h3 ? 8'h0 : _GEN_564; // @[d_cache.scala 233:31 249:25]
  wire [63:0] _GEN_590 = state == 3'h3 ? 64'h0 : _GEN_567; // @[d_cache.scala 233:31 252:25]
  wire [7:0] _GEN_591 = state == 3'h3 ? 8'h0 : _GEN_568; // @[d_cache.scala 233:31 253:25]
  wire  _GEN_593 = state == 3'h3 ? 1'h0 : _GEN_570; // @[d_cache.scala 233:31 255:26]
  wire  _GEN_594 = state == 3'h3 ? 1'h0 : _GEN_571; // @[d_cache.scala 233:31 256:26]
  wire  _GEN_595 = state == 3'h2 ? 1'h0 : _GEN_579; // @[d_cache.scala 209:33 210:27]
  wire [63:0] _GEN_596 = state == 3'h2 ? {{32'd0}, io_from_lsu_araddr} : _GEN_580; // @[d_cache.scala 209:33 211:26]
  wire [7:0] _GEN_597 = state == 3'h2 ? 8'h0 : _GEN_581; // @[d_cache.scala 209:33 212:25]
  wire  _GEN_600 = state == 3'h2 ? 1'h0 : _GEN_584; // @[d_cache.scala 209:33 215:26]
  wire [31:0] _GEN_601 = state == 3'h2 ? 32'h0 : _GEN_585; // @[d_cache.scala 209:33 216:26]
  wire  _GEN_602 = state == 3'h2 ? 1'h0 : _GEN_586; // @[d_cache.scala 209:33 217:27]
  wire [7:0] _GEN_603 = state == 3'h2 ? 8'h0 : _GEN_587; // @[d_cache.scala 209:33 218:25]
  wire [63:0] _GEN_606 = state == 3'h2 ? 64'h0 : _GEN_590; // @[d_cache.scala 209:33 221:25]
  wire [7:0] _GEN_607 = state == 3'h2 ? 8'h0 : _GEN_591; // @[d_cache.scala 209:33 222:25]
  wire  _GEN_609 = state == 3'h2 ? 1'h0 : _GEN_593; // @[d_cache.scala 209:33 224:26]
  wire  _GEN_610 = state == 3'h2 ? 1'h0 : _GEN_594; // @[d_cache.scala 209:33 225:26]
  wire [63:0] _GEN_611 = state == 3'h2 ? 64'h0 : _GEN_572; // @[d_cache.scala 209:33 226:25]
  wire  _GEN_613 = state == 3'h2 ? 1'h0 : _GEN_574; // @[d_cache.scala 209:33 228:26]
  wire  _GEN_617 = state == 3'h2 ? anyMatch : _GEN_577; // @[d_cache.scala 209:33 232:26]
  wire [63:0] _GEN_619 = state == 3'h1 ? {{32'd0}, io_from_lsu_araddr} : _GEN_596; // @[d_cache.scala 184:27 186:26]
  wire [1023:0] _GEN_637 = state == 3'h1 ? _io_to_lsu_rdata_T_1 : {{960'd0}, _GEN_611}; // @[d_cache.scala 184:27 201:25]
  wire [42:0] _GEN_588 = reset ? 43'h0 : _GEN_499; // @[d_cache.scala 71:{34,34}]
  assign cacheLine_MPORT_1_en = _T ? 1'h0 : _GEN_373;
  assign cacheLine_MPORT_1_addr = tagIndex[5:0];
  assign cacheLine_MPORT_1_data = cacheLine[cacheLine_MPORT_1_addr]; // @[d_cache.scala 24:24]
  assign cacheLine_write_back_data_MPORT_en = _T ? 1'h0 : _GEN_429;
  assign cacheLine_write_back_data_MPORT_addr = replaceIndex[5:0];
  assign cacheLine_write_back_data_MPORT_data = cacheLine[cacheLine_write_back_data_MPORT_addr]; // @[d_cache.scala 24:24]
  assign cacheLine_io_to_lsu_rdata_MPORT_en = state == 3'h1;
  assign cacheLine_io_to_lsu_rdata_MPORT_addr = tagIndex[5:0];
  assign cacheLine_io_to_lsu_rdata_MPORT_data = cacheLine[cacheLine_io_to_lsu_rdata_MPORT_addr]; // @[d_cache.scala 24:24]
  assign cacheLine_MPORT_data = _T_13[1023:0];
  assign cacheLine_MPORT_addr = tagIndex[5:0];
  assign cacheLine_MPORT_mask = 1'h1;
  assign cacheLine_MPORT_en = _T ? 1'h0 : _GEN_373;
  assign cacheLine_MPORT_3_data = {hi,lo};
  assign cacheLine_MPORT_3_addr = unvalidIndex[5:0];
  assign cacheLine_MPORT_3_mask = 1'h1;
  assign cacheLine_MPORT_3_en = _T ? 1'h0 : _GEN_396;
  assign cacheLine_MPORT_6_data = {hi,lo};
  assign cacheLine_MPORT_6_addr = replaceIndex[5:0];
  assign cacheLine_MPORT_6_mask = 1'h1;
  assign cacheLine_MPORT_6_en = _T ? 1'h0 : _GEN_420;
  assign validMem_valid_0_MPORT_en = 1'h1;
  assign validMem_valid_0_MPORT_addr = _valid_0_T_1[5:0];
  assign validMem_valid_0_MPORT_data = validMem[validMem_valid_0_MPORT_addr]; // @[d_cache.scala 25:23]
  assign validMem_valid_1_MPORT_en = 1'h1;
  assign validMem_valid_1_MPORT_addr = _valid_1_T_2[5:0];
  assign validMem_valid_1_MPORT_data = validMem[validMem_valid_1_MPORT_addr]; // @[d_cache.scala 25:23]
  assign validMem_valid_2_MPORT_en = 1'h1;
  assign validMem_valid_2_MPORT_addr = _valid_2_T_2[5:0];
  assign validMem_valid_2_MPORT_data = validMem[validMem_valid_2_MPORT_addr]; // @[d_cache.scala 25:23]
  assign validMem_valid_3_MPORT_en = 1'h1;
  assign validMem_valid_3_MPORT_addr = _valid_3_T_2[5:0];
  assign validMem_valid_3_MPORT_data = validMem[validMem_valid_3_MPORT_addr]; // @[d_cache.scala 25:23]
  assign validMem_MPORT_5_data = 1'h1;
  assign validMem_MPORT_5_addr = unvalidIndex[5:0];
  assign validMem_MPORT_5_mask = 1'h1;
  assign validMem_MPORT_5_en = _T ? 1'h0 : _GEN_396;
  assign validMem_MPORT_8_data = 1'h1;
  assign validMem_MPORT_8_addr = replaceIndex[5:0];
  assign validMem_MPORT_8_mask = 1'h1;
  assign validMem_MPORT_8_en = _T ? 1'h0 : _GEN_420;
  assign tagMem_tagMatch_0_MPORT_en = 1'h1;
  assign tagMem_tagMatch_0_MPORT_addr = _valid_0_T_1[5:0];
  assign tagMem_tagMatch_0_MPORT_data = tagMem[tagMem_tagMatch_0_MPORT_addr]; // @[d_cache.scala 28:21]
  assign tagMem_tagMatch_1_MPORT_en = 1'h1;
  assign tagMem_tagMatch_1_MPORT_addr = _valid_1_T_2[5:0];
  assign tagMem_tagMatch_1_MPORT_data = tagMem[tagMem_tagMatch_1_MPORT_addr]; // @[d_cache.scala 28:21]
  assign tagMem_tagMatch_2_MPORT_en = 1'h1;
  assign tagMem_tagMatch_2_MPORT_addr = _valid_2_T_2[5:0];
  assign tagMem_tagMatch_2_MPORT_data = tagMem[tagMem_tagMatch_2_MPORT_addr]; // @[d_cache.scala 28:21]
  assign tagMem_tagMatch_3_MPORT_en = 1'h1;
  assign tagMem_tagMatch_3_MPORT_addr = _valid_3_T_2[5:0];
  assign tagMem_tagMatch_3_MPORT_data = tagMem[tagMem_tagMatch_3_MPORT_addr]; // @[d_cache.scala 28:21]
  assign tagMem_write_back_addr_MPORT_en = _T ? 1'h0 : _GEN_429;
  assign tagMem_write_back_addr_MPORT_addr = replaceIndex[5:0];
  assign tagMem_write_back_addr_MPORT_data = tagMem[tagMem_write_back_addr_MPORT_addr]; // @[d_cache.scala 28:21]
  assign tagMem_MPORT_4_data = {{11'd0}, tag};
  assign tagMem_MPORT_4_addr = unvalidIndex[5:0];
  assign tagMem_MPORT_4_mask = 1'h1;
  assign tagMem_MPORT_4_en = _T ? 1'h0 : _GEN_396;
  assign tagMem_MPORT_7_data = {{11'd0}, tag};
  assign tagMem_MPORT_7_addr = replaceIndex[5:0];
  assign tagMem_MPORT_7_mask = 1'h1;
  assign tagMem_MPORT_7_en = _T ? 1'h0 : _GEN_420;
  assign dirtyMem_MPORT_9_en = _T ? 1'h0 : _GEN_420;
  assign dirtyMem_MPORT_9_addr = replaceIndex[5:0];
  assign dirtyMem_MPORT_9_data = dirtyMem[dirtyMem_MPORT_9_addr]; // @[d_cache.scala 29:23]
  assign dirtyMem_MPORT_2_data = 1'h1;
  assign dirtyMem_MPORT_2_addr = tagIndex[5:0];
  assign dirtyMem_MPORT_2_mask = 1'h1;
  assign dirtyMem_MPORT_2_en = _T ? 1'h0 : _GEN_373;
  assign dirtyMem_MPORT_10_data = 1'h0;
  assign dirtyMem_MPORT_10_addr = replaceIndex[5:0];
  assign dirtyMem_MPORT_10_mask = 1'h1;
  assign dirtyMem_MPORT_10_en = _T ? 1'h0 : _GEN_429;
  assign io_to_lsu_rdata = _GEN_637[63:0];
  assign io_to_lsu_rvalid = state == 3'h1 ? anyMatch : _GEN_613; // @[d_cache.scala 184:27 203:26]
  assign io_to_lsu_bvalid = state == 3'h1 ? 1'h0 : _GEN_617; // @[d_cache.scala 184:27 207:26]
  assign io_to_axi_araddr = _GEN_619[31:0];
  assign io_to_axi_arlen = state == 3'h1 ? 8'h0 : _GEN_597; // @[d_cache.scala 184:27 187:25]
  assign io_to_axi_arvalid = state == 3'h1 ? 1'h0 : _GEN_595; // @[d_cache.scala 184:27 185:27]
  assign io_to_axi_rready = state == 3'h1 ? 1'h0 : _GEN_600; // @[d_cache.scala 184:27 190:26]
  assign io_to_axi_awaddr = state == 3'h1 ? 32'h0 : _GEN_601; // @[d_cache.scala 184:27 191:26]
  assign io_to_axi_awlen = state == 3'h1 ? 8'h0 : _GEN_603; // @[d_cache.scala 184:27 193:25]
  assign io_to_axi_awvalid = state == 3'h1 ? 1'h0 : _GEN_602; // @[d_cache.scala 184:27 192:27]
  assign io_to_axi_wdata = state == 3'h1 ? 64'h0 : _GEN_606; // @[d_cache.scala 184:27 196:25]
  assign io_to_axi_wstrb = state == 3'h1 ? 8'h0 : _GEN_607; // @[d_cache.scala 184:27 197:25]
  assign io_to_axi_wvalid = state == 3'h1 ? 1'h0 : _GEN_609; // @[d_cache.scala 184:27 199:26]
  assign io_to_axi_bready = state == 3'h1 ? 1'h0 : _GEN_610; // @[d_cache.scala 184:27 200:26]
  always @(posedge clock) begin
    if (cacheLine_MPORT_en & cacheLine_MPORT_mask) begin
      cacheLine[cacheLine_MPORT_addr] <= cacheLine_MPORT_data; // @[d_cache.scala 24:24]
    end
    if (cacheLine_MPORT_3_en & cacheLine_MPORT_3_mask) begin
      cacheLine[cacheLine_MPORT_3_addr] <= cacheLine_MPORT_3_data; // @[d_cache.scala 24:24]
    end
    if (cacheLine_MPORT_6_en & cacheLine_MPORT_6_mask) begin
      cacheLine[cacheLine_MPORT_6_addr] <= cacheLine_MPORT_6_data; // @[d_cache.scala 24:24]
    end
    if (validMem_MPORT_5_en & validMem_MPORT_5_mask) begin
      validMem[validMem_MPORT_5_addr] <= validMem_MPORT_5_data; // @[d_cache.scala 25:23]
    end
    if (validMem_MPORT_8_en & validMem_MPORT_8_mask) begin
      validMem[validMem_MPORT_8_addr] <= validMem_MPORT_8_data; // @[d_cache.scala 25:23]
    end
    if (tagMem_MPORT_4_en & tagMem_MPORT_4_mask) begin
      tagMem[tagMem_MPORT_4_addr] <= tagMem_MPORT_4_data; // @[d_cache.scala 28:21]
    end
    if (tagMem_MPORT_7_en & tagMem_MPORT_7_mask) begin
      tagMem[tagMem_MPORT_7_addr] <= tagMem_MPORT_7_data; // @[d_cache.scala 28:21]
    end
    if (dirtyMem_MPORT_2_en & dirtyMem_MPORT_2_mask) begin
      dirtyMem[dirtyMem_MPORT_2_addr] <= dirtyMem_MPORT_2_data; // @[d_cache.scala 29:23]
    end
    if (dirtyMem_MPORT_10_en & dirtyMem_MPORT_10_mask) begin
      dirtyMem[dirtyMem_MPORT_10_addr] <= dirtyMem_MPORT_10_data; // @[d_cache.scala 29:23]
    end
    if (reset) begin // @[d_cache.scala 70:34]
      write_back_data <= 1024'h0; // @[d_cache.scala 70:34]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          write_back_data <= _GEN_296;
        end
      end
    end
    write_back_addr <= _GEN_588[31:0]; // @[d_cache.scala 71:{34,34}]
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_0 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_0 <= _GEN_242;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_1 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_1 <= _GEN_243;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_2 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_2 <= _GEN_244;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_3 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_3 <= _GEN_245;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_4 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_4 <= _GEN_246;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_5 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_5 <= _GEN_247;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_6 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_6 <= _GEN_248;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_7 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_7 <= _GEN_249;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_8 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_8 <= _GEN_250;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_9 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_9 <= _GEN_251;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_10 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_10 <= _GEN_252;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_11 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_11 <= _GEN_253;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_12 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_12 <= _GEN_254;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_13 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_13 <= _GEN_255;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_14 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_14 <= _GEN_256;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 75:31]
      receive_data_15 <= 64'h0; // @[d_cache.scala 75:31]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          receive_data_15 <= _GEN_257;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 76:30]
      receive_num <= 3'h0; // @[d_cache.scala 76:30]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (3'h1 == state) begin // @[d_cache.scala 101:18]
        if (!(anyMatch)) begin // @[d_cache.scala 112:27]
          receive_num <= 3'h0; // @[d_cache.scala 118:29]
        end
      end else if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
        receive_num <= _GEN_258;
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_0 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_0 <= _GEN_268;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_1 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_1 <= _GEN_269;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_2 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_2 <= _GEN_270;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_3 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_3 <= _GEN_271;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_4 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_4 <= _GEN_272;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_5 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_5 <= _GEN_273;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_6 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_6 <= _GEN_274;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_7 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_7 <= _GEN_275;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_8 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_8 <= _GEN_276;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_9 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_9 <= _GEN_277;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_10 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_10 <= _GEN_278;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_11 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_11 <= _GEN_279;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_12 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_12 <= _GEN_280;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_13 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_13 <= _GEN_281;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_14 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_14 <= _GEN_282;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 77:24]
      quene_15 <= 8'h0; // @[d_cache.scala 77:24]
    end else if (!(3'h0 == state)) begin // @[d_cache.scala 101:18]
      if (!(3'h1 == state)) begin // @[d_cache.scala 101:18]
        if (!(3'h2 == state)) begin // @[d_cache.scala 101:18]
          quene_15 <= _GEN_283;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 95:24]
      state <= 3'h0; // @[d_cache.scala 95:24]
    end else if (3'h0 == state) begin // @[d_cache.scala 101:18]
      if ((io_from_lsu_arvalid | io_from_lsu_awvalid) & io_from_lsu_araddr >= 32'ha0000000) begin // @[d_cache.scala 103:99]
        state <= 3'h0; // @[d_cache.scala 104:23]
      end else if (io_from_lsu_arvalid) begin // @[d_cache.scala 105:44]
        state <= 3'h1; // @[d_cache.scala 106:23]
      end else begin
        state <= _GEN_16;
      end
    end else if (3'h1 == state) begin // @[d_cache.scala 101:18]
      if (anyMatch) begin // @[d_cache.scala 112:27]
        state <= 3'h0;
      end else begin
        state <= 3'h3; // @[d_cache.scala 117:23]
      end
    end else if (3'h2 == state) begin // @[d_cache.scala 101:18]
      state <= _GEN_23;
    end else begin
      state <= _GEN_259;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {32{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    cacheLine[initvar] = _RAND_0[1023:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    validMem[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tagMem[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    dirtyMem[initvar] = _RAND_3[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {32{`RANDOM}};
  write_back_data = _RAND_4[1023:0];
  _RAND_5 = {1{`RANDOM}};
  write_back_addr = _RAND_5[31:0];
  _RAND_6 = {2{`RANDOM}};
  receive_data_0 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  receive_data_1 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  receive_data_2 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  receive_data_3 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  receive_data_4 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  receive_data_5 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  receive_data_6 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  receive_data_7 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  receive_data_8 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  receive_data_9 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  receive_data_10 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  receive_data_11 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  receive_data_12 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  receive_data_13 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  receive_data_14 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  receive_data_15 = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  receive_num = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  quene_0 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  quene_1 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  quene_2 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  quene_3 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  quene_4 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  quene_5 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  quene_6 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  quene_7 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  quene_8 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  quene_9 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  quene_10 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  quene_11 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  quene_12 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  quene_13 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  quene_14 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  quene_15 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  state = _RAND_39[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
