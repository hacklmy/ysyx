module D_CACHE(
  input         clock,
  input         reset,
  input  [31:0] io_from_lsu_araddr,
  input         io_from_lsu_arvalid,
  input  [31:0] io_from_lsu_awaddr,
  input         io_from_lsu_awvalid,
  input  [63:0] io_from_lsu_wdata,
  input  [7:0]  io_from_lsu_wstrb,
  input         io_from_lsu_wvalid,
  output [63:0] io_to_lsu_rdata,
  output        io_to_lsu_rvalid,
  output        io_to_lsu_wready,
  output [31:0] io_to_axi_araddr,
  output [7:0]  io_to_axi_arlen,
  output        io_to_axi_arvalid,
  output        io_to_axi_rready,
  output [31:0] io_to_axi_awaddr,
  output [7:0]  io_to_axi_awlen,
  output        io_to_axi_awvalid,
  output [63:0] io_to_axi_wdata,
  output [7:0]  io_to_axi_wstrb,
  output        io_to_axi_wvalid,
  output        io_to_axi_bready,
  input  [63:0] io_from_axi_rdata,
  input         io_from_axi_rlast,
  input         io_from_axi_rvalid,
  input         io_from_axi_wready,
  input         io_from_axi_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [511:0] _RAND_2;
  reg [511:0] _RAND_3;
  reg [511:0] _RAND_4;
  reg [511:0] _RAND_5;
  reg [511:0] _RAND_6;
  reg [511:0] _RAND_7;
  reg [511:0] _RAND_8;
  reg [511:0] _RAND_9;
  reg [511:0] _RAND_10;
  reg [511:0] _RAND_11;
  reg [511:0] _RAND_12;
  reg [511:0] _RAND_13;
  reg [511:0] _RAND_14;
  reg [511:0] _RAND_15;
  reg [511:0] _RAND_16;
  reg [511:0] _RAND_17;
  reg [511:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [511:0] _RAND_21;
  reg [511:0] _RAND_22;
  reg [511:0] _RAND_23;
  reg [511:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [511:0] _RAND_26;
  reg [511:0] _RAND_27;
  reg [511:0] _RAND_28;
  reg [511:0] _RAND_29;
  reg [511:0] _RAND_30;
  reg [511:0] _RAND_31;
  reg [511:0] _RAND_32;
  reg [511:0] _RAND_33;
  reg [511:0] _RAND_34;
  reg [511:0] _RAND_35;
  reg [511:0] _RAND_36;
  reg [511:0] _RAND_37;
  reg [511:0] _RAND_38;
  reg [511:0] _RAND_39;
  reg [511:0] _RAND_40;
  reg [511:0] _RAND_41;
  reg [511:0] _RAND_42;
  reg [511:0] _RAND_43;
  reg [511:0] _RAND_44;
  reg [511:0] _RAND_45;
  reg [511:0] _RAND_46;
  reg [511:0] _RAND_47;
  reg [511:0] _RAND_48;
  reg [511:0] _RAND_49;
  reg [511:0] _RAND_50;
  reg [511:0] _RAND_51;
  reg [511:0] _RAND_52;
  reg [511:0] _RAND_53;
  reg [511:0] _RAND_54;
  reg [511:0] _RAND_55;
  reg [511:0] _RAND_56;
  reg [511:0] _RAND_57;
  reg [511:0] _RAND_58;
  reg [511:0] _RAND_59;
  reg [511:0] _RAND_60;
  reg [511:0] _RAND_61;
  reg [511:0] _RAND_62;
  reg [511:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [511:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [63:0] _RAND_258;
  reg [63:0] _RAND_259;
  reg [63:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [63:0] _RAND_263;
  reg [63:0] _RAND_264;
  reg [63:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] ram_0_0; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_1; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_2; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_3; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_4; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_5; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_6; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_7; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_8; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_9; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_10; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_11; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_12; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_13; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_14; // @[d_cache.scala 19:24]
  reg [511:0] ram_0_15; // @[d_cache.scala 19:24]
  reg [511:0] ram_1_0; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_1; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_2; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_3; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_4; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_5; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_6; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_7; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_8; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_9; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_10; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_11; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_12; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_13; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_14; // @[d_cache.scala 20:24]
  reg [511:0] ram_1_15; // @[d_cache.scala 20:24]
  reg [511:0] ram_2_0; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_1; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_2; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_3; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_4; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_5; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_6; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_7; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_8; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_9; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_10; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_11; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_12; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_13; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_14; // @[d_cache.scala 21:24]
  reg [511:0] ram_2_15; // @[d_cache.scala 21:24]
  reg [511:0] ram_3_0; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_1; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_2; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_3; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_4; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_5; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_6; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_7; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_8; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_9; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_10; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_11; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_12; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_13; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_14; // @[d_cache.scala 22:24]
  reg [511:0] ram_3_15; // @[d_cache.scala 22:24]
  reg [31:0] tag_0_0; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_1; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_2; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_3; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_4; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_5; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_6; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_7; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_8; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_9; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_10; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_11; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_12; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_13; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_14; // @[d_cache.scala 24:24]
  reg [31:0] tag_0_15; // @[d_cache.scala 24:24]
  reg [31:0] tag_1_0; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_1; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_2; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_3; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_4; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_5; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_6; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_7; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_8; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_9; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_10; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_11; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_12; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_13; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_14; // @[d_cache.scala 25:24]
  reg [31:0] tag_1_15; // @[d_cache.scala 25:24]
  reg [31:0] tag_2_0; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_1; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_2; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_3; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_4; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_5; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_6; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_7; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_8; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_9; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_10; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_11; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_12; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_13; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_14; // @[d_cache.scala 26:24]
  reg [31:0] tag_2_15; // @[d_cache.scala 26:24]
  reg [31:0] tag_3_0; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_1; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_2; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_3; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_4; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_5; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_6; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_7; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_8; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_9; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_10; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_11; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_12; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_13; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_14; // @[d_cache.scala 27:24]
  reg [31:0] tag_3_15; // @[d_cache.scala 27:24]
  reg  valid_0_0; // @[d_cache.scala 29:26]
  reg  valid_0_1; // @[d_cache.scala 29:26]
  reg  valid_0_2; // @[d_cache.scala 29:26]
  reg  valid_0_3; // @[d_cache.scala 29:26]
  reg  valid_0_4; // @[d_cache.scala 29:26]
  reg  valid_0_5; // @[d_cache.scala 29:26]
  reg  valid_0_6; // @[d_cache.scala 29:26]
  reg  valid_0_7; // @[d_cache.scala 29:26]
  reg  valid_0_8; // @[d_cache.scala 29:26]
  reg  valid_0_9; // @[d_cache.scala 29:26]
  reg  valid_0_10; // @[d_cache.scala 29:26]
  reg  valid_0_11; // @[d_cache.scala 29:26]
  reg  valid_0_12; // @[d_cache.scala 29:26]
  reg  valid_0_13; // @[d_cache.scala 29:26]
  reg  valid_0_14; // @[d_cache.scala 29:26]
  reg  valid_0_15; // @[d_cache.scala 29:26]
  reg  valid_1_0; // @[d_cache.scala 30:26]
  reg  valid_1_1; // @[d_cache.scala 30:26]
  reg  valid_1_2; // @[d_cache.scala 30:26]
  reg  valid_1_3; // @[d_cache.scala 30:26]
  reg  valid_1_4; // @[d_cache.scala 30:26]
  reg  valid_1_5; // @[d_cache.scala 30:26]
  reg  valid_1_6; // @[d_cache.scala 30:26]
  reg  valid_1_7; // @[d_cache.scala 30:26]
  reg  valid_1_8; // @[d_cache.scala 30:26]
  reg  valid_1_9; // @[d_cache.scala 30:26]
  reg  valid_1_10; // @[d_cache.scala 30:26]
  reg  valid_1_11; // @[d_cache.scala 30:26]
  reg  valid_1_12; // @[d_cache.scala 30:26]
  reg  valid_1_13; // @[d_cache.scala 30:26]
  reg  valid_1_14; // @[d_cache.scala 30:26]
  reg  valid_1_15; // @[d_cache.scala 30:26]
  reg  valid_2_0; // @[d_cache.scala 31:26]
  reg  valid_2_1; // @[d_cache.scala 31:26]
  reg  valid_2_2; // @[d_cache.scala 31:26]
  reg  valid_2_3; // @[d_cache.scala 31:26]
  reg  valid_2_4; // @[d_cache.scala 31:26]
  reg  valid_2_5; // @[d_cache.scala 31:26]
  reg  valid_2_6; // @[d_cache.scala 31:26]
  reg  valid_2_7; // @[d_cache.scala 31:26]
  reg  valid_2_8; // @[d_cache.scala 31:26]
  reg  valid_2_9; // @[d_cache.scala 31:26]
  reg  valid_2_10; // @[d_cache.scala 31:26]
  reg  valid_2_11; // @[d_cache.scala 31:26]
  reg  valid_2_12; // @[d_cache.scala 31:26]
  reg  valid_2_13; // @[d_cache.scala 31:26]
  reg  valid_2_14; // @[d_cache.scala 31:26]
  reg  valid_2_15; // @[d_cache.scala 31:26]
  reg  valid_3_0; // @[d_cache.scala 32:26]
  reg  valid_3_1; // @[d_cache.scala 32:26]
  reg  valid_3_2; // @[d_cache.scala 32:26]
  reg  valid_3_3; // @[d_cache.scala 32:26]
  reg  valid_3_4; // @[d_cache.scala 32:26]
  reg  valid_3_5; // @[d_cache.scala 32:26]
  reg  valid_3_6; // @[d_cache.scala 32:26]
  reg  valid_3_7; // @[d_cache.scala 32:26]
  reg  valid_3_8; // @[d_cache.scala 32:26]
  reg  valid_3_9; // @[d_cache.scala 32:26]
  reg  valid_3_10; // @[d_cache.scala 32:26]
  reg  valid_3_11; // @[d_cache.scala 32:26]
  reg  valid_3_12; // @[d_cache.scala 32:26]
  reg  valid_3_13; // @[d_cache.scala 32:26]
  reg  valid_3_14; // @[d_cache.scala 32:26]
  reg  valid_3_15; // @[d_cache.scala 32:26]
  reg  dirty_0_0; // @[d_cache.scala 34:26]
  reg  dirty_0_1; // @[d_cache.scala 34:26]
  reg  dirty_0_2; // @[d_cache.scala 34:26]
  reg  dirty_0_3; // @[d_cache.scala 34:26]
  reg  dirty_0_4; // @[d_cache.scala 34:26]
  reg  dirty_0_5; // @[d_cache.scala 34:26]
  reg  dirty_0_6; // @[d_cache.scala 34:26]
  reg  dirty_0_7; // @[d_cache.scala 34:26]
  reg  dirty_0_8; // @[d_cache.scala 34:26]
  reg  dirty_0_9; // @[d_cache.scala 34:26]
  reg  dirty_0_10; // @[d_cache.scala 34:26]
  reg  dirty_0_11; // @[d_cache.scala 34:26]
  reg  dirty_0_12; // @[d_cache.scala 34:26]
  reg  dirty_0_13; // @[d_cache.scala 34:26]
  reg  dirty_0_14; // @[d_cache.scala 34:26]
  reg  dirty_0_15; // @[d_cache.scala 34:26]
  reg  dirty_1_0; // @[d_cache.scala 35:26]
  reg  dirty_1_1; // @[d_cache.scala 35:26]
  reg  dirty_1_2; // @[d_cache.scala 35:26]
  reg  dirty_1_3; // @[d_cache.scala 35:26]
  reg  dirty_1_4; // @[d_cache.scala 35:26]
  reg  dirty_1_5; // @[d_cache.scala 35:26]
  reg  dirty_1_6; // @[d_cache.scala 35:26]
  reg  dirty_1_7; // @[d_cache.scala 35:26]
  reg  dirty_1_8; // @[d_cache.scala 35:26]
  reg  dirty_1_9; // @[d_cache.scala 35:26]
  reg  dirty_1_10; // @[d_cache.scala 35:26]
  reg  dirty_1_11; // @[d_cache.scala 35:26]
  reg  dirty_1_12; // @[d_cache.scala 35:26]
  reg  dirty_1_13; // @[d_cache.scala 35:26]
  reg  dirty_1_14; // @[d_cache.scala 35:26]
  reg  dirty_1_15; // @[d_cache.scala 35:26]
  reg  dirty_2_0; // @[d_cache.scala 36:26]
  reg  dirty_2_1; // @[d_cache.scala 36:26]
  reg  dirty_2_2; // @[d_cache.scala 36:26]
  reg  dirty_2_3; // @[d_cache.scala 36:26]
  reg  dirty_2_4; // @[d_cache.scala 36:26]
  reg  dirty_2_5; // @[d_cache.scala 36:26]
  reg  dirty_2_6; // @[d_cache.scala 36:26]
  reg  dirty_2_7; // @[d_cache.scala 36:26]
  reg  dirty_2_8; // @[d_cache.scala 36:26]
  reg  dirty_2_9; // @[d_cache.scala 36:26]
  reg  dirty_2_10; // @[d_cache.scala 36:26]
  reg  dirty_2_11; // @[d_cache.scala 36:26]
  reg  dirty_2_12; // @[d_cache.scala 36:26]
  reg  dirty_2_13; // @[d_cache.scala 36:26]
  reg  dirty_2_14; // @[d_cache.scala 36:26]
  reg  dirty_2_15; // @[d_cache.scala 36:26]
  reg  dirty_3_0; // @[d_cache.scala 37:26]
  reg  dirty_3_1; // @[d_cache.scala 37:26]
  reg  dirty_3_2; // @[d_cache.scala 37:26]
  reg  dirty_3_3; // @[d_cache.scala 37:26]
  reg  dirty_3_4; // @[d_cache.scala 37:26]
  reg  dirty_3_5; // @[d_cache.scala 37:26]
  reg  dirty_3_6; // @[d_cache.scala 37:26]
  reg  dirty_3_7; // @[d_cache.scala 37:26]
  reg  dirty_3_8; // @[d_cache.scala 37:26]
  reg  dirty_3_9; // @[d_cache.scala 37:26]
  reg  dirty_3_10; // @[d_cache.scala 37:26]
  reg  dirty_3_11; // @[d_cache.scala 37:26]
  reg  dirty_3_12; // @[d_cache.scala 37:26]
  reg  dirty_3_13; // @[d_cache.scala 37:26]
  reg  dirty_3_14; // @[d_cache.scala 37:26]
  reg  dirty_3_15; // @[d_cache.scala 37:26]
  reg [511:0] write_back_data; // @[d_cache.scala 44:34]
  reg [31:0] write_back_addr; // @[d_cache.scala 45:34]
  reg [63:0] receive_data_0; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_1; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_2; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_3; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_4; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_5; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_6; // @[d_cache.scala 50:31]
  reg [63:0] receive_data_7; // @[d_cache.scala 50:31]
  reg [2:0] receive_num; // @[d_cache.scala 51:30]
  reg [7:0] quene_0; // @[d_cache.scala 52:24]
  reg [7:0] quene_1; // @[d_cache.scala 52:24]
  reg [7:0] quene_2; // @[d_cache.scala 52:24]
  reg [7:0] quene_3; // @[d_cache.scala 52:24]
  reg [7:0] quene_4; // @[d_cache.scala 52:24]
  reg [7:0] quene_5; // @[d_cache.scala 52:24]
  reg [7:0] quene_6; // @[d_cache.scala 52:24]
  reg [7:0] quene_7; // @[d_cache.scala 52:24]
  reg [7:0] quene_8; // @[d_cache.scala 52:24]
  reg [7:0] quene_9; // @[d_cache.scala 52:24]
  reg [7:0] quene_10; // @[d_cache.scala 52:24]
  reg [7:0] quene_11; // @[d_cache.scala 52:24]
  reg [7:0] quene_12; // @[d_cache.scala 52:24]
  reg [7:0] quene_13; // @[d_cache.scala 52:24]
  reg [7:0] quene_14; // @[d_cache.scala 52:24]
  reg [7:0] quene_15; // @[d_cache.scala 52:24]
  wire [5:0] offset = io_from_lsu_araddr[5:0]; // @[d_cache.scala 54:36]
  wire [3:0] index = io_from_lsu_araddr[9:6]; // @[d_cache.scala 55:35]
  wire [21:0] tag = io_from_lsu_araddr[31:10]; // @[d_cache.scala 56:33]
  wire [8:0] shift_bit = {offset, 3'h0}; // @[d_cache.scala 58:28]
  wire [63:0] _wmask_T_4 = io_from_lsu_wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[d_cache.scala 71:20]
  wire [63:0] _wmask_T_5 = io_from_lsu_wstrb == 8'hf ? 64'hffffffff : _wmask_T_4; // @[d_cache.scala 70:20]
  wire [63:0] _wmask_T_6 = io_from_lsu_wstrb == 8'h3 ? 64'hffff : _wmask_T_5; // @[d_cache.scala 69:20]
  wire [63:0] wmask = io_from_lsu_wstrb == 8'h1 ? 64'hff : _wmask_T_6; // @[d_cache.scala 68:20]
  wire [31:0] _GEN_1 = 4'h1 == index ? tag_0_1 : tag_0_0; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_2 = 4'h2 == index ? tag_0_2 : _GEN_1; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_3 = 4'h3 == index ? tag_0_3 : _GEN_2; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_4 = 4'h4 == index ? tag_0_4 : _GEN_3; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_5 = 4'h5 == index ? tag_0_5 : _GEN_4; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_6 = 4'h6 == index ? tag_0_6 : _GEN_5; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_7 = 4'h7 == index ? tag_0_7 : _GEN_6; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_8 = 4'h8 == index ? tag_0_8 : _GEN_7; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_9 = 4'h9 == index ? tag_0_9 : _GEN_8; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_10 = 4'ha == index ? tag_0_10 : _GEN_9; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_11 = 4'hb == index ? tag_0_11 : _GEN_10; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_12 = 4'hc == index ? tag_0_12 : _GEN_11; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_13 = 4'hd == index ? tag_0_13 : _GEN_12; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_14 = 4'he == index ? tag_0_14 : _GEN_13; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_15 = 4'hf == index ? tag_0_15 : _GEN_14; // @[d_cache.scala 91:{31,31}]
  wire [31:0] _GEN_5341 = {{10'd0}, tag}; // @[d_cache.scala 91:31]
  wire  _GEN_17 = 4'h1 == index ? valid_0_1 : valid_0_0; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_18 = 4'h2 == index ? valid_0_2 : _GEN_17; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_19 = 4'h3 == index ? valid_0_3 : _GEN_18; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_20 = 4'h4 == index ? valid_0_4 : _GEN_19; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_21 = 4'h5 == index ? valid_0_5 : _GEN_20; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_22 = 4'h6 == index ? valid_0_6 : _GEN_21; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_23 = 4'h7 == index ? valid_0_7 : _GEN_22; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_24 = 4'h8 == index ? valid_0_8 : _GEN_23; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_25 = 4'h9 == index ? valid_0_9 : _GEN_24; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_26 = 4'ha == index ? valid_0_10 : _GEN_25; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_27 = 4'hb == index ? valid_0_11 : _GEN_26; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_28 = 4'hc == index ? valid_0_12 : _GEN_27; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_29 = 4'hd == index ? valid_0_13 : _GEN_28; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_30 = 4'he == index ? valid_0_14 : _GEN_29; // @[d_cache.scala 91:{57,57}]
  wire  _GEN_31 = 4'hf == index ? valid_0_15 : _GEN_30; // @[d_cache.scala 91:{57,57}]
  wire  way0_hit = _GEN_15 == _GEN_5341 & _GEN_31; // @[d_cache.scala 91:40]
  wire [31:0] _GEN_33 = 4'h1 == index ? tag_1_1 : tag_1_0; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_34 = 4'h2 == index ? tag_1_2 : _GEN_33; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_35 = 4'h3 == index ? tag_1_3 : _GEN_34; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_36 = 4'h4 == index ? tag_1_4 : _GEN_35; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_37 = 4'h5 == index ? tag_1_5 : _GEN_36; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_38 = 4'h6 == index ? tag_1_6 : _GEN_37; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_39 = 4'h7 == index ? tag_1_7 : _GEN_38; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_40 = 4'h8 == index ? tag_1_8 : _GEN_39; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_41 = 4'h9 == index ? tag_1_9 : _GEN_40; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_42 = 4'ha == index ? tag_1_10 : _GEN_41; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_43 = 4'hb == index ? tag_1_11 : _GEN_42; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_44 = 4'hc == index ? tag_1_12 : _GEN_43; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_45 = 4'hd == index ? tag_1_13 : _GEN_44; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_46 = 4'he == index ? tag_1_14 : _GEN_45; // @[d_cache.scala 93:{31,31}]
  wire [31:0] _GEN_47 = 4'hf == index ? tag_1_15 : _GEN_46; // @[d_cache.scala 93:{31,31}]
  wire  _GEN_49 = 4'h1 == index ? valid_1_1 : valid_1_0; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_50 = 4'h2 == index ? valid_1_2 : _GEN_49; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_51 = 4'h3 == index ? valid_1_3 : _GEN_50; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_52 = 4'h4 == index ? valid_1_4 : _GEN_51; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_53 = 4'h5 == index ? valid_1_5 : _GEN_52; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_54 = 4'h6 == index ? valid_1_6 : _GEN_53; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_55 = 4'h7 == index ? valid_1_7 : _GEN_54; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_56 = 4'h8 == index ? valid_1_8 : _GEN_55; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_57 = 4'h9 == index ? valid_1_9 : _GEN_56; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_58 = 4'ha == index ? valid_1_10 : _GEN_57; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_59 = 4'hb == index ? valid_1_11 : _GEN_58; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_60 = 4'hc == index ? valid_1_12 : _GEN_59; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_61 = 4'hd == index ? valid_1_13 : _GEN_60; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_62 = 4'he == index ? valid_1_14 : _GEN_61; // @[d_cache.scala 93:{57,57}]
  wire  _GEN_63 = 4'hf == index ? valid_1_15 : _GEN_62; // @[d_cache.scala 93:{57,57}]
  wire  way1_hit = _GEN_47 == _GEN_5341 & _GEN_63; // @[d_cache.scala 93:40]
  wire [31:0] _GEN_65 = 4'h1 == index ? tag_2_1 : tag_2_0; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_66 = 4'h2 == index ? tag_2_2 : _GEN_65; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_67 = 4'h3 == index ? tag_2_3 : _GEN_66; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_68 = 4'h4 == index ? tag_2_4 : _GEN_67; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_69 = 4'h5 == index ? tag_2_5 : _GEN_68; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_70 = 4'h6 == index ? tag_2_6 : _GEN_69; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_71 = 4'h7 == index ? tag_2_7 : _GEN_70; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_72 = 4'h8 == index ? tag_2_8 : _GEN_71; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_73 = 4'h9 == index ? tag_2_9 : _GEN_72; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_74 = 4'ha == index ? tag_2_10 : _GEN_73; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_75 = 4'hb == index ? tag_2_11 : _GEN_74; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_76 = 4'hc == index ? tag_2_12 : _GEN_75; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_77 = 4'hd == index ? tag_2_13 : _GEN_76; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_78 = 4'he == index ? tag_2_14 : _GEN_77; // @[d_cache.scala 94:{31,31}]
  wire [31:0] _GEN_79 = 4'hf == index ? tag_2_15 : _GEN_78; // @[d_cache.scala 94:{31,31}]
  wire  _GEN_81 = 4'h1 == index ? valid_2_1 : valid_2_0; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_82 = 4'h2 == index ? valid_2_2 : _GEN_81; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_83 = 4'h3 == index ? valid_2_3 : _GEN_82; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_84 = 4'h4 == index ? valid_2_4 : _GEN_83; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_85 = 4'h5 == index ? valid_2_5 : _GEN_84; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_86 = 4'h6 == index ? valid_2_6 : _GEN_85; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_87 = 4'h7 == index ? valid_2_7 : _GEN_86; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_88 = 4'h8 == index ? valid_2_8 : _GEN_87; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_89 = 4'h9 == index ? valid_2_9 : _GEN_88; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_90 = 4'ha == index ? valid_2_10 : _GEN_89; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_91 = 4'hb == index ? valid_2_11 : _GEN_90; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_92 = 4'hc == index ? valid_2_12 : _GEN_91; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_93 = 4'hd == index ? valid_2_13 : _GEN_92; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_94 = 4'he == index ? valid_2_14 : _GEN_93; // @[d_cache.scala 94:{57,57}]
  wire  _GEN_95 = 4'hf == index ? valid_2_15 : _GEN_94; // @[d_cache.scala 94:{57,57}]
  wire  way2_hit = _GEN_79 == _GEN_5341 & _GEN_95; // @[d_cache.scala 94:40]
  wire [31:0] _GEN_97 = 4'h1 == index ? tag_3_1 : tag_3_0; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_98 = 4'h2 == index ? tag_3_2 : _GEN_97; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_99 = 4'h3 == index ? tag_3_3 : _GEN_98; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_100 = 4'h4 == index ? tag_3_4 : _GEN_99; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_101 = 4'h5 == index ? tag_3_5 : _GEN_100; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_102 = 4'h6 == index ? tag_3_6 : _GEN_101; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_103 = 4'h7 == index ? tag_3_7 : _GEN_102; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_104 = 4'h8 == index ? tag_3_8 : _GEN_103; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_105 = 4'h9 == index ? tag_3_9 : _GEN_104; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_106 = 4'ha == index ? tag_3_10 : _GEN_105; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_107 = 4'hb == index ? tag_3_11 : _GEN_106; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_108 = 4'hc == index ? tag_3_12 : _GEN_107; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_109 = 4'hd == index ? tag_3_13 : _GEN_108; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_110 = 4'he == index ? tag_3_14 : _GEN_109; // @[d_cache.scala 95:{31,31}]
  wire [31:0] _GEN_111 = 4'hf == index ? tag_3_15 : _GEN_110; // @[d_cache.scala 95:{31,31}]
  wire  _GEN_113 = 4'h1 == index ? valid_3_1 : valid_3_0; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_114 = 4'h2 == index ? valid_3_2 : _GEN_113; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_115 = 4'h3 == index ? valid_3_3 : _GEN_114; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_116 = 4'h4 == index ? valid_3_4 : _GEN_115; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_117 = 4'h5 == index ? valid_3_5 : _GEN_116; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_118 = 4'h6 == index ? valid_3_6 : _GEN_117; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_119 = 4'h7 == index ? valid_3_7 : _GEN_118; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_120 = 4'h8 == index ? valid_3_8 : _GEN_119; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_121 = 4'h9 == index ? valid_3_9 : _GEN_120; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_122 = 4'ha == index ? valid_3_10 : _GEN_121; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_123 = 4'hb == index ? valid_3_11 : _GEN_122; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_124 = 4'hc == index ? valid_3_12 : _GEN_123; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_125 = 4'hd == index ? valid_3_13 : _GEN_124; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_126 = 4'he == index ? valid_3_14 : _GEN_125; // @[d_cache.scala 95:{57,57}]
  wire  _GEN_127 = 4'hf == index ? valid_3_15 : _GEN_126; // @[d_cache.scala 95:{57,57}]
  wire  way3_hit = _GEN_111 == _GEN_5341 & _GEN_127; // @[d_cache.scala 95:40]
  wire [2:0] _unuse_way_T_4 = ~_GEN_127 ? 3'h4 : 3'h0; // @[d_cache.scala 98:108]
  wire [2:0] _unuse_way_T_5 = ~_GEN_95 ? 3'h3 : _unuse_way_T_4; // @[d_cache.scala 98:79]
  wire [2:0] _unuse_way_T_6 = ~_GEN_63 ? 3'h2 : _unuse_way_T_5; // @[d_cache.scala 98:50]
  wire [2:0] unuse_way = ~_GEN_31 ? 3'h1 : _unuse_way_T_6; // @[d_cache.scala 98:21]
  reg [3:0] state; // @[d_cache.scala 100:24]
  wire  _T_1 = io_from_lsu_araddr >= 32'ha0000000; // @[d_cache.scala 108:41]
  wire [3:0] _GEN_129 = _T_1 ? 4'h8 : 4'h2; // @[d_cache.scala 114:58 115:27 117:27]
  wire  _T_6 = way0_hit | way1_hit | way2_hit | way3_hit; // @[d_cache.scala 123:46]
  wire [63:0] _ram_0_T = io_from_lsu_wdata & wmask; // @[d_cache.scala 135:53]
  wire [574:0] _GEN_5704 = {{511'd0}, _ram_0_T}; // @[d_cache.scala 135:62]
  wire [574:0] _ram_0_T_1 = _GEN_5704 << shift_bit; // @[d_cache.scala 135:62]
  wire [574:0] _GEN_5705 = {{511'd0}, wmask}; // @[d_cache.scala 135:102]
  wire [574:0] _ram_0_T_2 = _GEN_5705 << shift_bit; // @[d_cache.scala 135:102]
  wire [574:0] _ram_0_T_3 = ~_ram_0_T_2; // @[d_cache.scala 135:94]
  wire [511:0] _GEN_136 = 4'h1 == index ? ram_0_1 : ram_0_0; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_137 = 4'h2 == index ? ram_0_2 : _GEN_136; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_138 = 4'h3 == index ? ram_0_3 : _GEN_137; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_139 = 4'h4 == index ? ram_0_4 : _GEN_138; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_140 = 4'h5 == index ? ram_0_5 : _GEN_139; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_141 = 4'h6 == index ? ram_0_6 : _GEN_140; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_142 = 4'h7 == index ? ram_0_7 : _GEN_141; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_143 = 4'h8 == index ? ram_0_8 : _GEN_142; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_144 = 4'h9 == index ? ram_0_9 : _GEN_143; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_145 = 4'ha == index ? ram_0_10 : _GEN_144; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_146 = 4'hb == index ? ram_0_11 : _GEN_145; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_147 = 4'hc == index ? ram_0_12 : _GEN_146; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_148 = 4'hd == index ? ram_0_13 : _GEN_147; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_149 = 4'he == index ? ram_0_14 : _GEN_148; // @[d_cache.scala 135:{92,92}]
  wire [511:0] _GEN_150 = 4'hf == index ? ram_0_15 : _GEN_149; // @[d_cache.scala 135:{92,92}]
  wire [574:0] _GEN_5350 = {{63'd0}, _GEN_150}; // @[d_cache.scala 135:92]
  wire [574:0] _ram_0_T_4 = _GEN_5350 & _ram_0_T_3; // @[d_cache.scala 135:92]
  wire [574:0] _ram_0_T_5 = _ram_0_T_1 | _ram_0_T_4; // @[d_cache.scala 135:76]
  wire [511:0] _GEN_151 = 4'h0 == index ? _ram_0_T_5[511:0] : ram_0_0; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_152 = 4'h1 == index ? _ram_0_T_5[511:0] : ram_0_1; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_153 = 4'h2 == index ? _ram_0_T_5[511:0] : ram_0_2; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_154 = 4'h3 == index ? _ram_0_T_5[511:0] : ram_0_3; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_155 = 4'h4 == index ? _ram_0_T_5[511:0] : ram_0_4; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_156 = 4'h5 == index ? _ram_0_T_5[511:0] : ram_0_5; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_157 = 4'h6 == index ? _ram_0_T_5[511:0] : ram_0_6; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_158 = 4'h7 == index ? _ram_0_T_5[511:0] : ram_0_7; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_159 = 4'h8 == index ? _ram_0_T_5[511:0] : ram_0_8; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_160 = 4'h9 == index ? _ram_0_T_5[511:0] : ram_0_9; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_161 = 4'ha == index ? _ram_0_T_5[511:0] : ram_0_10; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_162 = 4'hb == index ? _ram_0_T_5[511:0] : ram_0_11; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_163 = 4'hc == index ? _ram_0_T_5[511:0] : ram_0_12; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_164 = 4'hd == index ? _ram_0_T_5[511:0] : ram_0_13; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_165 = 4'he == index ? _ram_0_T_5[511:0] : ram_0_14; // @[d_cache.scala 135:{30,30} 19:24]
  wire [511:0] _GEN_166 = 4'hf == index ? _ram_0_T_5[511:0] : ram_0_15; // @[d_cache.scala 135:{30,30} 19:24]
  wire  _GEN_5351 = 4'h0 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_167 = 4'h0 == index | dirty_0_0; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5356 = 4'h1 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_168 = 4'h1 == index | dirty_0_1; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5357 = 4'h2 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_169 = 4'h2 == index | dirty_0_2; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5361 = 4'h3 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_170 = 4'h3 == index | dirty_0_3; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5365 = 4'h4 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_171 = 4'h4 == index | dirty_0_4; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5367 = 4'h5 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_172 = 4'h5 == index | dirty_0_5; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5369 = 4'h6 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_173 = 4'h6 == index | dirty_0_6; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5370 = 4'h7 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_174 = 4'h7 == index | dirty_0_7; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5374 = 4'h8 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_175 = 4'h8 == index | dirty_0_8; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5375 = 4'h9 == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_176 = 4'h9 == index | dirty_0_9; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5380 = 4'ha == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_177 = 4'ha == index | dirty_0_10; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5381 = 4'hb == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_178 = 4'hb == index | dirty_0_11; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5384 = 4'hc == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_179 = 4'hc == index | dirty_0_12; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5388 = 4'hd == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_180 = 4'hd == index | dirty_0_13; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5390 = 4'he == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_181 = 4'he == index | dirty_0_14; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_5392 = 4'hf == index; // @[d_cache.scala 136:{32,32} 34:26]
  wire  _GEN_182 = 4'hf == index | dirty_0_15; // @[d_cache.scala 136:{32,32} 34:26]
  wire [511:0] _GEN_184 = 4'h1 == index ? ram_1_1 : ram_1_0; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_185 = 4'h2 == index ? ram_1_2 : _GEN_184; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_186 = 4'h3 == index ? ram_1_3 : _GEN_185; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_187 = 4'h4 == index ? ram_1_4 : _GEN_186; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_188 = 4'h5 == index ? ram_1_5 : _GEN_187; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_189 = 4'h6 == index ? ram_1_6 : _GEN_188; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_190 = 4'h7 == index ? ram_1_7 : _GEN_189; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_191 = 4'h8 == index ? ram_1_8 : _GEN_190; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_192 = 4'h9 == index ? ram_1_9 : _GEN_191; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_193 = 4'ha == index ? ram_1_10 : _GEN_192; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_194 = 4'hb == index ? ram_1_11 : _GEN_193; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_195 = 4'hc == index ? ram_1_12 : _GEN_194; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_196 = 4'hd == index ? ram_1_13 : _GEN_195; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_197 = 4'he == index ? ram_1_14 : _GEN_196; // @[d_cache.scala 139:{92,92}]
  wire [511:0] _GEN_198 = 4'hf == index ? ram_1_15 : _GEN_197; // @[d_cache.scala 139:{92,92}]
  wire [574:0] _GEN_5393 = {{63'd0}, _GEN_198}; // @[d_cache.scala 139:92]
  wire [574:0] _ram_1_T_4 = _GEN_5393 & _ram_0_T_3; // @[d_cache.scala 139:92]
  wire [574:0] _ram_1_T_5 = _ram_0_T_1 | _ram_1_T_4; // @[d_cache.scala 139:76]
  wire [511:0] _GEN_199 = 4'h0 == index ? _ram_1_T_5[511:0] : ram_1_0; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_200 = 4'h1 == index ? _ram_1_T_5[511:0] : ram_1_1; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_201 = 4'h2 == index ? _ram_1_T_5[511:0] : ram_1_2; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_202 = 4'h3 == index ? _ram_1_T_5[511:0] : ram_1_3; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_203 = 4'h4 == index ? _ram_1_T_5[511:0] : ram_1_4; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_204 = 4'h5 == index ? _ram_1_T_5[511:0] : ram_1_5; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_205 = 4'h6 == index ? _ram_1_T_5[511:0] : ram_1_6; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_206 = 4'h7 == index ? _ram_1_T_5[511:0] : ram_1_7; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_207 = 4'h8 == index ? _ram_1_T_5[511:0] : ram_1_8; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_208 = 4'h9 == index ? _ram_1_T_5[511:0] : ram_1_9; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_209 = 4'ha == index ? _ram_1_T_5[511:0] : ram_1_10; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_210 = 4'hb == index ? _ram_1_T_5[511:0] : ram_1_11; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_211 = 4'hc == index ? _ram_1_T_5[511:0] : ram_1_12; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_212 = 4'hd == index ? _ram_1_T_5[511:0] : ram_1_13; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_213 = 4'he == index ? _ram_1_T_5[511:0] : ram_1_14; // @[d_cache.scala 139:{30,30} 20:24]
  wire [511:0] _GEN_214 = 4'hf == index ? _ram_1_T_5[511:0] : ram_1_15; // @[d_cache.scala 139:{30,30} 20:24]
  wire  _GEN_215 = _GEN_5351 | dirty_1_0; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_216 = _GEN_5356 | dirty_1_1; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_217 = _GEN_5357 | dirty_1_2; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_218 = _GEN_5361 | dirty_1_3; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_219 = _GEN_5365 | dirty_1_4; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_220 = _GEN_5367 | dirty_1_5; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_221 = _GEN_5369 | dirty_1_6; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_222 = _GEN_5370 | dirty_1_7; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_223 = _GEN_5374 | dirty_1_8; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_224 = _GEN_5375 | dirty_1_9; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_225 = _GEN_5380 | dirty_1_10; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_226 = _GEN_5381 | dirty_1_11; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_227 = _GEN_5384 | dirty_1_12; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_228 = _GEN_5388 | dirty_1_13; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_229 = _GEN_5390 | dirty_1_14; // @[d_cache.scala 140:{32,32} 35:26]
  wire  _GEN_230 = _GEN_5392 | dirty_1_15; // @[d_cache.scala 140:{32,32} 35:26]
  wire [511:0] _GEN_232 = 4'h1 == index ? ram_2_1 : ram_2_0; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_233 = 4'h2 == index ? ram_2_2 : _GEN_232; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_234 = 4'h3 == index ? ram_2_3 : _GEN_233; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_235 = 4'h4 == index ? ram_2_4 : _GEN_234; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_236 = 4'h5 == index ? ram_2_5 : _GEN_235; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_237 = 4'h6 == index ? ram_2_6 : _GEN_236; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_238 = 4'h7 == index ? ram_2_7 : _GEN_237; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_239 = 4'h8 == index ? ram_2_8 : _GEN_238; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_240 = 4'h9 == index ? ram_2_9 : _GEN_239; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_241 = 4'ha == index ? ram_2_10 : _GEN_240; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_242 = 4'hb == index ? ram_2_11 : _GEN_241; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_243 = 4'hc == index ? ram_2_12 : _GEN_242; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_244 = 4'hd == index ? ram_2_13 : _GEN_243; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_245 = 4'he == index ? ram_2_14 : _GEN_244; // @[d_cache.scala 143:{92,92}]
  wire [511:0] _GEN_246 = 4'hf == index ? ram_2_15 : _GEN_245; // @[d_cache.scala 143:{92,92}]
  wire [574:0] _GEN_5442 = {{63'd0}, _GEN_246}; // @[d_cache.scala 143:92]
  wire [574:0] _ram_2_T_4 = _GEN_5442 & _ram_0_T_3; // @[d_cache.scala 143:92]
  wire [574:0] _ram_2_T_5 = _ram_0_T_1 | _ram_2_T_4; // @[d_cache.scala 143:76]
  wire [511:0] _GEN_247 = 4'h0 == index ? _ram_2_T_5[511:0] : ram_2_0; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_248 = 4'h1 == index ? _ram_2_T_5[511:0] : ram_2_1; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_249 = 4'h2 == index ? _ram_2_T_5[511:0] : ram_2_2; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_250 = 4'h3 == index ? _ram_2_T_5[511:0] : ram_2_3; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_251 = 4'h4 == index ? _ram_2_T_5[511:0] : ram_2_4; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_252 = 4'h5 == index ? _ram_2_T_5[511:0] : ram_2_5; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_253 = 4'h6 == index ? _ram_2_T_5[511:0] : ram_2_6; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_254 = 4'h7 == index ? _ram_2_T_5[511:0] : ram_2_7; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_255 = 4'h8 == index ? _ram_2_T_5[511:0] : ram_2_8; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_256 = 4'h9 == index ? _ram_2_T_5[511:0] : ram_2_9; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_257 = 4'ha == index ? _ram_2_T_5[511:0] : ram_2_10; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_258 = 4'hb == index ? _ram_2_T_5[511:0] : ram_2_11; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_259 = 4'hc == index ? _ram_2_T_5[511:0] : ram_2_12; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_260 = 4'hd == index ? _ram_2_T_5[511:0] : ram_2_13; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_261 = 4'he == index ? _ram_2_T_5[511:0] : ram_2_14; // @[d_cache.scala 143:{30,30} 21:24]
  wire [511:0] _GEN_262 = 4'hf == index ? _ram_2_T_5[511:0] : ram_2_15; // @[d_cache.scala 143:{30,30} 21:24]
  wire  _GEN_263 = _GEN_5351 | dirty_2_0; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_264 = _GEN_5356 | dirty_2_1; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_265 = _GEN_5357 | dirty_2_2; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_266 = _GEN_5361 | dirty_2_3; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_267 = _GEN_5365 | dirty_2_4; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_268 = _GEN_5367 | dirty_2_5; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_269 = _GEN_5369 | dirty_2_6; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_270 = _GEN_5370 | dirty_2_7; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_271 = _GEN_5374 | dirty_2_8; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_272 = _GEN_5375 | dirty_2_9; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_273 = _GEN_5380 | dirty_2_10; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_274 = _GEN_5381 | dirty_2_11; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_275 = _GEN_5384 | dirty_2_12; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_276 = _GEN_5388 | dirty_2_13; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_277 = _GEN_5390 | dirty_2_14; // @[d_cache.scala 144:{32,32} 36:26]
  wire  _GEN_278 = _GEN_5392 | dirty_2_15; // @[d_cache.scala 144:{32,32} 36:26]
  wire [511:0] _GEN_280 = 4'h1 == index ? ram_3_1 : ram_3_0; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_281 = 4'h2 == index ? ram_3_2 : _GEN_280; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_282 = 4'h3 == index ? ram_3_3 : _GEN_281; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_283 = 4'h4 == index ? ram_3_4 : _GEN_282; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_284 = 4'h5 == index ? ram_3_5 : _GEN_283; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_285 = 4'h6 == index ? ram_3_6 : _GEN_284; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_286 = 4'h7 == index ? ram_3_7 : _GEN_285; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_287 = 4'h8 == index ? ram_3_8 : _GEN_286; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_288 = 4'h9 == index ? ram_3_9 : _GEN_287; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_289 = 4'ha == index ? ram_3_10 : _GEN_288; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_290 = 4'hb == index ? ram_3_11 : _GEN_289; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_291 = 4'hc == index ? ram_3_12 : _GEN_290; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_292 = 4'hd == index ? ram_3_13 : _GEN_291; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_293 = 4'he == index ? ram_3_14 : _GEN_292; // @[d_cache.scala 147:{92,92}]
  wire [511:0] _GEN_294 = 4'hf == index ? ram_3_15 : _GEN_293; // @[d_cache.scala 147:{92,92}]
  wire [574:0] _GEN_5480 = {{63'd0}, _GEN_294}; // @[d_cache.scala 147:92]
  wire [574:0] _ram_3_T_4 = _GEN_5480 & _ram_0_T_3; // @[d_cache.scala 147:92]
  wire [574:0] _ram_3_T_5 = _ram_0_T_1 | _ram_3_T_4; // @[d_cache.scala 147:76]
  wire [511:0] _GEN_295 = 4'h0 == index ? _ram_3_T_5[511:0] : ram_3_0; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_296 = 4'h1 == index ? _ram_3_T_5[511:0] : ram_3_1; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_297 = 4'h2 == index ? _ram_3_T_5[511:0] : ram_3_2; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_298 = 4'h3 == index ? _ram_3_T_5[511:0] : ram_3_3; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_299 = 4'h4 == index ? _ram_3_T_5[511:0] : ram_3_4; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_300 = 4'h5 == index ? _ram_3_T_5[511:0] : ram_3_5; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_301 = 4'h6 == index ? _ram_3_T_5[511:0] : ram_3_6; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_302 = 4'h7 == index ? _ram_3_T_5[511:0] : ram_3_7; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_303 = 4'h8 == index ? _ram_3_T_5[511:0] : ram_3_8; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_304 = 4'h9 == index ? _ram_3_T_5[511:0] : ram_3_9; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_305 = 4'ha == index ? _ram_3_T_5[511:0] : ram_3_10; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_306 = 4'hb == index ? _ram_3_T_5[511:0] : ram_3_11; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_307 = 4'hc == index ? _ram_3_T_5[511:0] : ram_3_12; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_308 = 4'hd == index ? _ram_3_T_5[511:0] : ram_3_13; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_309 = 4'he == index ? _ram_3_T_5[511:0] : ram_3_14; // @[d_cache.scala 147:{30,30} 22:24]
  wire [511:0] _GEN_310 = 4'hf == index ? _ram_3_T_5[511:0] : ram_3_15; // @[d_cache.scala 147:{30,30} 22:24]
  wire  _GEN_311 = _GEN_5351 | dirty_3_0; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_312 = _GEN_5356 | dirty_3_1; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_313 = _GEN_5357 | dirty_3_2; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_314 = _GEN_5361 | dirty_3_3; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_315 = _GEN_5365 | dirty_3_4; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_316 = _GEN_5367 | dirty_3_5; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_317 = _GEN_5369 | dirty_3_6; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_318 = _GEN_5370 | dirty_3_7; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_319 = _GEN_5374 | dirty_3_8; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_320 = _GEN_5375 | dirty_3_9; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_321 = _GEN_5380 | dirty_3_10; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_322 = _GEN_5381 | dirty_3_11; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_323 = _GEN_5384 | dirty_3_12; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_324 = _GEN_5388 | dirty_3_13; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_325 = _GEN_5390 | dirty_3_14; // @[d_cache.scala 148:{32,32} 37:26]
  wire  _GEN_326 = _GEN_5392 | dirty_3_15; // @[d_cache.scala 148:{32,32} 37:26]
  wire [3:0] _GEN_327 = way3_hit ? 4'h0 : 4'h4; // @[d_cache.scala 145:33 146:23 150:23]
  wire [511:0] _GEN_328 = way3_hit ? _GEN_295 : ram_3_0; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_329 = way3_hit ? _GEN_296 : ram_3_1; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_330 = way3_hit ? _GEN_297 : ram_3_2; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_331 = way3_hit ? _GEN_298 : ram_3_3; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_332 = way3_hit ? _GEN_299 : ram_3_4; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_333 = way3_hit ? _GEN_300 : ram_3_5; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_334 = way3_hit ? _GEN_301 : ram_3_6; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_335 = way3_hit ? _GEN_302 : ram_3_7; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_336 = way3_hit ? _GEN_303 : ram_3_8; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_337 = way3_hit ? _GEN_304 : ram_3_9; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_338 = way3_hit ? _GEN_305 : ram_3_10; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_339 = way3_hit ? _GEN_306 : ram_3_11; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_340 = way3_hit ? _GEN_307 : ram_3_12; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_341 = way3_hit ? _GEN_308 : ram_3_13; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_342 = way3_hit ? _GEN_309 : ram_3_14; // @[d_cache.scala 145:33 22:24]
  wire [511:0] _GEN_343 = way3_hit ? _GEN_310 : ram_3_15; // @[d_cache.scala 145:33 22:24]
  wire  _GEN_344 = way3_hit ? _GEN_311 : dirty_3_0; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_345 = way3_hit ? _GEN_312 : dirty_3_1; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_346 = way3_hit ? _GEN_313 : dirty_3_2; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_347 = way3_hit ? _GEN_314 : dirty_3_3; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_348 = way3_hit ? _GEN_315 : dirty_3_4; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_349 = way3_hit ? _GEN_316 : dirty_3_5; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_350 = way3_hit ? _GEN_317 : dirty_3_6; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_351 = way3_hit ? _GEN_318 : dirty_3_7; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_352 = way3_hit ? _GEN_319 : dirty_3_8; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_353 = way3_hit ? _GEN_320 : dirty_3_9; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_354 = way3_hit ? _GEN_321 : dirty_3_10; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_355 = way3_hit ? _GEN_322 : dirty_3_11; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_356 = way3_hit ? _GEN_323 : dirty_3_12; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_357 = way3_hit ? _GEN_324 : dirty_3_13; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_358 = way3_hit ? _GEN_325 : dirty_3_14; // @[d_cache.scala 145:33 37:26]
  wire  _GEN_359 = way3_hit ? _GEN_326 : dirty_3_15; // @[d_cache.scala 145:33 37:26]
  wire [3:0] _GEN_360 = way2_hit ? 4'h0 : _GEN_327; // @[d_cache.scala 141:33 142:23]
  wire [511:0] _GEN_361 = way2_hit ? _GEN_247 : ram_2_0; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_362 = way2_hit ? _GEN_248 : ram_2_1; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_363 = way2_hit ? _GEN_249 : ram_2_2; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_364 = way2_hit ? _GEN_250 : ram_2_3; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_365 = way2_hit ? _GEN_251 : ram_2_4; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_366 = way2_hit ? _GEN_252 : ram_2_5; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_367 = way2_hit ? _GEN_253 : ram_2_6; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_368 = way2_hit ? _GEN_254 : ram_2_7; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_369 = way2_hit ? _GEN_255 : ram_2_8; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_370 = way2_hit ? _GEN_256 : ram_2_9; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_371 = way2_hit ? _GEN_257 : ram_2_10; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_372 = way2_hit ? _GEN_258 : ram_2_11; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_373 = way2_hit ? _GEN_259 : ram_2_12; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_374 = way2_hit ? _GEN_260 : ram_2_13; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_375 = way2_hit ? _GEN_261 : ram_2_14; // @[d_cache.scala 141:33 21:24]
  wire [511:0] _GEN_376 = way2_hit ? _GEN_262 : ram_2_15; // @[d_cache.scala 141:33 21:24]
  wire  _GEN_377 = way2_hit ? _GEN_263 : dirty_2_0; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_378 = way2_hit ? _GEN_264 : dirty_2_1; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_379 = way2_hit ? _GEN_265 : dirty_2_2; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_380 = way2_hit ? _GEN_266 : dirty_2_3; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_381 = way2_hit ? _GEN_267 : dirty_2_4; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_382 = way2_hit ? _GEN_268 : dirty_2_5; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_383 = way2_hit ? _GEN_269 : dirty_2_6; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_384 = way2_hit ? _GEN_270 : dirty_2_7; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_385 = way2_hit ? _GEN_271 : dirty_2_8; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_386 = way2_hit ? _GEN_272 : dirty_2_9; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_387 = way2_hit ? _GEN_273 : dirty_2_10; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_388 = way2_hit ? _GEN_274 : dirty_2_11; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_389 = way2_hit ? _GEN_275 : dirty_2_12; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_390 = way2_hit ? _GEN_276 : dirty_2_13; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_391 = way2_hit ? _GEN_277 : dirty_2_14; // @[d_cache.scala 141:33 36:26]
  wire  _GEN_392 = way2_hit ? _GEN_278 : dirty_2_15; // @[d_cache.scala 141:33 36:26]
  wire [511:0] _GEN_393 = way2_hit ? ram_3_0 : _GEN_328; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_394 = way2_hit ? ram_3_1 : _GEN_329; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_395 = way2_hit ? ram_3_2 : _GEN_330; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_396 = way2_hit ? ram_3_3 : _GEN_331; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_397 = way2_hit ? ram_3_4 : _GEN_332; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_398 = way2_hit ? ram_3_5 : _GEN_333; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_399 = way2_hit ? ram_3_6 : _GEN_334; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_400 = way2_hit ? ram_3_7 : _GEN_335; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_401 = way2_hit ? ram_3_8 : _GEN_336; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_402 = way2_hit ? ram_3_9 : _GEN_337; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_403 = way2_hit ? ram_3_10 : _GEN_338; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_404 = way2_hit ? ram_3_11 : _GEN_339; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_405 = way2_hit ? ram_3_12 : _GEN_340; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_406 = way2_hit ? ram_3_13 : _GEN_341; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_407 = way2_hit ? ram_3_14 : _GEN_342; // @[d_cache.scala 141:33 22:24]
  wire [511:0] _GEN_408 = way2_hit ? ram_3_15 : _GEN_343; // @[d_cache.scala 141:33 22:24]
  wire  _GEN_409 = way2_hit ? dirty_3_0 : _GEN_344; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_410 = way2_hit ? dirty_3_1 : _GEN_345; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_411 = way2_hit ? dirty_3_2 : _GEN_346; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_412 = way2_hit ? dirty_3_3 : _GEN_347; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_413 = way2_hit ? dirty_3_4 : _GEN_348; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_414 = way2_hit ? dirty_3_5 : _GEN_349; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_415 = way2_hit ? dirty_3_6 : _GEN_350; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_416 = way2_hit ? dirty_3_7 : _GEN_351; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_417 = way2_hit ? dirty_3_8 : _GEN_352; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_418 = way2_hit ? dirty_3_9 : _GEN_353; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_419 = way2_hit ? dirty_3_10 : _GEN_354; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_420 = way2_hit ? dirty_3_11 : _GEN_355; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_421 = way2_hit ? dirty_3_12 : _GEN_356; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_422 = way2_hit ? dirty_3_13 : _GEN_357; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_423 = way2_hit ? dirty_3_14 : _GEN_358; // @[d_cache.scala 141:33 37:26]
  wire  _GEN_424 = way2_hit ? dirty_3_15 : _GEN_359; // @[d_cache.scala 141:33 37:26]
  wire [3:0] _GEN_425 = way1_hit ? 4'h0 : _GEN_360; // @[d_cache.scala 137:33 138:23]
  wire [511:0] _GEN_426 = way1_hit ? _GEN_199 : ram_1_0; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_427 = way1_hit ? _GEN_200 : ram_1_1; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_428 = way1_hit ? _GEN_201 : ram_1_2; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_429 = way1_hit ? _GEN_202 : ram_1_3; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_430 = way1_hit ? _GEN_203 : ram_1_4; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_431 = way1_hit ? _GEN_204 : ram_1_5; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_432 = way1_hit ? _GEN_205 : ram_1_6; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_433 = way1_hit ? _GEN_206 : ram_1_7; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_434 = way1_hit ? _GEN_207 : ram_1_8; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_435 = way1_hit ? _GEN_208 : ram_1_9; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_436 = way1_hit ? _GEN_209 : ram_1_10; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_437 = way1_hit ? _GEN_210 : ram_1_11; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_438 = way1_hit ? _GEN_211 : ram_1_12; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_439 = way1_hit ? _GEN_212 : ram_1_13; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_440 = way1_hit ? _GEN_213 : ram_1_14; // @[d_cache.scala 137:33 20:24]
  wire [511:0] _GEN_441 = way1_hit ? _GEN_214 : ram_1_15; // @[d_cache.scala 137:33 20:24]
  wire  _GEN_442 = way1_hit ? _GEN_215 : dirty_1_0; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_443 = way1_hit ? _GEN_216 : dirty_1_1; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_444 = way1_hit ? _GEN_217 : dirty_1_2; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_445 = way1_hit ? _GEN_218 : dirty_1_3; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_446 = way1_hit ? _GEN_219 : dirty_1_4; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_447 = way1_hit ? _GEN_220 : dirty_1_5; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_448 = way1_hit ? _GEN_221 : dirty_1_6; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_449 = way1_hit ? _GEN_222 : dirty_1_7; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_450 = way1_hit ? _GEN_223 : dirty_1_8; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_451 = way1_hit ? _GEN_224 : dirty_1_9; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_452 = way1_hit ? _GEN_225 : dirty_1_10; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_453 = way1_hit ? _GEN_226 : dirty_1_11; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_454 = way1_hit ? _GEN_227 : dirty_1_12; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_455 = way1_hit ? _GEN_228 : dirty_1_13; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_456 = way1_hit ? _GEN_229 : dirty_1_14; // @[d_cache.scala 137:33 35:26]
  wire  _GEN_457 = way1_hit ? _GEN_230 : dirty_1_15; // @[d_cache.scala 137:33 35:26]
  wire [511:0] _GEN_458 = way1_hit ? ram_2_0 : _GEN_361; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_459 = way1_hit ? ram_2_1 : _GEN_362; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_460 = way1_hit ? ram_2_2 : _GEN_363; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_461 = way1_hit ? ram_2_3 : _GEN_364; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_462 = way1_hit ? ram_2_4 : _GEN_365; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_463 = way1_hit ? ram_2_5 : _GEN_366; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_464 = way1_hit ? ram_2_6 : _GEN_367; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_465 = way1_hit ? ram_2_7 : _GEN_368; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_466 = way1_hit ? ram_2_8 : _GEN_369; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_467 = way1_hit ? ram_2_9 : _GEN_370; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_468 = way1_hit ? ram_2_10 : _GEN_371; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_469 = way1_hit ? ram_2_11 : _GEN_372; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_470 = way1_hit ? ram_2_12 : _GEN_373; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_471 = way1_hit ? ram_2_13 : _GEN_374; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_472 = way1_hit ? ram_2_14 : _GEN_375; // @[d_cache.scala 137:33 21:24]
  wire [511:0] _GEN_473 = way1_hit ? ram_2_15 : _GEN_376; // @[d_cache.scala 137:33 21:24]
  wire  _GEN_474 = way1_hit ? dirty_2_0 : _GEN_377; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_475 = way1_hit ? dirty_2_1 : _GEN_378; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_476 = way1_hit ? dirty_2_2 : _GEN_379; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_477 = way1_hit ? dirty_2_3 : _GEN_380; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_478 = way1_hit ? dirty_2_4 : _GEN_381; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_479 = way1_hit ? dirty_2_5 : _GEN_382; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_480 = way1_hit ? dirty_2_6 : _GEN_383; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_481 = way1_hit ? dirty_2_7 : _GEN_384; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_482 = way1_hit ? dirty_2_8 : _GEN_385; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_483 = way1_hit ? dirty_2_9 : _GEN_386; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_484 = way1_hit ? dirty_2_10 : _GEN_387; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_485 = way1_hit ? dirty_2_11 : _GEN_388; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_486 = way1_hit ? dirty_2_12 : _GEN_389; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_487 = way1_hit ? dirty_2_13 : _GEN_390; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_488 = way1_hit ? dirty_2_14 : _GEN_391; // @[d_cache.scala 137:33 36:26]
  wire  _GEN_489 = way1_hit ? dirty_2_15 : _GEN_392; // @[d_cache.scala 137:33 36:26]
  wire [511:0] _GEN_490 = way1_hit ? ram_3_0 : _GEN_393; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_491 = way1_hit ? ram_3_1 : _GEN_394; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_492 = way1_hit ? ram_3_2 : _GEN_395; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_493 = way1_hit ? ram_3_3 : _GEN_396; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_494 = way1_hit ? ram_3_4 : _GEN_397; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_495 = way1_hit ? ram_3_5 : _GEN_398; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_496 = way1_hit ? ram_3_6 : _GEN_399; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_497 = way1_hit ? ram_3_7 : _GEN_400; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_498 = way1_hit ? ram_3_8 : _GEN_401; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_499 = way1_hit ? ram_3_9 : _GEN_402; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_500 = way1_hit ? ram_3_10 : _GEN_403; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_501 = way1_hit ? ram_3_11 : _GEN_404; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_502 = way1_hit ? ram_3_12 : _GEN_405; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_503 = way1_hit ? ram_3_13 : _GEN_406; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_504 = way1_hit ? ram_3_14 : _GEN_407; // @[d_cache.scala 137:33 22:24]
  wire [511:0] _GEN_505 = way1_hit ? ram_3_15 : _GEN_408; // @[d_cache.scala 137:33 22:24]
  wire  _GEN_506 = way1_hit ? dirty_3_0 : _GEN_409; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_507 = way1_hit ? dirty_3_1 : _GEN_410; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_508 = way1_hit ? dirty_3_2 : _GEN_411; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_509 = way1_hit ? dirty_3_3 : _GEN_412; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_510 = way1_hit ? dirty_3_4 : _GEN_413; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_511 = way1_hit ? dirty_3_5 : _GEN_414; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_512 = way1_hit ? dirty_3_6 : _GEN_415; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_513 = way1_hit ? dirty_3_7 : _GEN_416; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_514 = way1_hit ? dirty_3_8 : _GEN_417; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_515 = way1_hit ? dirty_3_9 : _GEN_418; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_516 = way1_hit ? dirty_3_10 : _GEN_419; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_517 = way1_hit ? dirty_3_11 : _GEN_420; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_518 = way1_hit ? dirty_3_12 : _GEN_421; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_519 = way1_hit ? dirty_3_13 : _GEN_422; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_520 = way1_hit ? dirty_3_14 : _GEN_423; // @[d_cache.scala 137:33 37:26]
  wire  _GEN_521 = way1_hit ? dirty_3_15 : _GEN_424; // @[d_cache.scala 137:33 37:26]
  wire [3:0] _GEN_522 = way0_hit ? 4'h0 : _GEN_425; // @[d_cache.scala 133:27 134:23]
  wire [511:0] _GEN_523 = way0_hit ? _GEN_151 : ram_0_0; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_524 = way0_hit ? _GEN_152 : ram_0_1; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_525 = way0_hit ? _GEN_153 : ram_0_2; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_526 = way0_hit ? _GEN_154 : ram_0_3; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_527 = way0_hit ? _GEN_155 : ram_0_4; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_528 = way0_hit ? _GEN_156 : ram_0_5; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_529 = way0_hit ? _GEN_157 : ram_0_6; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_530 = way0_hit ? _GEN_158 : ram_0_7; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_531 = way0_hit ? _GEN_159 : ram_0_8; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_532 = way0_hit ? _GEN_160 : ram_0_9; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_533 = way0_hit ? _GEN_161 : ram_0_10; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_534 = way0_hit ? _GEN_162 : ram_0_11; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_535 = way0_hit ? _GEN_163 : ram_0_12; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_536 = way0_hit ? _GEN_164 : ram_0_13; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_537 = way0_hit ? _GEN_165 : ram_0_14; // @[d_cache.scala 133:27 19:24]
  wire [511:0] _GEN_538 = way0_hit ? _GEN_166 : ram_0_15; // @[d_cache.scala 133:27 19:24]
  wire  _GEN_539 = way0_hit ? _GEN_167 : dirty_0_0; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_540 = way0_hit ? _GEN_168 : dirty_0_1; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_541 = way0_hit ? _GEN_169 : dirty_0_2; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_542 = way0_hit ? _GEN_170 : dirty_0_3; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_543 = way0_hit ? _GEN_171 : dirty_0_4; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_544 = way0_hit ? _GEN_172 : dirty_0_5; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_545 = way0_hit ? _GEN_173 : dirty_0_6; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_546 = way0_hit ? _GEN_174 : dirty_0_7; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_547 = way0_hit ? _GEN_175 : dirty_0_8; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_548 = way0_hit ? _GEN_176 : dirty_0_9; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_549 = way0_hit ? _GEN_177 : dirty_0_10; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_550 = way0_hit ? _GEN_178 : dirty_0_11; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_551 = way0_hit ? _GEN_179 : dirty_0_12; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_552 = way0_hit ? _GEN_180 : dirty_0_13; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_553 = way0_hit ? _GEN_181 : dirty_0_14; // @[d_cache.scala 133:27 34:26]
  wire  _GEN_554 = way0_hit ? _GEN_182 : dirty_0_15; // @[d_cache.scala 133:27 34:26]
  wire [511:0] _GEN_555 = way0_hit ? ram_1_0 : _GEN_426; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_556 = way0_hit ? ram_1_1 : _GEN_427; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_557 = way0_hit ? ram_1_2 : _GEN_428; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_558 = way0_hit ? ram_1_3 : _GEN_429; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_559 = way0_hit ? ram_1_4 : _GEN_430; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_560 = way0_hit ? ram_1_5 : _GEN_431; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_561 = way0_hit ? ram_1_6 : _GEN_432; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_562 = way0_hit ? ram_1_7 : _GEN_433; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_563 = way0_hit ? ram_1_8 : _GEN_434; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_564 = way0_hit ? ram_1_9 : _GEN_435; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_565 = way0_hit ? ram_1_10 : _GEN_436; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_566 = way0_hit ? ram_1_11 : _GEN_437; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_567 = way0_hit ? ram_1_12 : _GEN_438; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_568 = way0_hit ? ram_1_13 : _GEN_439; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_569 = way0_hit ? ram_1_14 : _GEN_440; // @[d_cache.scala 133:27 20:24]
  wire [511:0] _GEN_570 = way0_hit ? ram_1_15 : _GEN_441; // @[d_cache.scala 133:27 20:24]
  wire  _GEN_571 = way0_hit ? dirty_1_0 : _GEN_442; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_572 = way0_hit ? dirty_1_1 : _GEN_443; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_573 = way0_hit ? dirty_1_2 : _GEN_444; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_574 = way0_hit ? dirty_1_3 : _GEN_445; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_575 = way0_hit ? dirty_1_4 : _GEN_446; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_576 = way0_hit ? dirty_1_5 : _GEN_447; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_577 = way0_hit ? dirty_1_6 : _GEN_448; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_578 = way0_hit ? dirty_1_7 : _GEN_449; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_579 = way0_hit ? dirty_1_8 : _GEN_450; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_580 = way0_hit ? dirty_1_9 : _GEN_451; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_581 = way0_hit ? dirty_1_10 : _GEN_452; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_582 = way0_hit ? dirty_1_11 : _GEN_453; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_583 = way0_hit ? dirty_1_12 : _GEN_454; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_584 = way0_hit ? dirty_1_13 : _GEN_455; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_585 = way0_hit ? dirty_1_14 : _GEN_456; // @[d_cache.scala 133:27 35:26]
  wire  _GEN_586 = way0_hit ? dirty_1_15 : _GEN_457; // @[d_cache.scala 133:27 35:26]
  wire [511:0] _GEN_587 = way0_hit ? ram_2_0 : _GEN_458; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_588 = way0_hit ? ram_2_1 : _GEN_459; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_589 = way0_hit ? ram_2_2 : _GEN_460; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_590 = way0_hit ? ram_2_3 : _GEN_461; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_591 = way0_hit ? ram_2_4 : _GEN_462; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_592 = way0_hit ? ram_2_5 : _GEN_463; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_593 = way0_hit ? ram_2_6 : _GEN_464; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_594 = way0_hit ? ram_2_7 : _GEN_465; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_595 = way0_hit ? ram_2_8 : _GEN_466; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_596 = way0_hit ? ram_2_9 : _GEN_467; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_597 = way0_hit ? ram_2_10 : _GEN_468; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_598 = way0_hit ? ram_2_11 : _GEN_469; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_599 = way0_hit ? ram_2_12 : _GEN_470; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_600 = way0_hit ? ram_2_13 : _GEN_471; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_601 = way0_hit ? ram_2_14 : _GEN_472; // @[d_cache.scala 133:27 21:24]
  wire [511:0] _GEN_602 = way0_hit ? ram_2_15 : _GEN_473; // @[d_cache.scala 133:27 21:24]
  wire  _GEN_603 = way0_hit ? dirty_2_0 : _GEN_474; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_604 = way0_hit ? dirty_2_1 : _GEN_475; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_605 = way0_hit ? dirty_2_2 : _GEN_476; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_606 = way0_hit ? dirty_2_3 : _GEN_477; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_607 = way0_hit ? dirty_2_4 : _GEN_478; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_608 = way0_hit ? dirty_2_5 : _GEN_479; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_609 = way0_hit ? dirty_2_6 : _GEN_480; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_610 = way0_hit ? dirty_2_7 : _GEN_481; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_611 = way0_hit ? dirty_2_8 : _GEN_482; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_612 = way0_hit ? dirty_2_9 : _GEN_483; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_613 = way0_hit ? dirty_2_10 : _GEN_484; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_614 = way0_hit ? dirty_2_11 : _GEN_485; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_615 = way0_hit ? dirty_2_12 : _GEN_486; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_616 = way0_hit ? dirty_2_13 : _GEN_487; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_617 = way0_hit ? dirty_2_14 : _GEN_488; // @[d_cache.scala 133:27 36:26]
  wire  _GEN_618 = way0_hit ? dirty_2_15 : _GEN_489; // @[d_cache.scala 133:27 36:26]
  wire [511:0] _GEN_619 = way0_hit ? ram_3_0 : _GEN_490; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_620 = way0_hit ? ram_3_1 : _GEN_491; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_621 = way0_hit ? ram_3_2 : _GEN_492; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_622 = way0_hit ? ram_3_3 : _GEN_493; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_623 = way0_hit ? ram_3_4 : _GEN_494; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_624 = way0_hit ? ram_3_5 : _GEN_495; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_625 = way0_hit ? ram_3_6 : _GEN_496; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_626 = way0_hit ? ram_3_7 : _GEN_497; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_627 = way0_hit ? ram_3_8 : _GEN_498; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_628 = way0_hit ? ram_3_9 : _GEN_499; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_629 = way0_hit ? ram_3_10 : _GEN_500; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_630 = way0_hit ? ram_3_11 : _GEN_501; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_631 = way0_hit ? ram_3_12 : _GEN_502; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_632 = way0_hit ? ram_3_13 : _GEN_503; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_633 = way0_hit ? ram_3_14 : _GEN_504; // @[d_cache.scala 133:27 22:24]
  wire [511:0] _GEN_634 = way0_hit ? ram_3_15 : _GEN_505; // @[d_cache.scala 133:27 22:24]
  wire  _GEN_635 = way0_hit ? dirty_3_0 : _GEN_506; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_636 = way0_hit ? dirty_3_1 : _GEN_507; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_637 = way0_hit ? dirty_3_2 : _GEN_508; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_638 = way0_hit ? dirty_3_3 : _GEN_509; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_639 = way0_hit ? dirty_3_4 : _GEN_510; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_640 = way0_hit ? dirty_3_5 : _GEN_511; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_641 = way0_hit ? dirty_3_6 : _GEN_512; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_642 = way0_hit ? dirty_3_7 : _GEN_513; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_643 = way0_hit ? dirty_3_8 : _GEN_514; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_644 = way0_hit ? dirty_3_9 : _GEN_515; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_645 = way0_hit ? dirty_3_10 : _GEN_516; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_646 = way0_hit ? dirty_3_11 : _GEN_517; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_647 = way0_hit ? dirty_3_12 : _GEN_518; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_648 = way0_hit ? dirty_3_13 : _GEN_519; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_649 = way0_hit ? dirty_3_14 : _GEN_520; // @[d_cache.scala 133:27 37:26]
  wire  _GEN_650 = way0_hit ? dirty_3_15 : _GEN_521; // @[d_cache.scala 133:27 37:26]
  wire [63:0] _GEN_651 = 3'h0 == receive_num ? io_from_axi_rdata : receive_data_0; // @[d_cache.scala 155:{43,43} 50:31]
  wire [63:0] _GEN_652 = 3'h1 == receive_num ? io_from_axi_rdata : receive_data_1; // @[d_cache.scala 155:{43,43} 50:31]
  wire [63:0] _GEN_653 = 3'h2 == receive_num ? io_from_axi_rdata : receive_data_2; // @[d_cache.scala 155:{43,43} 50:31]
  wire [63:0] _GEN_654 = 3'h3 == receive_num ? io_from_axi_rdata : receive_data_3; // @[d_cache.scala 155:{43,43} 50:31]
  wire [63:0] _GEN_655 = 3'h4 == receive_num ? io_from_axi_rdata : receive_data_4; // @[d_cache.scala 155:{43,43} 50:31]
  wire [63:0] _GEN_656 = 3'h5 == receive_num ? io_from_axi_rdata : receive_data_5; // @[d_cache.scala 155:{43,43} 50:31]
  wire [63:0] _GEN_657 = 3'h6 == receive_num ? io_from_axi_rdata : receive_data_6; // @[d_cache.scala 155:{43,43} 50:31]
  wire [63:0] _GEN_658 = 3'h7 == receive_num ? io_from_axi_rdata : receive_data_7; // @[d_cache.scala 155:{43,43} 50:31]
  wire [2:0] _receive_num_T_1 = receive_num + 3'h1; // @[d_cache.scala 156:44]
  wire [3:0] _GEN_659 = io_from_axi_rlast ? 4'h5 : state; // @[d_cache.scala 100:24 157:40 158:27]
  wire [63:0] _GEN_660 = io_from_axi_rvalid ? _GEN_651 : receive_data_0; // @[d_cache.scala 154:37 50:31]
  wire [63:0] _GEN_661 = io_from_axi_rvalid ? _GEN_652 : receive_data_1; // @[d_cache.scala 154:37 50:31]
  wire [63:0] _GEN_662 = io_from_axi_rvalid ? _GEN_653 : receive_data_2; // @[d_cache.scala 154:37 50:31]
  wire [63:0] _GEN_663 = io_from_axi_rvalid ? _GEN_654 : receive_data_3; // @[d_cache.scala 154:37 50:31]
  wire [63:0] _GEN_664 = io_from_axi_rvalid ? _GEN_655 : receive_data_4; // @[d_cache.scala 154:37 50:31]
  wire [63:0] _GEN_665 = io_from_axi_rvalid ? _GEN_656 : receive_data_5; // @[d_cache.scala 154:37 50:31]
  wire [63:0] _GEN_666 = io_from_axi_rvalid ? _GEN_657 : receive_data_6; // @[d_cache.scala 154:37 50:31]
  wire [63:0] _GEN_667 = io_from_axi_rvalid ? _GEN_658 : receive_data_7; // @[d_cache.scala 154:37 50:31]
  wire [2:0] _GEN_668 = io_from_axi_rvalid ? _receive_num_T_1 : receive_num; // @[d_cache.scala 154:37 156:29 51:30]
  wire [3:0] _GEN_669 = io_from_axi_rvalid ? _GEN_659 : state; // @[d_cache.scala 100:24 154:37]
  wire [3:0] _GEN_670 = io_from_axi_bvalid ? 4'h0 : state; // @[d_cache.scala 163:37 164:23 100:24]
  wire [511:0] _ram_0_T_6 = {receive_data_7,receive_data_6,receive_data_5,receive_data_4,receive_data_3,receive_data_2,
    receive_data_1,receive_data_0}; // @[Cat.scala 31:58]
  wire [511:0] _GEN_671 = 4'h0 == index ? _ram_0_T_6 : ram_0_0; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_672 = 4'h1 == index ? _ram_0_T_6 : ram_0_1; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_673 = 4'h2 == index ? _ram_0_T_6 : ram_0_2; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_674 = 4'h3 == index ? _ram_0_T_6 : ram_0_3; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_675 = 4'h4 == index ? _ram_0_T_6 : ram_0_4; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_676 = 4'h5 == index ? _ram_0_T_6 : ram_0_5; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_677 = 4'h6 == index ? _ram_0_T_6 : ram_0_6; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_678 = 4'h7 == index ? _ram_0_T_6 : ram_0_7; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_679 = 4'h8 == index ? _ram_0_T_6 : ram_0_8; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_680 = 4'h9 == index ? _ram_0_T_6 : ram_0_9; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_681 = 4'ha == index ? _ram_0_T_6 : ram_0_10; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_682 = 4'hb == index ? _ram_0_T_6 : ram_0_11; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_683 = 4'hc == index ? _ram_0_T_6 : ram_0_12; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_684 = 4'hd == index ? _ram_0_T_6 : ram_0_13; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_685 = 4'he == index ? _ram_0_T_6 : ram_0_14; // @[d_cache.scala 170:{30,30} 19:24]
  wire [511:0] _GEN_686 = 4'hf == index ? _ram_0_T_6 : ram_0_15; // @[d_cache.scala 170:{30,30} 19:24]
  wire [31:0] _GEN_687 = 4'h0 == index ? _GEN_5341 : tag_0_0; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_688 = 4'h1 == index ? _GEN_5341 : tag_0_1; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_689 = 4'h2 == index ? _GEN_5341 : tag_0_2; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_690 = 4'h3 == index ? _GEN_5341 : tag_0_3; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_691 = 4'h4 == index ? _GEN_5341 : tag_0_4; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_692 = 4'h5 == index ? _GEN_5341 : tag_0_5; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_693 = 4'h6 == index ? _GEN_5341 : tag_0_6; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_694 = 4'h7 == index ? _GEN_5341 : tag_0_7; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_695 = 4'h8 == index ? _GEN_5341 : tag_0_8; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_696 = 4'h9 == index ? _GEN_5341 : tag_0_9; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_697 = 4'ha == index ? _GEN_5341 : tag_0_10; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_698 = 4'hb == index ? _GEN_5341 : tag_0_11; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_699 = 4'hc == index ? _GEN_5341 : tag_0_12; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_700 = 4'hd == index ? _GEN_5341 : tag_0_13; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_701 = 4'he == index ? _GEN_5341 : tag_0_14; // @[d_cache.scala 171:{30,30} 24:24]
  wire [31:0] _GEN_702 = 4'hf == index ? _GEN_5341 : tag_0_15; // @[d_cache.scala 171:{30,30} 24:24]
  wire  _GEN_703 = _GEN_5351 | valid_0_0; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_704 = _GEN_5356 | valid_0_1; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_705 = _GEN_5357 | valid_0_2; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_706 = _GEN_5361 | valid_0_3; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_707 = _GEN_5365 | valid_0_4; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_708 = _GEN_5367 | valid_0_5; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_709 = _GEN_5369 | valid_0_6; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_710 = _GEN_5370 | valid_0_7; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_711 = _GEN_5374 | valid_0_8; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_712 = _GEN_5375 | valid_0_9; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_713 = _GEN_5380 | valid_0_10; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_714 = _GEN_5381 | valid_0_11; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_715 = _GEN_5384 | valid_0_12; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_716 = _GEN_5388 | valid_0_13; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_717 = _GEN_5390 | valid_0_14; // @[d_cache.scala 172:{32,32} 29:26]
  wire  _GEN_718 = _GEN_5392 | valid_0_15; // @[d_cache.scala 172:{32,32} 29:26]
  wire [7:0] _GEN_720 = 4'h1 == index ? quene_1 : quene_0; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_721 = 4'h2 == index ? quene_2 : _GEN_720; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_722 = 4'h3 == index ? quene_3 : _GEN_721; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_723 = 4'h4 == index ? quene_4 : _GEN_722; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_724 = 4'h5 == index ? quene_5 : _GEN_723; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_725 = 4'h6 == index ? quene_6 : _GEN_724; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_726 = 4'h7 == index ? quene_7 : _GEN_725; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_727 = 4'h8 == index ? quene_8 : _GEN_726; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_728 = 4'h9 == index ? quene_9 : _GEN_727; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_729 = 4'ha == index ? quene_10 : _GEN_728; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_730 = 4'hb == index ? quene_11 : _GEN_729; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_731 = 4'hc == index ? quene_12 : _GEN_730; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_732 = 4'hd == index ? quene_13 : _GEN_731; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_733 = 4'he == index ? quene_14 : _GEN_732; // @[d_cache.scala 173:{46,46}]
  wire [7:0] _GEN_734 = 4'hf == index ? quene_15 : _GEN_733; // @[d_cache.scala 173:{46,46}]
  wire [9:0] _GEN_5513 = {_GEN_734, 2'h0}; // @[d_cache.scala 173:46]
  wire [10:0] _quene_T = {{1'd0}, _GEN_5513}; // @[d_cache.scala 173:46]
  wire [7:0] _GEN_735 = 4'h0 == index ? _quene_T[7:0] : quene_0; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_736 = 4'h1 == index ? _quene_T[7:0] : quene_1; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_737 = 4'h2 == index ? _quene_T[7:0] : quene_2; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_738 = 4'h3 == index ? _quene_T[7:0] : quene_3; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_739 = 4'h4 == index ? _quene_T[7:0] : quene_4; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_740 = 4'h5 == index ? _quene_T[7:0] : quene_5; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_741 = 4'h6 == index ? _quene_T[7:0] : quene_6; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_742 = 4'h7 == index ? _quene_T[7:0] : quene_7; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_743 = 4'h8 == index ? _quene_T[7:0] : quene_8; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_744 = 4'h9 == index ? _quene_T[7:0] : quene_9; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_745 = 4'ha == index ? _quene_T[7:0] : quene_10; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_746 = 4'hb == index ? _quene_T[7:0] : quene_11; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_747 = 4'hc == index ? _quene_T[7:0] : quene_12; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_748 = 4'hd == index ? _quene_T[7:0] : quene_13; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_749 = 4'he == index ? _quene_T[7:0] : quene_14; // @[d_cache.scala 173:{30,30} 52:24]
  wire [7:0] _GEN_750 = 4'hf == index ? _quene_T[7:0] : quene_15; // @[d_cache.scala 173:{30,30} 52:24]
  wire [511:0] _GEN_751 = 4'h0 == index ? _ram_0_T_6 : ram_1_0; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_752 = 4'h1 == index ? _ram_0_T_6 : ram_1_1; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_753 = 4'h2 == index ? _ram_0_T_6 : ram_1_2; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_754 = 4'h3 == index ? _ram_0_T_6 : ram_1_3; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_755 = 4'h4 == index ? _ram_0_T_6 : ram_1_4; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_756 = 4'h5 == index ? _ram_0_T_6 : ram_1_5; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_757 = 4'h6 == index ? _ram_0_T_6 : ram_1_6; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_758 = 4'h7 == index ? _ram_0_T_6 : ram_1_7; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_759 = 4'h8 == index ? _ram_0_T_6 : ram_1_8; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_760 = 4'h9 == index ? _ram_0_T_6 : ram_1_9; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_761 = 4'ha == index ? _ram_0_T_6 : ram_1_10; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_762 = 4'hb == index ? _ram_0_T_6 : ram_1_11; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_763 = 4'hc == index ? _ram_0_T_6 : ram_1_12; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_764 = 4'hd == index ? _ram_0_T_6 : ram_1_13; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_765 = 4'he == index ? _ram_0_T_6 : ram_1_14; // @[d_cache.scala 176:{30,30} 20:24]
  wire [511:0] _GEN_766 = 4'hf == index ? _ram_0_T_6 : ram_1_15; // @[d_cache.scala 176:{30,30} 20:24]
  wire [31:0] _GEN_767 = 4'h0 == index ? _GEN_5341 : tag_1_0; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_768 = 4'h1 == index ? _GEN_5341 : tag_1_1; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_769 = 4'h2 == index ? _GEN_5341 : tag_1_2; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_770 = 4'h3 == index ? _GEN_5341 : tag_1_3; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_771 = 4'h4 == index ? _GEN_5341 : tag_1_4; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_772 = 4'h5 == index ? _GEN_5341 : tag_1_5; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_773 = 4'h6 == index ? _GEN_5341 : tag_1_6; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_774 = 4'h7 == index ? _GEN_5341 : tag_1_7; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_775 = 4'h8 == index ? _GEN_5341 : tag_1_8; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_776 = 4'h9 == index ? _GEN_5341 : tag_1_9; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_777 = 4'ha == index ? _GEN_5341 : tag_1_10; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_778 = 4'hb == index ? _GEN_5341 : tag_1_11; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_779 = 4'hc == index ? _GEN_5341 : tag_1_12; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_780 = 4'hd == index ? _GEN_5341 : tag_1_13; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_781 = 4'he == index ? _GEN_5341 : tag_1_14; // @[d_cache.scala 177:{30,30} 25:24]
  wire [31:0] _GEN_782 = 4'hf == index ? _GEN_5341 : tag_1_15; // @[d_cache.scala 177:{30,30} 25:24]
  wire  _GEN_783 = _GEN_5351 | valid_1_0; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_784 = _GEN_5356 | valid_1_1; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_785 = _GEN_5357 | valid_1_2; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_786 = _GEN_5361 | valid_1_3; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_787 = _GEN_5365 | valid_1_4; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_788 = _GEN_5367 | valid_1_5; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_789 = _GEN_5369 | valid_1_6; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_790 = _GEN_5370 | valid_1_7; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_791 = _GEN_5374 | valid_1_8; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_792 = _GEN_5375 | valid_1_9; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_793 = _GEN_5380 | valid_1_10; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_794 = _GEN_5381 | valid_1_11; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_795 = _GEN_5384 | valid_1_12; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_796 = _GEN_5388 | valid_1_13; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_797 = _GEN_5390 | valid_1_14; // @[d_cache.scala 178:{32,32} 30:26]
  wire  _GEN_798 = _GEN_5392 | valid_1_15; // @[d_cache.scala 178:{32,32} 30:26]
  wire [10:0] _quene_T_2 = _quene_T | 11'h1; // @[d_cache.scala 179:55]
  wire [7:0] _GEN_799 = 4'h0 == index ? _quene_T_2[7:0] : quene_0; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_800 = 4'h1 == index ? _quene_T_2[7:0] : quene_1; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_801 = 4'h2 == index ? _quene_T_2[7:0] : quene_2; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_802 = 4'h3 == index ? _quene_T_2[7:0] : quene_3; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_803 = 4'h4 == index ? _quene_T_2[7:0] : quene_4; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_804 = 4'h5 == index ? _quene_T_2[7:0] : quene_5; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_805 = 4'h6 == index ? _quene_T_2[7:0] : quene_6; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_806 = 4'h7 == index ? _quene_T_2[7:0] : quene_7; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_807 = 4'h8 == index ? _quene_T_2[7:0] : quene_8; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_808 = 4'h9 == index ? _quene_T_2[7:0] : quene_9; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_809 = 4'ha == index ? _quene_T_2[7:0] : quene_10; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_810 = 4'hb == index ? _quene_T_2[7:0] : quene_11; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_811 = 4'hc == index ? _quene_T_2[7:0] : quene_12; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_812 = 4'hd == index ? _quene_T_2[7:0] : quene_13; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_813 = 4'he == index ? _quene_T_2[7:0] : quene_14; // @[d_cache.scala 179:{30,30} 52:24]
  wire [7:0] _GEN_814 = 4'hf == index ? _quene_T_2[7:0] : quene_15; // @[d_cache.scala 179:{30,30} 52:24]
  wire [511:0] _GEN_815 = 4'h0 == index ? _ram_0_T_6 : ram_2_0; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_816 = 4'h1 == index ? _ram_0_T_6 : ram_2_1; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_817 = 4'h2 == index ? _ram_0_T_6 : ram_2_2; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_818 = 4'h3 == index ? _ram_0_T_6 : ram_2_3; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_819 = 4'h4 == index ? _ram_0_T_6 : ram_2_4; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_820 = 4'h5 == index ? _ram_0_T_6 : ram_2_5; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_821 = 4'h6 == index ? _ram_0_T_6 : ram_2_6; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_822 = 4'h7 == index ? _ram_0_T_6 : ram_2_7; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_823 = 4'h8 == index ? _ram_0_T_6 : ram_2_8; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_824 = 4'h9 == index ? _ram_0_T_6 : ram_2_9; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_825 = 4'ha == index ? _ram_0_T_6 : ram_2_10; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_826 = 4'hb == index ? _ram_0_T_6 : ram_2_11; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_827 = 4'hc == index ? _ram_0_T_6 : ram_2_12; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_828 = 4'hd == index ? _ram_0_T_6 : ram_2_13; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_829 = 4'he == index ? _ram_0_T_6 : ram_2_14; // @[d_cache.scala 182:{30,30} 21:24]
  wire [511:0] _GEN_830 = 4'hf == index ? _ram_0_T_6 : ram_2_15; // @[d_cache.scala 182:{30,30} 21:24]
  wire [31:0] _GEN_831 = 4'h0 == index ? _GEN_5341 : tag_2_0; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_832 = 4'h1 == index ? _GEN_5341 : tag_2_1; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_833 = 4'h2 == index ? _GEN_5341 : tag_2_2; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_834 = 4'h3 == index ? _GEN_5341 : tag_2_3; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_835 = 4'h4 == index ? _GEN_5341 : tag_2_4; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_836 = 4'h5 == index ? _GEN_5341 : tag_2_5; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_837 = 4'h6 == index ? _GEN_5341 : tag_2_6; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_838 = 4'h7 == index ? _GEN_5341 : tag_2_7; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_839 = 4'h8 == index ? _GEN_5341 : tag_2_8; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_840 = 4'h9 == index ? _GEN_5341 : tag_2_9; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_841 = 4'ha == index ? _GEN_5341 : tag_2_10; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_842 = 4'hb == index ? _GEN_5341 : tag_2_11; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_843 = 4'hc == index ? _GEN_5341 : tag_2_12; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_844 = 4'hd == index ? _GEN_5341 : tag_2_13; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_845 = 4'he == index ? _GEN_5341 : tag_2_14; // @[d_cache.scala 183:{30,30} 26:24]
  wire [31:0] _GEN_846 = 4'hf == index ? _GEN_5341 : tag_2_15; // @[d_cache.scala 183:{30,30} 26:24]
  wire  _GEN_847 = _GEN_5351 | valid_2_0; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_848 = _GEN_5356 | valid_2_1; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_849 = _GEN_5357 | valid_2_2; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_850 = _GEN_5361 | valid_2_3; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_851 = _GEN_5365 | valid_2_4; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_852 = _GEN_5367 | valid_2_5; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_853 = _GEN_5369 | valid_2_6; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_854 = _GEN_5370 | valid_2_7; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_855 = _GEN_5374 | valid_2_8; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_856 = _GEN_5375 | valid_2_9; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_857 = _GEN_5380 | valid_2_10; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_858 = _GEN_5381 | valid_2_11; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_859 = _GEN_5384 | valid_2_12; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_860 = _GEN_5388 | valid_2_13; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_861 = _GEN_5390 | valid_2_14; // @[d_cache.scala 184:{32,32} 31:26]
  wire  _GEN_862 = _GEN_5392 | valid_2_15; // @[d_cache.scala 184:{32,32} 31:26]
  wire [10:0] _quene_T_4 = _quene_T | 11'h2; // @[d_cache.scala 185:55]
  wire [7:0] _GEN_863 = 4'h0 == index ? _quene_T_4[7:0] : quene_0; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_864 = 4'h1 == index ? _quene_T_4[7:0] : quene_1; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_865 = 4'h2 == index ? _quene_T_4[7:0] : quene_2; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_866 = 4'h3 == index ? _quene_T_4[7:0] : quene_3; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_867 = 4'h4 == index ? _quene_T_4[7:0] : quene_4; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_868 = 4'h5 == index ? _quene_T_4[7:0] : quene_5; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_869 = 4'h6 == index ? _quene_T_4[7:0] : quene_6; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_870 = 4'h7 == index ? _quene_T_4[7:0] : quene_7; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_871 = 4'h8 == index ? _quene_T_4[7:0] : quene_8; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_872 = 4'h9 == index ? _quene_T_4[7:0] : quene_9; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_873 = 4'ha == index ? _quene_T_4[7:0] : quene_10; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_874 = 4'hb == index ? _quene_T_4[7:0] : quene_11; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_875 = 4'hc == index ? _quene_T_4[7:0] : quene_12; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_876 = 4'hd == index ? _quene_T_4[7:0] : quene_13; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_877 = 4'he == index ? _quene_T_4[7:0] : quene_14; // @[d_cache.scala 185:{30,30} 52:24]
  wire [7:0] _GEN_878 = 4'hf == index ? _quene_T_4[7:0] : quene_15; // @[d_cache.scala 185:{30,30} 52:24]
  wire [511:0] _GEN_879 = 4'h0 == index ? _ram_0_T_6 : ram_3_0; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_880 = 4'h1 == index ? _ram_0_T_6 : ram_3_1; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_881 = 4'h2 == index ? _ram_0_T_6 : ram_3_2; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_882 = 4'h3 == index ? _ram_0_T_6 : ram_3_3; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_883 = 4'h4 == index ? _ram_0_T_6 : ram_3_4; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_884 = 4'h5 == index ? _ram_0_T_6 : ram_3_5; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_885 = 4'h6 == index ? _ram_0_T_6 : ram_3_6; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_886 = 4'h7 == index ? _ram_0_T_6 : ram_3_7; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_887 = 4'h8 == index ? _ram_0_T_6 : ram_3_8; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_888 = 4'h9 == index ? _ram_0_T_6 : ram_3_9; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_889 = 4'ha == index ? _ram_0_T_6 : ram_3_10; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_890 = 4'hb == index ? _ram_0_T_6 : ram_3_11; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_891 = 4'hc == index ? _ram_0_T_6 : ram_3_12; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_892 = 4'hd == index ? _ram_0_T_6 : ram_3_13; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_893 = 4'he == index ? _ram_0_T_6 : ram_3_14; // @[d_cache.scala 188:{30,30} 22:24]
  wire [511:0] _GEN_894 = 4'hf == index ? _ram_0_T_6 : ram_3_15; // @[d_cache.scala 188:{30,30} 22:24]
  wire [31:0] _GEN_895 = 4'h0 == index ? _GEN_5341 : tag_3_0; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_896 = 4'h1 == index ? _GEN_5341 : tag_3_1; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_897 = 4'h2 == index ? _GEN_5341 : tag_3_2; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_898 = 4'h3 == index ? _GEN_5341 : tag_3_3; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_899 = 4'h4 == index ? _GEN_5341 : tag_3_4; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_900 = 4'h5 == index ? _GEN_5341 : tag_3_5; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_901 = 4'h6 == index ? _GEN_5341 : tag_3_6; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_902 = 4'h7 == index ? _GEN_5341 : tag_3_7; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_903 = 4'h8 == index ? _GEN_5341 : tag_3_8; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_904 = 4'h9 == index ? _GEN_5341 : tag_3_9; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_905 = 4'ha == index ? _GEN_5341 : tag_3_10; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_906 = 4'hb == index ? _GEN_5341 : tag_3_11; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_907 = 4'hc == index ? _GEN_5341 : tag_3_12; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_908 = 4'hd == index ? _GEN_5341 : tag_3_13; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_909 = 4'he == index ? _GEN_5341 : tag_3_14; // @[d_cache.scala 189:{30,30} 27:24]
  wire [31:0] _GEN_910 = 4'hf == index ? _GEN_5341 : tag_3_15; // @[d_cache.scala 189:{30,30} 27:24]
  wire  _GEN_911 = _GEN_5351 | valid_3_0; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_912 = _GEN_5356 | valid_3_1; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_913 = _GEN_5357 | valid_3_2; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_914 = _GEN_5361 | valid_3_3; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_915 = _GEN_5365 | valid_3_4; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_916 = _GEN_5367 | valid_3_5; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_917 = _GEN_5369 | valid_3_6; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_918 = _GEN_5370 | valid_3_7; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_919 = _GEN_5374 | valid_3_8; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_920 = _GEN_5375 | valid_3_9; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_921 = _GEN_5380 | valid_3_10; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_922 = _GEN_5381 | valid_3_11; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_923 = _GEN_5384 | valid_3_12; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_924 = _GEN_5388 | valid_3_13; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_925 = _GEN_5390 | valid_3_14; // @[d_cache.scala 190:{32,32} 32:26]
  wire  _GEN_926 = _GEN_5392 | valid_3_15; // @[d_cache.scala 190:{32,32} 32:26]
  wire [10:0] _quene_T_6 = _quene_T | 11'h3; // @[d_cache.scala 191:55]
  wire [7:0] _GEN_927 = 4'h0 == index ? _quene_T_6[7:0] : quene_0; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_928 = 4'h1 == index ? _quene_T_6[7:0] : quene_1; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_929 = 4'h2 == index ? _quene_T_6[7:0] : quene_2; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_930 = 4'h3 == index ? _quene_T_6[7:0] : quene_3; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_931 = 4'h4 == index ? _quene_T_6[7:0] : quene_4; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_932 = 4'h5 == index ? _quene_T_6[7:0] : quene_5; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_933 = 4'h6 == index ? _quene_T_6[7:0] : quene_6; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_934 = 4'h7 == index ? _quene_T_6[7:0] : quene_7; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_935 = 4'h8 == index ? _quene_T_6[7:0] : quene_8; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_936 = 4'h9 == index ? _quene_T_6[7:0] : quene_9; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_937 = 4'ha == index ? _quene_T_6[7:0] : quene_10; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_938 = 4'hb == index ? _quene_T_6[7:0] : quene_11; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_939 = 4'hc == index ? _quene_T_6[7:0] : quene_12; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_940 = 4'hd == index ? _quene_T_6[7:0] : quene_13; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_941 = 4'he == index ? _quene_T_6[7:0] : quene_14; // @[d_cache.scala 191:{30,30} 52:24]
  wire [7:0] _GEN_942 = 4'hf == index ? _quene_T_6[7:0] : quene_15; // @[d_cache.scala 191:{30,30} 52:24]
  wire  _GEN_944 = 4'h1 == index ? dirty_0_1 : dirty_0_0; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_945 = 4'h2 == index ? dirty_0_2 : _GEN_944; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_946 = 4'h3 == index ? dirty_0_3 : _GEN_945; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_947 = 4'h4 == index ? dirty_0_4 : _GEN_946; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_948 = 4'h5 == index ? dirty_0_5 : _GEN_947; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_949 = 4'h6 == index ? dirty_0_6 : _GEN_948; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_950 = 4'h7 == index ? dirty_0_7 : _GEN_949; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_951 = 4'h8 == index ? dirty_0_8 : _GEN_950; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_952 = 4'h9 == index ? dirty_0_9 : _GEN_951; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_953 = 4'ha == index ? dirty_0_10 : _GEN_952; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_954 = 4'hb == index ? dirty_0_11 : _GEN_953; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_955 = 4'hc == index ? dirty_0_12 : _GEN_954; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_956 = 4'hd == index ? dirty_0_13 : _GEN_955; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_957 = 4'he == index ? dirty_0_14 : _GEN_956; // @[d_cache.scala 194:{40,40}]
  wire  _GEN_958 = 4'hf == index ? dirty_0_15 : _GEN_957; // @[d_cache.scala 194:{40,40}]
  wire [41:0] _write_back_addr_T_1 = {_GEN_15,index,6'h0}; // @[Cat.scala 31:58]
  wire  _GEN_991 = 4'h0 == index ? 1'h0 : dirty_0_0; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_992 = 4'h1 == index ? 1'h0 : dirty_0_1; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_993 = 4'h2 == index ? 1'h0 : dirty_0_2; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_994 = 4'h3 == index ? 1'h0 : dirty_0_3; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_995 = 4'h4 == index ? 1'h0 : dirty_0_4; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_996 = 4'h5 == index ? 1'h0 : dirty_0_5; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_997 = 4'h6 == index ? 1'h0 : dirty_0_6; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_998 = 4'h7 == index ? 1'h0 : dirty_0_7; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_999 = 4'h8 == index ? 1'h0 : dirty_0_8; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_1000 = 4'h9 == index ? 1'h0 : dirty_0_9; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_1001 = 4'ha == index ? 1'h0 : dirty_0_10; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_1002 = 4'hb == index ? 1'h0 : dirty_0_11; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_1003 = 4'hc == index ? 1'h0 : dirty_0_12; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_1004 = 4'hd == index ? 1'h0 : dirty_0_13; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_1005 = 4'he == index ? 1'h0 : dirty_0_14; // @[d_cache.scala 199:{40,40} 34:26]
  wire  _GEN_1006 = 4'hf == index ? 1'h0 : dirty_0_15; // @[d_cache.scala 199:{40,40} 34:26]
  wire [511:0] _GEN_1103 = _GEN_958 ? _GEN_150 : write_back_data; // @[d_cache.scala 194:47 195:41 44:34]
  wire [41:0] _GEN_1104 = _GEN_958 ? _write_back_addr_T_1 : {{10'd0}, write_back_addr}; // @[d_cache.scala 194:47 196:41 45:34]
  wire [511:0] _GEN_1105 = _GEN_958 ? _GEN_671 : _GEN_671; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1106 = _GEN_958 ? _GEN_672 : _GEN_672; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1107 = _GEN_958 ? _GEN_673 : _GEN_673; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1108 = _GEN_958 ? _GEN_674 : _GEN_674; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1109 = _GEN_958 ? _GEN_675 : _GEN_675; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1110 = _GEN_958 ? _GEN_676 : _GEN_676; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1111 = _GEN_958 ? _GEN_677 : _GEN_677; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1112 = _GEN_958 ? _GEN_678 : _GEN_678; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1113 = _GEN_958 ? _GEN_679 : _GEN_679; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1114 = _GEN_958 ? _GEN_680 : _GEN_680; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1115 = _GEN_958 ? _GEN_681 : _GEN_681; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1116 = _GEN_958 ? _GEN_682 : _GEN_682; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1117 = _GEN_958 ? _GEN_683 : _GEN_683; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1118 = _GEN_958 ? _GEN_684 : _GEN_684; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1119 = _GEN_958 ? _GEN_685 : _GEN_685; // @[d_cache.scala 194:47]
  wire [511:0] _GEN_1120 = _GEN_958 ? _GEN_686 : _GEN_686; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1121 = _GEN_958 ? _GEN_687 : _GEN_687; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1122 = _GEN_958 ? _GEN_688 : _GEN_688; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1123 = _GEN_958 ? _GEN_689 : _GEN_689; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1124 = _GEN_958 ? _GEN_690 : _GEN_690; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1125 = _GEN_958 ? _GEN_691 : _GEN_691; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1126 = _GEN_958 ? _GEN_692 : _GEN_692; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1127 = _GEN_958 ? _GEN_693 : _GEN_693; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1128 = _GEN_958 ? _GEN_694 : _GEN_694; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1129 = _GEN_958 ? _GEN_695 : _GEN_695; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1130 = _GEN_958 ? _GEN_696 : _GEN_696; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1131 = _GEN_958 ? _GEN_697 : _GEN_697; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1132 = _GEN_958 ? _GEN_698 : _GEN_698; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1133 = _GEN_958 ? _GEN_699 : _GEN_699; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1134 = _GEN_958 ? _GEN_700 : _GEN_700; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1135 = _GEN_958 ? _GEN_701 : _GEN_701; // @[d_cache.scala 194:47]
  wire [31:0] _GEN_1136 = _GEN_958 ? _GEN_702 : _GEN_702; // @[d_cache.scala 194:47]
  wire  _GEN_1137 = _GEN_958 ? _GEN_991 : dirty_0_0; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1138 = _GEN_958 ? _GEN_992 : dirty_0_1; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1139 = _GEN_958 ? _GEN_993 : dirty_0_2; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1140 = _GEN_958 ? _GEN_994 : dirty_0_3; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1141 = _GEN_958 ? _GEN_995 : dirty_0_4; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1142 = _GEN_958 ? _GEN_996 : dirty_0_5; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1143 = _GEN_958 ? _GEN_997 : dirty_0_6; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1144 = _GEN_958 ? _GEN_998 : dirty_0_7; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1145 = _GEN_958 ? _GEN_999 : dirty_0_8; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1146 = _GEN_958 ? _GEN_1000 : dirty_0_9; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1147 = _GEN_958 ? _GEN_1001 : dirty_0_10; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1148 = _GEN_958 ? _GEN_1002 : dirty_0_11; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1149 = _GEN_958 ? _GEN_1003 : dirty_0_12; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1150 = _GEN_958 ? _GEN_1004 : dirty_0_13; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1151 = _GEN_958 ? _GEN_1005 : dirty_0_14; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1152 = _GEN_958 ? _GEN_1006 : dirty_0_15; // @[d_cache.scala 194:47 34:26]
  wire  _GEN_1153 = _GEN_958 ? _GEN_703 : _GEN_703; // @[d_cache.scala 194:47]
  wire  _GEN_1154 = _GEN_958 ? _GEN_704 : _GEN_704; // @[d_cache.scala 194:47]
  wire  _GEN_1155 = _GEN_958 ? _GEN_705 : _GEN_705; // @[d_cache.scala 194:47]
  wire  _GEN_1156 = _GEN_958 ? _GEN_706 : _GEN_706; // @[d_cache.scala 194:47]
  wire  _GEN_1157 = _GEN_958 ? _GEN_707 : _GEN_707; // @[d_cache.scala 194:47]
  wire  _GEN_1158 = _GEN_958 ? _GEN_708 : _GEN_708; // @[d_cache.scala 194:47]
  wire  _GEN_1159 = _GEN_958 ? _GEN_709 : _GEN_709; // @[d_cache.scala 194:47]
  wire  _GEN_1160 = _GEN_958 ? _GEN_710 : _GEN_710; // @[d_cache.scala 194:47]
  wire  _GEN_1161 = _GEN_958 ? _GEN_711 : _GEN_711; // @[d_cache.scala 194:47]
  wire  _GEN_1162 = _GEN_958 ? _GEN_712 : _GEN_712; // @[d_cache.scala 194:47]
  wire  _GEN_1163 = _GEN_958 ? _GEN_713 : _GEN_713; // @[d_cache.scala 194:47]
  wire  _GEN_1164 = _GEN_958 ? _GEN_714 : _GEN_714; // @[d_cache.scala 194:47]
  wire  _GEN_1165 = _GEN_958 ? _GEN_715 : _GEN_715; // @[d_cache.scala 194:47]
  wire  _GEN_1166 = _GEN_958 ? _GEN_716 : _GEN_716; // @[d_cache.scala 194:47]
  wire  _GEN_1167 = _GEN_958 ? _GEN_717 : _GEN_717; // @[d_cache.scala 194:47]
  wire  _GEN_1168 = _GEN_958 ? _GEN_718 : _GEN_718; // @[d_cache.scala 194:47]
  wire [3:0] _GEN_1169 = _GEN_958 ? 4'h6 : 4'h1; // @[d_cache.scala 194:47 201:31 204:31]
  wire [7:0] _GEN_1170 = _GEN_958 ? _GEN_735 : _GEN_735; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1171 = _GEN_958 ? _GEN_736 : _GEN_736; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1172 = _GEN_958 ? _GEN_737 : _GEN_737; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1173 = _GEN_958 ? _GEN_738 : _GEN_738; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1174 = _GEN_958 ? _GEN_739 : _GEN_739; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1175 = _GEN_958 ? _GEN_740 : _GEN_740; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1176 = _GEN_958 ? _GEN_741 : _GEN_741; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1177 = _GEN_958 ? _GEN_742 : _GEN_742; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1178 = _GEN_958 ? _GEN_743 : _GEN_743; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1179 = _GEN_958 ? _GEN_744 : _GEN_744; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1180 = _GEN_958 ? _GEN_745 : _GEN_745; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1181 = _GEN_958 ? _GEN_746 : _GEN_746; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1182 = _GEN_958 ? _GEN_747 : _GEN_747; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1183 = _GEN_958 ? _GEN_748 : _GEN_748; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1184 = _GEN_958 ? _GEN_749 : _GEN_749; // @[d_cache.scala 194:47]
  wire [7:0] _GEN_1185 = _GEN_958 ? _GEN_750 : _GEN_750; // @[d_cache.scala 194:47]
  wire  _GEN_1187 = 4'h1 == index ? dirty_1_1 : dirty_1_0; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1188 = 4'h2 == index ? dirty_1_2 : _GEN_1187; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1189 = 4'h3 == index ? dirty_1_3 : _GEN_1188; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1190 = 4'h4 == index ? dirty_1_4 : _GEN_1189; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1191 = 4'h5 == index ? dirty_1_5 : _GEN_1190; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1192 = 4'h6 == index ? dirty_1_6 : _GEN_1191; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1193 = 4'h7 == index ? dirty_1_7 : _GEN_1192; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1194 = 4'h8 == index ? dirty_1_8 : _GEN_1193; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1195 = 4'h9 == index ? dirty_1_9 : _GEN_1194; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1196 = 4'ha == index ? dirty_1_10 : _GEN_1195; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1197 = 4'hb == index ? dirty_1_11 : _GEN_1196; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1198 = 4'hc == index ? dirty_1_12 : _GEN_1197; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1199 = 4'hd == index ? dirty_1_13 : _GEN_1198; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1200 = 4'he == index ? dirty_1_14 : _GEN_1199; // @[d_cache.scala 211:{40,40}]
  wire  _GEN_1201 = 4'hf == index ? dirty_1_15 : _GEN_1200; // @[d_cache.scala 211:{40,40}]
  wire [41:0] _write_back_addr_T_3 = {_GEN_47,index,6'h0}; // @[Cat.scala 31:58]
  wire  _GEN_1234 = 4'h0 == index ? 1'h0 : dirty_1_0; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1235 = 4'h1 == index ? 1'h0 : dirty_1_1; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1236 = 4'h2 == index ? 1'h0 : dirty_1_2; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1237 = 4'h3 == index ? 1'h0 : dirty_1_3; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1238 = 4'h4 == index ? 1'h0 : dirty_1_4; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1239 = 4'h5 == index ? 1'h0 : dirty_1_5; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1240 = 4'h6 == index ? 1'h0 : dirty_1_6; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1241 = 4'h7 == index ? 1'h0 : dirty_1_7; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1242 = 4'h8 == index ? 1'h0 : dirty_1_8; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1243 = 4'h9 == index ? 1'h0 : dirty_1_9; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1244 = 4'ha == index ? 1'h0 : dirty_1_10; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1245 = 4'hb == index ? 1'h0 : dirty_1_11; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1246 = 4'hc == index ? 1'h0 : dirty_1_12; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1247 = 4'hd == index ? 1'h0 : dirty_1_13; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1248 = 4'he == index ? 1'h0 : dirty_1_14; // @[d_cache.scala 216:{40,40} 35:26]
  wire  _GEN_1249 = 4'hf == index ? 1'h0 : dirty_1_15; // @[d_cache.scala 216:{40,40} 35:26]
  wire [511:0] _GEN_1346 = _GEN_1201 ? _GEN_198 : write_back_data; // @[d_cache.scala 211:47 212:41 44:34]
  wire [41:0] _GEN_1347 = _GEN_1201 ? _write_back_addr_T_3 : {{10'd0}, write_back_addr}; // @[d_cache.scala 211:47 213:41 45:34]
  wire [511:0] _GEN_1348 = _GEN_1201 ? _GEN_751 : _GEN_751; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1349 = _GEN_1201 ? _GEN_752 : _GEN_752; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1350 = _GEN_1201 ? _GEN_753 : _GEN_753; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1351 = _GEN_1201 ? _GEN_754 : _GEN_754; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1352 = _GEN_1201 ? _GEN_755 : _GEN_755; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1353 = _GEN_1201 ? _GEN_756 : _GEN_756; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1354 = _GEN_1201 ? _GEN_757 : _GEN_757; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1355 = _GEN_1201 ? _GEN_758 : _GEN_758; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1356 = _GEN_1201 ? _GEN_759 : _GEN_759; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1357 = _GEN_1201 ? _GEN_760 : _GEN_760; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1358 = _GEN_1201 ? _GEN_761 : _GEN_761; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1359 = _GEN_1201 ? _GEN_762 : _GEN_762; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1360 = _GEN_1201 ? _GEN_763 : _GEN_763; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1361 = _GEN_1201 ? _GEN_764 : _GEN_764; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1362 = _GEN_1201 ? _GEN_765 : _GEN_765; // @[d_cache.scala 211:47]
  wire [511:0] _GEN_1363 = _GEN_1201 ? _GEN_766 : _GEN_766; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1364 = _GEN_1201 ? _GEN_767 : _GEN_767; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1365 = _GEN_1201 ? _GEN_768 : _GEN_768; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1366 = _GEN_1201 ? _GEN_769 : _GEN_769; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1367 = _GEN_1201 ? _GEN_770 : _GEN_770; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1368 = _GEN_1201 ? _GEN_771 : _GEN_771; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1369 = _GEN_1201 ? _GEN_772 : _GEN_772; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1370 = _GEN_1201 ? _GEN_773 : _GEN_773; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1371 = _GEN_1201 ? _GEN_774 : _GEN_774; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1372 = _GEN_1201 ? _GEN_775 : _GEN_775; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1373 = _GEN_1201 ? _GEN_776 : _GEN_776; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1374 = _GEN_1201 ? _GEN_777 : _GEN_777; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1375 = _GEN_1201 ? _GEN_778 : _GEN_778; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1376 = _GEN_1201 ? _GEN_779 : _GEN_779; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1377 = _GEN_1201 ? _GEN_780 : _GEN_780; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1378 = _GEN_1201 ? _GEN_781 : _GEN_781; // @[d_cache.scala 211:47]
  wire [31:0] _GEN_1379 = _GEN_1201 ? _GEN_782 : _GEN_782; // @[d_cache.scala 211:47]
  wire  _GEN_1380 = _GEN_1201 ? _GEN_1234 : dirty_1_0; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1381 = _GEN_1201 ? _GEN_1235 : dirty_1_1; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1382 = _GEN_1201 ? _GEN_1236 : dirty_1_2; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1383 = _GEN_1201 ? _GEN_1237 : dirty_1_3; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1384 = _GEN_1201 ? _GEN_1238 : dirty_1_4; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1385 = _GEN_1201 ? _GEN_1239 : dirty_1_5; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1386 = _GEN_1201 ? _GEN_1240 : dirty_1_6; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1387 = _GEN_1201 ? _GEN_1241 : dirty_1_7; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1388 = _GEN_1201 ? _GEN_1242 : dirty_1_8; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1389 = _GEN_1201 ? _GEN_1243 : dirty_1_9; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1390 = _GEN_1201 ? _GEN_1244 : dirty_1_10; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1391 = _GEN_1201 ? _GEN_1245 : dirty_1_11; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1392 = _GEN_1201 ? _GEN_1246 : dirty_1_12; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1393 = _GEN_1201 ? _GEN_1247 : dirty_1_13; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1394 = _GEN_1201 ? _GEN_1248 : dirty_1_14; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1395 = _GEN_1201 ? _GEN_1249 : dirty_1_15; // @[d_cache.scala 211:47 35:26]
  wire  _GEN_1396 = _GEN_1201 ? _GEN_783 : _GEN_783; // @[d_cache.scala 211:47]
  wire  _GEN_1397 = _GEN_1201 ? _GEN_784 : _GEN_784; // @[d_cache.scala 211:47]
  wire  _GEN_1398 = _GEN_1201 ? _GEN_785 : _GEN_785; // @[d_cache.scala 211:47]
  wire  _GEN_1399 = _GEN_1201 ? _GEN_786 : _GEN_786; // @[d_cache.scala 211:47]
  wire  _GEN_1400 = _GEN_1201 ? _GEN_787 : _GEN_787; // @[d_cache.scala 211:47]
  wire  _GEN_1401 = _GEN_1201 ? _GEN_788 : _GEN_788; // @[d_cache.scala 211:47]
  wire  _GEN_1402 = _GEN_1201 ? _GEN_789 : _GEN_789; // @[d_cache.scala 211:47]
  wire  _GEN_1403 = _GEN_1201 ? _GEN_790 : _GEN_790; // @[d_cache.scala 211:47]
  wire  _GEN_1404 = _GEN_1201 ? _GEN_791 : _GEN_791; // @[d_cache.scala 211:47]
  wire  _GEN_1405 = _GEN_1201 ? _GEN_792 : _GEN_792; // @[d_cache.scala 211:47]
  wire  _GEN_1406 = _GEN_1201 ? _GEN_793 : _GEN_793; // @[d_cache.scala 211:47]
  wire  _GEN_1407 = _GEN_1201 ? _GEN_794 : _GEN_794; // @[d_cache.scala 211:47]
  wire  _GEN_1408 = _GEN_1201 ? _GEN_795 : _GEN_795; // @[d_cache.scala 211:47]
  wire  _GEN_1409 = _GEN_1201 ? _GEN_796 : _GEN_796; // @[d_cache.scala 211:47]
  wire  _GEN_1410 = _GEN_1201 ? _GEN_797 : _GEN_797; // @[d_cache.scala 211:47]
  wire  _GEN_1411 = _GEN_1201 ? _GEN_798 : _GEN_798; // @[d_cache.scala 211:47]
  wire [3:0] _GEN_1412 = _GEN_1201 ? 4'h6 : 4'h1; // @[d_cache.scala 211:47 218:31 221:31]
  wire [7:0] _GEN_1413 = _GEN_1201 ? _GEN_799 : _GEN_799; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1414 = _GEN_1201 ? _GEN_800 : _GEN_800; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1415 = _GEN_1201 ? _GEN_801 : _GEN_801; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1416 = _GEN_1201 ? _GEN_802 : _GEN_802; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1417 = _GEN_1201 ? _GEN_803 : _GEN_803; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1418 = _GEN_1201 ? _GEN_804 : _GEN_804; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1419 = _GEN_1201 ? _GEN_805 : _GEN_805; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1420 = _GEN_1201 ? _GEN_806 : _GEN_806; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1421 = _GEN_1201 ? _GEN_807 : _GEN_807; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1422 = _GEN_1201 ? _GEN_808 : _GEN_808; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1423 = _GEN_1201 ? _GEN_809 : _GEN_809; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1424 = _GEN_1201 ? _GEN_810 : _GEN_810; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1425 = _GEN_1201 ? _GEN_811 : _GEN_811; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1426 = _GEN_1201 ? _GEN_812 : _GEN_812; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1427 = _GEN_1201 ? _GEN_813 : _GEN_813; // @[d_cache.scala 211:47]
  wire [7:0] _GEN_1428 = _GEN_1201 ? _GEN_814 : _GEN_814; // @[d_cache.scala 211:47]
  wire  _GEN_1430 = 4'h1 == index ? dirty_2_1 : dirty_2_0; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1431 = 4'h2 == index ? dirty_2_2 : _GEN_1430; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1432 = 4'h3 == index ? dirty_2_3 : _GEN_1431; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1433 = 4'h4 == index ? dirty_2_4 : _GEN_1432; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1434 = 4'h5 == index ? dirty_2_5 : _GEN_1433; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1435 = 4'h6 == index ? dirty_2_6 : _GEN_1434; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1436 = 4'h7 == index ? dirty_2_7 : _GEN_1435; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1437 = 4'h8 == index ? dirty_2_8 : _GEN_1436; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1438 = 4'h9 == index ? dirty_2_9 : _GEN_1437; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1439 = 4'ha == index ? dirty_2_10 : _GEN_1438; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1440 = 4'hb == index ? dirty_2_11 : _GEN_1439; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1441 = 4'hc == index ? dirty_2_12 : _GEN_1440; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1442 = 4'hd == index ? dirty_2_13 : _GEN_1441; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1443 = 4'he == index ? dirty_2_14 : _GEN_1442; // @[d_cache.scala 228:{40,40}]
  wire  _GEN_1444 = 4'hf == index ? dirty_2_15 : _GEN_1443; // @[d_cache.scala 228:{40,40}]
  wire [41:0] _write_back_addr_T_5 = {_GEN_79,index,6'h0}; // @[Cat.scala 31:58]
  wire  _GEN_1477 = 4'h0 == index ? 1'h0 : dirty_2_0; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1478 = 4'h1 == index ? 1'h0 : dirty_2_1; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1479 = 4'h2 == index ? 1'h0 : dirty_2_2; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1480 = 4'h3 == index ? 1'h0 : dirty_2_3; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1481 = 4'h4 == index ? 1'h0 : dirty_2_4; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1482 = 4'h5 == index ? 1'h0 : dirty_2_5; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1483 = 4'h6 == index ? 1'h0 : dirty_2_6; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1484 = 4'h7 == index ? 1'h0 : dirty_2_7; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1485 = 4'h8 == index ? 1'h0 : dirty_2_8; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1486 = 4'h9 == index ? 1'h0 : dirty_2_9; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1487 = 4'ha == index ? 1'h0 : dirty_2_10; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1488 = 4'hb == index ? 1'h0 : dirty_2_11; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1489 = 4'hc == index ? 1'h0 : dirty_2_12; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1490 = 4'hd == index ? 1'h0 : dirty_2_13; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1491 = 4'he == index ? 1'h0 : dirty_2_14; // @[d_cache.scala 233:{40,40} 36:26]
  wire  _GEN_1492 = 4'hf == index ? 1'h0 : dirty_2_15; // @[d_cache.scala 233:{40,40} 36:26]
  wire [511:0] _GEN_1589 = _GEN_1444 ? _GEN_246 : write_back_data; // @[d_cache.scala 228:47 229:41 44:34]
  wire [41:0] _GEN_1590 = _GEN_1444 ? _write_back_addr_T_5 : {{10'd0}, write_back_addr}; // @[d_cache.scala 228:47 230:41 45:34]
  wire [511:0] _GEN_1591 = _GEN_1444 ? _GEN_815 : _GEN_815; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1592 = _GEN_1444 ? _GEN_816 : _GEN_816; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1593 = _GEN_1444 ? _GEN_817 : _GEN_817; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1594 = _GEN_1444 ? _GEN_818 : _GEN_818; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1595 = _GEN_1444 ? _GEN_819 : _GEN_819; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1596 = _GEN_1444 ? _GEN_820 : _GEN_820; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1597 = _GEN_1444 ? _GEN_821 : _GEN_821; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1598 = _GEN_1444 ? _GEN_822 : _GEN_822; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1599 = _GEN_1444 ? _GEN_823 : _GEN_823; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1600 = _GEN_1444 ? _GEN_824 : _GEN_824; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1601 = _GEN_1444 ? _GEN_825 : _GEN_825; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1602 = _GEN_1444 ? _GEN_826 : _GEN_826; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1603 = _GEN_1444 ? _GEN_827 : _GEN_827; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1604 = _GEN_1444 ? _GEN_828 : _GEN_828; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1605 = _GEN_1444 ? _GEN_829 : _GEN_829; // @[d_cache.scala 228:47]
  wire [511:0] _GEN_1606 = _GEN_1444 ? _GEN_830 : _GEN_830; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1607 = _GEN_1444 ? _GEN_831 : _GEN_831; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1608 = _GEN_1444 ? _GEN_832 : _GEN_832; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1609 = _GEN_1444 ? _GEN_833 : _GEN_833; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1610 = _GEN_1444 ? _GEN_834 : _GEN_834; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1611 = _GEN_1444 ? _GEN_835 : _GEN_835; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1612 = _GEN_1444 ? _GEN_836 : _GEN_836; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1613 = _GEN_1444 ? _GEN_837 : _GEN_837; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1614 = _GEN_1444 ? _GEN_838 : _GEN_838; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1615 = _GEN_1444 ? _GEN_839 : _GEN_839; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1616 = _GEN_1444 ? _GEN_840 : _GEN_840; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1617 = _GEN_1444 ? _GEN_841 : _GEN_841; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1618 = _GEN_1444 ? _GEN_842 : _GEN_842; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1619 = _GEN_1444 ? _GEN_843 : _GEN_843; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1620 = _GEN_1444 ? _GEN_844 : _GEN_844; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1621 = _GEN_1444 ? _GEN_845 : _GEN_845; // @[d_cache.scala 228:47]
  wire [31:0] _GEN_1622 = _GEN_1444 ? _GEN_846 : _GEN_846; // @[d_cache.scala 228:47]
  wire  _GEN_1623 = _GEN_1444 ? _GEN_1477 : dirty_2_0; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1624 = _GEN_1444 ? _GEN_1478 : dirty_2_1; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1625 = _GEN_1444 ? _GEN_1479 : dirty_2_2; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1626 = _GEN_1444 ? _GEN_1480 : dirty_2_3; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1627 = _GEN_1444 ? _GEN_1481 : dirty_2_4; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1628 = _GEN_1444 ? _GEN_1482 : dirty_2_5; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1629 = _GEN_1444 ? _GEN_1483 : dirty_2_6; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1630 = _GEN_1444 ? _GEN_1484 : dirty_2_7; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1631 = _GEN_1444 ? _GEN_1485 : dirty_2_8; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1632 = _GEN_1444 ? _GEN_1486 : dirty_2_9; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1633 = _GEN_1444 ? _GEN_1487 : dirty_2_10; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1634 = _GEN_1444 ? _GEN_1488 : dirty_2_11; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1635 = _GEN_1444 ? _GEN_1489 : dirty_2_12; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1636 = _GEN_1444 ? _GEN_1490 : dirty_2_13; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1637 = _GEN_1444 ? _GEN_1491 : dirty_2_14; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1638 = _GEN_1444 ? _GEN_1492 : dirty_2_15; // @[d_cache.scala 228:47 36:26]
  wire  _GEN_1639 = _GEN_1444 ? _GEN_847 : _GEN_847; // @[d_cache.scala 228:47]
  wire  _GEN_1640 = _GEN_1444 ? _GEN_848 : _GEN_848; // @[d_cache.scala 228:47]
  wire  _GEN_1641 = _GEN_1444 ? _GEN_849 : _GEN_849; // @[d_cache.scala 228:47]
  wire  _GEN_1642 = _GEN_1444 ? _GEN_850 : _GEN_850; // @[d_cache.scala 228:47]
  wire  _GEN_1643 = _GEN_1444 ? _GEN_851 : _GEN_851; // @[d_cache.scala 228:47]
  wire  _GEN_1644 = _GEN_1444 ? _GEN_852 : _GEN_852; // @[d_cache.scala 228:47]
  wire  _GEN_1645 = _GEN_1444 ? _GEN_853 : _GEN_853; // @[d_cache.scala 228:47]
  wire  _GEN_1646 = _GEN_1444 ? _GEN_854 : _GEN_854; // @[d_cache.scala 228:47]
  wire  _GEN_1647 = _GEN_1444 ? _GEN_855 : _GEN_855; // @[d_cache.scala 228:47]
  wire  _GEN_1648 = _GEN_1444 ? _GEN_856 : _GEN_856; // @[d_cache.scala 228:47]
  wire  _GEN_1649 = _GEN_1444 ? _GEN_857 : _GEN_857; // @[d_cache.scala 228:47]
  wire  _GEN_1650 = _GEN_1444 ? _GEN_858 : _GEN_858; // @[d_cache.scala 228:47]
  wire  _GEN_1651 = _GEN_1444 ? _GEN_859 : _GEN_859; // @[d_cache.scala 228:47]
  wire  _GEN_1652 = _GEN_1444 ? _GEN_860 : _GEN_860; // @[d_cache.scala 228:47]
  wire  _GEN_1653 = _GEN_1444 ? _GEN_861 : _GEN_861; // @[d_cache.scala 228:47]
  wire  _GEN_1654 = _GEN_1444 ? _GEN_862 : _GEN_862; // @[d_cache.scala 228:47]
  wire [3:0] _GEN_1655 = _GEN_1444 ? 4'h6 : 4'h1; // @[d_cache.scala 228:47 235:31 238:31]
  wire [7:0] _GEN_1656 = _GEN_1444 ? _GEN_863 : _GEN_863; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1657 = _GEN_1444 ? _GEN_864 : _GEN_864; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1658 = _GEN_1444 ? _GEN_865 : _GEN_865; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1659 = _GEN_1444 ? _GEN_866 : _GEN_866; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1660 = _GEN_1444 ? _GEN_867 : _GEN_867; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1661 = _GEN_1444 ? _GEN_868 : _GEN_868; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1662 = _GEN_1444 ? _GEN_869 : _GEN_869; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1663 = _GEN_1444 ? _GEN_870 : _GEN_870; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1664 = _GEN_1444 ? _GEN_871 : _GEN_871; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1665 = _GEN_1444 ? _GEN_872 : _GEN_872; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1666 = _GEN_1444 ? _GEN_873 : _GEN_873; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1667 = _GEN_1444 ? _GEN_874 : _GEN_874; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1668 = _GEN_1444 ? _GEN_875 : _GEN_875; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1669 = _GEN_1444 ? _GEN_876 : _GEN_876; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1670 = _GEN_1444 ? _GEN_877 : _GEN_877; // @[d_cache.scala 228:47]
  wire [7:0] _GEN_1671 = _GEN_1444 ? _GEN_878 : _GEN_878; // @[d_cache.scala 228:47]
  wire  _GEN_1673 = 4'h1 == index ? dirty_3_1 : dirty_3_0; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1674 = 4'h2 == index ? dirty_3_2 : _GEN_1673; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1675 = 4'h3 == index ? dirty_3_3 : _GEN_1674; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1676 = 4'h4 == index ? dirty_3_4 : _GEN_1675; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1677 = 4'h5 == index ? dirty_3_5 : _GEN_1676; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1678 = 4'h6 == index ? dirty_3_6 : _GEN_1677; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1679 = 4'h7 == index ? dirty_3_7 : _GEN_1678; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1680 = 4'h8 == index ? dirty_3_8 : _GEN_1679; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1681 = 4'h9 == index ? dirty_3_9 : _GEN_1680; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1682 = 4'ha == index ? dirty_3_10 : _GEN_1681; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1683 = 4'hb == index ? dirty_3_11 : _GEN_1682; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1684 = 4'hc == index ? dirty_3_12 : _GEN_1683; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1685 = 4'hd == index ? dirty_3_13 : _GEN_1684; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1686 = 4'he == index ? dirty_3_14 : _GEN_1685; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1687 = 4'hf == index ? dirty_3_15 : _GEN_1686; // @[d_cache.scala 245:{40,40}]
  wire  _GEN_1720 = 4'h0 == index ? 1'h0 : dirty_3_0; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1721 = 4'h1 == index ? 1'h0 : dirty_3_1; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1722 = 4'h2 == index ? 1'h0 : dirty_3_2; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1723 = 4'h3 == index ? 1'h0 : dirty_3_3; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1724 = 4'h4 == index ? 1'h0 : dirty_3_4; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1725 = 4'h5 == index ? 1'h0 : dirty_3_5; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1726 = 4'h6 == index ? 1'h0 : dirty_3_6; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1727 = 4'h7 == index ? 1'h0 : dirty_3_7; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1728 = 4'h8 == index ? 1'h0 : dirty_3_8; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1729 = 4'h9 == index ? 1'h0 : dirty_3_9; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1730 = 4'ha == index ? 1'h0 : dirty_3_10; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1731 = 4'hb == index ? 1'h0 : dirty_3_11; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1732 = 4'hc == index ? 1'h0 : dirty_3_12; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1733 = 4'hd == index ? 1'h0 : dirty_3_13; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1734 = 4'he == index ? 1'h0 : dirty_3_14; // @[d_cache.scala 250:{40,40} 37:26]
  wire  _GEN_1735 = 4'hf == index ? 1'h0 : dirty_3_15; // @[d_cache.scala 250:{40,40} 37:26]
  wire [511:0] _GEN_1832 = _GEN_1687 ? _GEN_294 : write_back_data; // @[d_cache.scala 245:47 246:41 44:34]
  wire [41:0] _GEN_1833 = _GEN_1687 ? _write_back_addr_T_3 : {{10'd0}, write_back_addr}; // @[d_cache.scala 245:47 247:41 45:34]
  wire [511:0] _GEN_1834 = _GEN_1687 ? _GEN_879 : _GEN_879; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1835 = _GEN_1687 ? _GEN_880 : _GEN_880; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1836 = _GEN_1687 ? _GEN_881 : _GEN_881; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1837 = _GEN_1687 ? _GEN_882 : _GEN_882; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1838 = _GEN_1687 ? _GEN_883 : _GEN_883; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1839 = _GEN_1687 ? _GEN_884 : _GEN_884; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1840 = _GEN_1687 ? _GEN_885 : _GEN_885; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1841 = _GEN_1687 ? _GEN_886 : _GEN_886; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1842 = _GEN_1687 ? _GEN_887 : _GEN_887; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1843 = _GEN_1687 ? _GEN_888 : _GEN_888; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1844 = _GEN_1687 ? _GEN_889 : _GEN_889; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1845 = _GEN_1687 ? _GEN_890 : _GEN_890; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1846 = _GEN_1687 ? _GEN_891 : _GEN_891; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1847 = _GEN_1687 ? _GEN_892 : _GEN_892; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1848 = _GEN_1687 ? _GEN_893 : _GEN_893; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1849 = _GEN_1687 ? _GEN_894 : _GEN_894; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1850 = _GEN_1687 ? _GEN_895 : _GEN_895; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1851 = _GEN_1687 ? _GEN_896 : _GEN_896; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1852 = _GEN_1687 ? _GEN_897 : _GEN_897; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1853 = _GEN_1687 ? _GEN_898 : _GEN_898; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1854 = _GEN_1687 ? _GEN_899 : _GEN_899; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1855 = _GEN_1687 ? _GEN_900 : _GEN_900; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1856 = _GEN_1687 ? _GEN_901 : _GEN_901; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1857 = _GEN_1687 ? _GEN_902 : _GEN_902; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1858 = _GEN_1687 ? _GEN_903 : _GEN_903; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1859 = _GEN_1687 ? _GEN_904 : _GEN_904; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1860 = _GEN_1687 ? _GEN_905 : _GEN_905; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1861 = _GEN_1687 ? _GEN_906 : _GEN_906; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1862 = _GEN_1687 ? _GEN_907 : _GEN_907; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1863 = _GEN_1687 ? _GEN_908 : _GEN_908; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1864 = _GEN_1687 ? _GEN_909 : _GEN_909; // @[d_cache.scala 245:47]
  wire [31:0] _GEN_1865 = _GEN_1687 ? _GEN_910 : _GEN_910; // @[d_cache.scala 245:47]
  wire  _GEN_1866 = _GEN_1687 ? _GEN_1720 : dirty_3_0; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1867 = _GEN_1687 ? _GEN_1721 : dirty_3_1; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1868 = _GEN_1687 ? _GEN_1722 : dirty_3_2; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1869 = _GEN_1687 ? _GEN_1723 : dirty_3_3; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1870 = _GEN_1687 ? _GEN_1724 : dirty_3_4; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1871 = _GEN_1687 ? _GEN_1725 : dirty_3_5; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1872 = _GEN_1687 ? _GEN_1726 : dirty_3_6; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1873 = _GEN_1687 ? _GEN_1727 : dirty_3_7; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1874 = _GEN_1687 ? _GEN_1728 : dirty_3_8; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1875 = _GEN_1687 ? _GEN_1729 : dirty_3_9; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1876 = _GEN_1687 ? _GEN_1730 : dirty_3_10; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1877 = _GEN_1687 ? _GEN_1731 : dirty_3_11; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1878 = _GEN_1687 ? _GEN_1732 : dirty_3_12; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1879 = _GEN_1687 ? _GEN_1733 : dirty_3_13; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1880 = _GEN_1687 ? _GEN_1734 : dirty_3_14; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1881 = _GEN_1687 ? _GEN_1735 : dirty_3_15; // @[d_cache.scala 245:47 37:26]
  wire  _GEN_1882 = _GEN_1687 ? _GEN_911 : _GEN_911; // @[d_cache.scala 245:47]
  wire  _GEN_1883 = _GEN_1687 ? _GEN_912 : _GEN_912; // @[d_cache.scala 245:47]
  wire  _GEN_1884 = _GEN_1687 ? _GEN_913 : _GEN_913; // @[d_cache.scala 245:47]
  wire  _GEN_1885 = _GEN_1687 ? _GEN_914 : _GEN_914; // @[d_cache.scala 245:47]
  wire  _GEN_1886 = _GEN_1687 ? _GEN_915 : _GEN_915; // @[d_cache.scala 245:47]
  wire  _GEN_1887 = _GEN_1687 ? _GEN_916 : _GEN_916; // @[d_cache.scala 245:47]
  wire  _GEN_1888 = _GEN_1687 ? _GEN_917 : _GEN_917; // @[d_cache.scala 245:47]
  wire  _GEN_1889 = _GEN_1687 ? _GEN_918 : _GEN_918; // @[d_cache.scala 245:47]
  wire  _GEN_1890 = _GEN_1687 ? _GEN_919 : _GEN_919; // @[d_cache.scala 245:47]
  wire  _GEN_1891 = _GEN_1687 ? _GEN_920 : _GEN_920; // @[d_cache.scala 245:47]
  wire  _GEN_1892 = _GEN_1687 ? _GEN_921 : _GEN_921; // @[d_cache.scala 245:47]
  wire  _GEN_1893 = _GEN_1687 ? _GEN_922 : _GEN_922; // @[d_cache.scala 245:47]
  wire  _GEN_1894 = _GEN_1687 ? _GEN_923 : _GEN_923; // @[d_cache.scala 245:47]
  wire  _GEN_1895 = _GEN_1687 ? _GEN_924 : _GEN_924; // @[d_cache.scala 245:47]
  wire  _GEN_1896 = _GEN_1687 ? _GEN_925 : _GEN_925; // @[d_cache.scala 245:47]
  wire  _GEN_1897 = _GEN_1687 ? _GEN_926 : _GEN_926; // @[d_cache.scala 245:47]
  wire [3:0] _GEN_1898 = _GEN_1687 ? 4'h6 : 4'h1; // @[d_cache.scala 245:47 252:31 255:31]
  wire [7:0] _GEN_1899 = _GEN_1687 ? _GEN_927 : _GEN_927; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1900 = _GEN_1687 ? _GEN_928 : _GEN_928; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1901 = _GEN_1687 ? _GEN_929 : _GEN_929; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1902 = _GEN_1687 ? _GEN_930 : _GEN_930; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1903 = _GEN_1687 ? _GEN_931 : _GEN_931; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1904 = _GEN_1687 ? _GEN_932 : _GEN_932; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1905 = _GEN_1687 ? _GEN_933 : _GEN_933; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1906 = _GEN_1687 ? _GEN_934 : _GEN_934; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1907 = _GEN_1687 ? _GEN_935 : _GEN_935; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1908 = _GEN_1687 ? _GEN_936 : _GEN_936; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1909 = _GEN_1687 ? _GEN_937 : _GEN_937; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1910 = _GEN_1687 ? _GEN_938 : _GEN_938; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1911 = _GEN_1687 ? _GEN_939 : _GEN_939; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1912 = _GEN_1687 ? _GEN_940 : _GEN_940; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1913 = _GEN_1687 ? _GEN_941 : _GEN_941; // @[d_cache.scala 245:47]
  wire [7:0] _GEN_1914 = _GEN_1687 ? _GEN_942 : _GEN_942; // @[d_cache.scala 245:47]
  wire [511:0] _GEN_1915 = _GEN_734[7:6] == 2'h2 ? _GEN_1589 : _GEN_1832; // @[d_cache.scala 227:52]
  wire [41:0] _GEN_1916 = _GEN_734[7:6] == 2'h2 ? _GEN_1590 : _GEN_1833; // @[d_cache.scala 227:52]
  wire [511:0] _GEN_1917 = _GEN_734[7:6] == 2'h2 ? _GEN_1591 : ram_2_0; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1918 = _GEN_734[7:6] == 2'h2 ? _GEN_1592 : ram_2_1; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1919 = _GEN_734[7:6] == 2'h2 ? _GEN_1593 : ram_2_2; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1920 = _GEN_734[7:6] == 2'h2 ? _GEN_1594 : ram_2_3; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1921 = _GEN_734[7:6] == 2'h2 ? _GEN_1595 : ram_2_4; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1922 = _GEN_734[7:6] == 2'h2 ? _GEN_1596 : ram_2_5; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1923 = _GEN_734[7:6] == 2'h2 ? _GEN_1597 : ram_2_6; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1924 = _GEN_734[7:6] == 2'h2 ? _GEN_1598 : ram_2_7; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1925 = _GEN_734[7:6] == 2'h2 ? _GEN_1599 : ram_2_8; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1926 = _GEN_734[7:6] == 2'h2 ? _GEN_1600 : ram_2_9; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1927 = _GEN_734[7:6] == 2'h2 ? _GEN_1601 : ram_2_10; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1928 = _GEN_734[7:6] == 2'h2 ? _GEN_1602 : ram_2_11; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1929 = _GEN_734[7:6] == 2'h2 ? _GEN_1603 : ram_2_12; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1930 = _GEN_734[7:6] == 2'h2 ? _GEN_1604 : ram_2_13; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1931 = _GEN_734[7:6] == 2'h2 ? _GEN_1605 : ram_2_14; // @[d_cache.scala 21:24 227:52]
  wire [511:0] _GEN_1932 = _GEN_734[7:6] == 2'h2 ? _GEN_1606 : ram_2_15; // @[d_cache.scala 21:24 227:52]
  wire [31:0] _GEN_1933 = _GEN_734[7:6] == 2'h2 ? _GEN_1607 : tag_2_0; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1934 = _GEN_734[7:6] == 2'h2 ? _GEN_1608 : tag_2_1; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1935 = _GEN_734[7:6] == 2'h2 ? _GEN_1609 : tag_2_2; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1936 = _GEN_734[7:6] == 2'h2 ? _GEN_1610 : tag_2_3; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1937 = _GEN_734[7:6] == 2'h2 ? _GEN_1611 : tag_2_4; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1938 = _GEN_734[7:6] == 2'h2 ? _GEN_1612 : tag_2_5; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1939 = _GEN_734[7:6] == 2'h2 ? _GEN_1613 : tag_2_6; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1940 = _GEN_734[7:6] == 2'h2 ? _GEN_1614 : tag_2_7; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1941 = _GEN_734[7:6] == 2'h2 ? _GEN_1615 : tag_2_8; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1942 = _GEN_734[7:6] == 2'h2 ? _GEN_1616 : tag_2_9; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1943 = _GEN_734[7:6] == 2'h2 ? _GEN_1617 : tag_2_10; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1944 = _GEN_734[7:6] == 2'h2 ? _GEN_1618 : tag_2_11; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1945 = _GEN_734[7:6] == 2'h2 ? _GEN_1619 : tag_2_12; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1946 = _GEN_734[7:6] == 2'h2 ? _GEN_1620 : tag_2_13; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1947 = _GEN_734[7:6] == 2'h2 ? _GEN_1621 : tag_2_14; // @[d_cache.scala 227:52 26:24]
  wire [31:0] _GEN_1948 = _GEN_734[7:6] == 2'h2 ? _GEN_1622 : tag_2_15; // @[d_cache.scala 227:52 26:24]
  wire  _GEN_1949 = _GEN_734[7:6] == 2'h2 ? _GEN_1623 : dirty_2_0; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1950 = _GEN_734[7:6] == 2'h2 ? _GEN_1624 : dirty_2_1; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1951 = _GEN_734[7:6] == 2'h2 ? _GEN_1625 : dirty_2_2; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1952 = _GEN_734[7:6] == 2'h2 ? _GEN_1626 : dirty_2_3; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1953 = _GEN_734[7:6] == 2'h2 ? _GEN_1627 : dirty_2_4; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1954 = _GEN_734[7:6] == 2'h2 ? _GEN_1628 : dirty_2_5; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1955 = _GEN_734[7:6] == 2'h2 ? _GEN_1629 : dirty_2_6; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1956 = _GEN_734[7:6] == 2'h2 ? _GEN_1630 : dirty_2_7; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1957 = _GEN_734[7:6] == 2'h2 ? _GEN_1631 : dirty_2_8; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1958 = _GEN_734[7:6] == 2'h2 ? _GEN_1632 : dirty_2_9; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1959 = _GEN_734[7:6] == 2'h2 ? _GEN_1633 : dirty_2_10; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1960 = _GEN_734[7:6] == 2'h2 ? _GEN_1634 : dirty_2_11; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1961 = _GEN_734[7:6] == 2'h2 ? _GEN_1635 : dirty_2_12; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1962 = _GEN_734[7:6] == 2'h2 ? _GEN_1636 : dirty_2_13; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1963 = _GEN_734[7:6] == 2'h2 ? _GEN_1637 : dirty_2_14; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1964 = _GEN_734[7:6] == 2'h2 ? _GEN_1638 : dirty_2_15; // @[d_cache.scala 227:52 36:26]
  wire  _GEN_1965 = _GEN_734[7:6] == 2'h2 ? _GEN_1639 : valid_2_0; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1966 = _GEN_734[7:6] == 2'h2 ? _GEN_1640 : valid_2_1; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1967 = _GEN_734[7:6] == 2'h2 ? _GEN_1641 : valid_2_2; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1968 = _GEN_734[7:6] == 2'h2 ? _GEN_1642 : valid_2_3; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1969 = _GEN_734[7:6] == 2'h2 ? _GEN_1643 : valid_2_4; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1970 = _GEN_734[7:6] == 2'h2 ? _GEN_1644 : valid_2_5; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1971 = _GEN_734[7:6] == 2'h2 ? _GEN_1645 : valid_2_6; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1972 = _GEN_734[7:6] == 2'h2 ? _GEN_1646 : valid_2_7; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1973 = _GEN_734[7:6] == 2'h2 ? _GEN_1647 : valid_2_8; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1974 = _GEN_734[7:6] == 2'h2 ? _GEN_1648 : valid_2_9; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1975 = _GEN_734[7:6] == 2'h2 ? _GEN_1649 : valid_2_10; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1976 = _GEN_734[7:6] == 2'h2 ? _GEN_1650 : valid_2_11; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1977 = _GEN_734[7:6] == 2'h2 ? _GEN_1651 : valid_2_12; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1978 = _GEN_734[7:6] == 2'h2 ? _GEN_1652 : valid_2_13; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1979 = _GEN_734[7:6] == 2'h2 ? _GEN_1653 : valid_2_14; // @[d_cache.scala 227:52 31:26]
  wire  _GEN_1980 = _GEN_734[7:6] == 2'h2 ? _GEN_1654 : valid_2_15; // @[d_cache.scala 227:52 31:26]
  wire [3:0] _GEN_1981 = _GEN_734[7:6] == 2'h2 ? _GEN_1655 : _GEN_1898; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1982 = _GEN_734[7:6] == 2'h2 ? _GEN_1656 : _GEN_1899; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1983 = _GEN_734[7:6] == 2'h2 ? _GEN_1657 : _GEN_1900; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1984 = _GEN_734[7:6] == 2'h2 ? _GEN_1658 : _GEN_1901; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1985 = _GEN_734[7:6] == 2'h2 ? _GEN_1659 : _GEN_1902; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1986 = _GEN_734[7:6] == 2'h2 ? _GEN_1660 : _GEN_1903; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1987 = _GEN_734[7:6] == 2'h2 ? _GEN_1661 : _GEN_1904; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1988 = _GEN_734[7:6] == 2'h2 ? _GEN_1662 : _GEN_1905; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1989 = _GEN_734[7:6] == 2'h2 ? _GEN_1663 : _GEN_1906; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1990 = _GEN_734[7:6] == 2'h2 ? _GEN_1664 : _GEN_1907; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1991 = _GEN_734[7:6] == 2'h2 ? _GEN_1665 : _GEN_1908; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1992 = _GEN_734[7:6] == 2'h2 ? _GEN_1666 : _GEN_1909; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1993 = _GEN_734[7:6] == 2'h2 ? _GEN_1667 : _GEN_1910; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1994 = _GEN_734[7:6] == 2'h2 ? _GEN_1668 : _GEN_1911; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1995 = _GEN_734[7:6] == 2'h2 ? _GEN_1669 : _GEN_1912; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1996 = _GEN_734[7:6] == 2'h2 ? _GEN_1670 : _GEN_1913; // @[d_cache.scala 227:52]
  wire [7:0] _GEN_1997 = _GEN_734[7:6] == 2'h2 ? _GEN_1671 : _GEN_1914; // @[d_cache.scala 227:52]
  wire [511:0] _GEN_1998 = _GEN_734[7:6] == 2'h2 ? ram_3_0 : _GEN_1834; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_1999 = _GEN_734[7:6] == 2'h2 ? ram_3_1 : _GEN_1835; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2000 = _GEN_734[7:6] == 2'h2 ? ram_3_2 : _GEN_1836; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2001 = _GEN_734[7:6] == 2'h2 ? ram_3_3 : _GEN_1837; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2002 = _GEN_734[7:6] == 2'h2 ? ram_3_4 : _GEN_1838; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2003 = _GEN_734[7:6] == 2'h2 ? ram_3_5 : _GEN_1839; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2004 = _GEN_734[7:6] == 2'h2 ? ram_3_6 : _GEN_1840; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2005 = _GEN_734[7:6] == 2'h2 ? ram_3_7 : _GEN_1841; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2006 = _GEN_734[7:6] == 2'h2 ? ram_3_8 : _GEN_1842; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2007 = _GEN_734[7:6] == 2'h2 ? ram_3_9 : _GEN_1843; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2008 = _GEN_734[7:6] == 2'h2 ? ram_3_10 : _GEN_1844; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2009 = _GEN_734[7:6] == 2'h2 ? ram_3_11 : _GEN_1845; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2010 = _GEN_734[7:6] == 2'h2 ? ram_3_12 : _GEN_1846; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2011 = _GEN_734[7:6] == 2'h2 ? ram_3_13 : _GEN_1847; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2012 = _GEN_734[7:6] == 2'h2 ? ram_3_14 : _GEN_1848; // @[d_cache.scala 22:24 227:52]
  wire [511:0] _GEN_2013 = _GEN_734[7:6] == 2'h2 ? ram_3_15 : _GEN_1849; // @[d_cache.scala 22:24 227:52]
  wire [31:0] _GEN_2014 = _GEN_734[7:6] == 2'h2 ? tag_3_0 : _GEN_1850; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2015 = _GEN_734[7:6] == 2'h2 ? tag_3_1 : _GEN_1851; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2016 = _GEN_734[7:6] == 2'h2 ? tag_3_2 : _GEN_1852; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2017 = _GEN_734[7:6] == 2'h2 ? tag_3_3 : _GEN_1853; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2018 = _GEN_734[7:6] == 2'h2 ? tag_3_4 : _GEN_1854; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2019 = _GEN_734[7:6] == 2'h2 ? tag_3_5 : _GEN_1855; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2020 = _GEN_734[7:6] == 2'h2 ? tag_3_6 : _GEN_1856; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2021 = _GEN_734[7:6] == 2'h2 ? tag_3_7 : _GEN_1857; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2022 = _GEN_734[7:6] == 2'h2 ? tag_3_8 : _GEN_1858; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2023 = _GEN_734[7:6] == 2'h2 ? tag_3_9 : _GEN_1859; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2024 = _GEN_734[7:6] == 2'h2 ? tag_3_10 : _GEN_1860; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2025 = _GEN_734[7:6] == 2'h2 ? tag_3_11 : _GEN_1861; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2026 = _GEN_734[7:6] == 2'h2 ? tag_3_12 : _GEN_1862; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2027 = _GEN_734[7:6] == 2'h2 ? tag_3_13 : _GEN_1863; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2028 = _GEN_734[7:6] == 2'h2 ? tag_3_14 : _GEN_1864; // @[d_cache.scala 227:52 27:24]
  wire [31:0] _GEN_2029 = _GEN_734[7:6] == 2'h2 ? tag_3_15 : _GEN_1865; // @[d_cache.scala 227:52 27:24]
  wire  _GEN_2030 = _GEN_734[7:6] == 2'h2 ? dirty_3_0 : _GEN_1866; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2031 = _GEN_734[7:6] == 2'h2 ? dirty_3_1 : _GEN_1867; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2032 = _GEN_734[7:6] == 2'h2 ? dirty_3_2 : _GEN_1868; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2033 = _GEN_734[7:6] == 2'h2 ? dirty_3_3 : _GEN_1869; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2034 = _GEN_734[7:6] == 2'h2 ? dirty_3_4 : _GEN_1870; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2035 = _GEN_734[7:6] == 2'h2 ? dirty_3_5 : _GEN_1871; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2036 = _GEN_734[7:6] == 2'h2 ? dirty_3_6 : _GEN_1872; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2037 = _GEN_734[7:6] == 2'h2 ? dirty_3_7 : _GEN_1873; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2038 = _GEN_734[7:6] == 2'h2 ? dirty_3_8 : _GEN_1874; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2039 = _GEN_734[7:6] == 2'h2 ? dirty_3_9 : _GEN_1875; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2040 = _GEN_734[7:6] == 2'h2 ? dirty_3_10 : _GEN_1876; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2041 = _GEN_734[7:6] == 2'h2 ? dirty_3_11 : _GEN_1877; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2042 = _GEN_734[7:6] == 2'h2 ? dirty_3_12 : _GEN_1878; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2043 = _GEN_734[7:6] == 2'h2 ? dirty_3_13 : _GEN_1879; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2044 = _GEN_734[7:6] == 2'h2 ? dirty_3_14 : _GEN_1880; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2045 = _GEN_734[7:6] == 2'h2 ? dirty_3_15 : _GEN_1881; // @[d_cache.scala 227:52 37:26]
  wire  _GEN_2046 = _GEN_734[7:6] == 2'h2 ? valid_3_0 : _GEN_1882; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2047 = _GEN_734[7:6] == 2'h2 ? valid_3_1 : _GEN_1883; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2048 = _GEN_734[7:6] == 2'h2 ? valid_3_2 : _GEN_1884; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2049 = _GEN_734[7:6] == 2'h2 ? valid_3_3 : _GEN_1885; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2050 = _GEN_734[7:6] == 2'h2 ? valid_3_4 : _GEN_1886; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2051 = _GEN_734[7:6] == 2'h2 ? valid_3_5 : _GEN_1887; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2052 = _GEN_734[7:6] == 2'h2 ? valid_3_6 : _GEN_1888; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2053 = _GEN_734[7:6] == 2'h2 ? valid_3_7 : _GEN_1889; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2054 = _GEN_734[7:6] == 2'h2 ? valid_3_8 : _GEN_1890; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2055 = _GEN_734[7:6] == 2'h2 ? valid_3_9 : _GEN_1891; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2056 = _GEN_734[7:6] == 2'h2 ? valid_3_10 : _GEN_1892; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2057 = _GEN_734[7:6] == 2'h2 ? valid_3_11 : _GEN_1893; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2058 = _GEN_734[7:6] == 2'h2 ? valid_3_12 : _GEN_1894; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2059 = _GEN_734[7:6] == 2'h2 ? valid_3_13 : _GEN_1895; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2060 = _GEN_734[7:6] == 2'h2 ? valid_3_14 : _GEN_1896; // @[d_cache.scala 227:52 32:26]
  wire  _GEN_2061 = _GEN_734[7:6] == 2'h2 ? valid_3_15 : _GEN_1897; // @[d_cache.scala 227:52 32:26]
  wire [511:0] _GEN_2062 = _GEN_734[7:6] == 2'h1 ? _GEN_1346 : _GEN_1915; // @[d_cache.scala 210:52]
  wire [41:0] _GEN_2063 = _GEN_734[7:6] == 2'h1 ? _GEN_1347 : _GEN_1916; // @[d_cache.scala 210:52]
  wire [511:0] _GEN_2064 = _GEN_734[7:6] == 2'h1 ? _GEN_1348 : ram_1_0; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2065 = _GEN_734[7:6] == 2'h1 ? _GEN_1349 : ram_1_1; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2066 = _GEN_734[7:6] == 2'h1 ? _GEN_1350 : ram_1_2; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2067 = _GEN_734[7:6] == 2'h1 ? _GEN_1351 : ram_1_3; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2068 = _GEN_734[7:6] == 2'h1 ? _GEN_1352 : ram_1_4; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2069 = _GEN_734[7:6] == 2'h1 ? _GEN_1353 : ram_1_5; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2070 = _GEN_734[7:6] == 2'h1 ? _GEN_1354 : ram_1_6; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2071 = _GEN_734[7:6] == 2'h1 ? _GEN_1355 : ram_1_7; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2072 = _GEN_734[7:6] == 2'h1 ? _GEN_1356 : ram_1_8; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2073 = _GEN_734[7:6] == 2'h1 ? _GEN_1357 : ram_1_9; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2074 = _GEN_734[7:6] == 2'h1 ? _GEN_1358 : ram_1_10; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2075 = _GEN_734[7:6] == 2'h1 ? _GEN_1359 : ram_1_11; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2076 = _GEN_734[7:6] == 2'h1 ? _GEN_1360 : ram_1_12; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2077 = _GEN_734[7:6] == 2'h1 ? _GEN_1361 : ram_1_13; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2078 = _GEN_734[7:6] == 2'h1 ? _GEN_1362 : ram_1_14; // @[d_cache.scala 20:24 210:52]
  wire [511:0] _GEN_2079 = _GEN_734[7:6] == 2'h1 ? _GEN_1363 : ram_1_15; // @[d_cache.scala 20:24 210:52]
  wire [31:0] _GEN_2080 = _GEN_734[7:6] == 2'h1 ? _GEN_1364 : tag_1_0; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2081 = _GEN_734[7:6] == 2'h1 ? _GEN_1365 : tag_1_1; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2082 = _GEN_734[7:6] == 2'h1 ? _GEN_1366 : tag_1_2; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2083 = _GEN_734[7:6] == 2'h1 ? _GEN_1367 : tag_1_3; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2084 = _GEN_734[7:6] == 2'h1 ? _GEN_1368 : tag_1_4; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2085 = _GEN_734[7:6] == 2'h1 ? _GEN_1369 : tag_1_5; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2086 = _GEN_734[7:6] == 2'h1 ? _GEN_1370 : tag_1_6; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2087 = _GEN_734[7:6] == 2'h1 ? _GEN_1371 : tag_1_7; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2088 = _GEN_734[7:6] == 2'h1 ? _GEN_1372 : tag_1_8; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2089 = _GEN_734[7:6] == 2'h1 ? _GEN_1373 : tag_1_9; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2090 = _GEN_734[7:6] == 2'h1 ? _GEN_1374 : tag_1_10; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2091 = _GEN_734[7:6] == 2'h1 ? _GEN_1375 : tag_1_11; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2092 = _GEN_734[7:6] == 2'h1 ? _GEN_1376 : tag_1_12; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2093 = _GEN_734[7:6] == 2'h1 ? _GEN_1377 : tag_1_13; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2094 = _GEN_734[7:6] == 2'h1 ? _GEN_1378 : tag_1_14; // @[d_cache.scala 210:52 25:24]
  wire [31:0] _GEN_2095 = _GEN_734[7:6] == 2'h1 ? _GEN_1379 : tag_1_15; // @[d_cache.scala 210:52 25:24]
  wire  _GEN_2096 = _GEN_734[7:6] == 2'h1 ? _GEN_1380 : dirty_1_0; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2097 = _GEN_734[7:6] == 2'h1 ? _GEN_1381 : dirty_1_1; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2098 = _GEN_734[7:6] == 2'h1 ? _GEN_1382 : dirty_1_2; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2099 = _GEN_734[7:6] == 2'h1 ? _GEN_1383 : dirty_1_3; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2100 = _GEN_734[7:6] == 2'h1 ? _GEN_1384 : dirty_1_4; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2101 = _GEN_734[7:6] == 2'h1 ? _GEN_1385 : dirty_1_5; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2102 = _GEN_734[7:6] == 2'h1 ? _GEN_1386 : dirty_1_6; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2103 = _GEN_734[7:6] == 2'h1 ? _GEN_1387 : dirty_1_7; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2104 = _GEN_734[7:6] == 2'h1 ? _GEN_1388 : dirty_1_8; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2105 = _GEN_734[7:6] == 2'h1 ? _GEN_1389 : dirty_1_9; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2106 = _GEN_734[7:6] == 2'h1 ? _GEN_1390 : dirty_1_10; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2107 = _GEN_734[7:6] == 2'h1 ? _GEN_1391 : dirty_1_11; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2108 = _GEN_734[7:6] == 2'h1 ? _GEN_1392 : dirty_1_12; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2109 = _GEN_734[7:6] == 2'h1 ? _GEN_1393 : dirty_1_13; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2110 = _GEN_734[7:6] == 2'h1 ? _GEN_1394 : dirty_1_14; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2111 = _GEN_734[7:6] == 2'h1 ? _GEN_1395 : dirty_1_15; // @[d_cache.scala 210:52 35:26]
  wire  _GEN_2112 = _GEN_734[7:6] == 2'h1 ? _GEN_1396 : valid_1_0; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2113 = _GEN_734[7:6] == 2'h1 ? _GEN_1397 : valid_1_1; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2114 = _GEN_734[7:6] == 2'h1 ? _GEN_1398 : valid_1_2; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2115 = _GEN_734[7:6] == 2'h1 ? _GEN_1399 : valid_1_3; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2116 = _GEN_734[7:6] == 2'h1 ? _GEN_1400 : valid_1_4; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2117 = _GEN_734[7:6] == 2'h1 ? _GEN_1401 : valid_1_5; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2118 = _GEN_734[7:6] == 2'h1 ? _GEN_1402 : valid_1_6; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2119 = _GEN_734[7:6] == 2'h1 ? _GEN_1403 : valid_1_7; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2120 = _GEN_734[7:6] == 2'h1 ? _GEN_1404 : valid_1_8; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2121 = _GEN_734[7:6] == 2'h1 ? _GEN_1405 : valid_1_9; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2122 = _GEN_734[7:6] == 2'h1 ? _GEN_1406 : valid_1_10; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2123 = _GEN_734[7:6] == 2'h1 ? _GEN_1407 : valid_1_11; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2124 = _GEN_734[7:6] == 2'h1 ? _GEN_1408 : valid_1_12; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2125 = _GEN_734[7:6] == 2'h1 ? _GEN_1409 : valid_1_13; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2126 = _GEN_734[7:6] == 2'h1 ? _GEN_1410 : valid_1_14; // @[d_cache.scala 210:52 30:26]
  wire  _GEN_2127 = _GEN_734[7:6] == 2'h1 ? _GEN_1411 : valid_1_15; // @[d_cache.scala 210:52 30:26]
  wire [3:0] _GEN_2128 = _GEN_734[7:6] == 2'h1 ? _GEN_1412 : _GEN_1981; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2129 = _GEN_734[7:6] == 2'h1 ? _GEN_1413 : _GEN_1982; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2130 = _GEN_734[7:6] == 2'h1 ? _GEN_1414 : _GEN_1983; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2131 = _GEN_734[7:6] == 2'h1 ? _GEN_1415 : _GEN_1984; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2132 = _GEN_734[7:6] == 2'h1 ? _GEN_1416 : _GEN_1985; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2133 = _GEN_734[7:6] == 2'h1 ? _GEN_1417 : _GEN_1986; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2134 = _GEN_734[7:6] == 2'h1 ? _GEN_1418 : _GEN_1987; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2135 = _GEN_734[7:6] == 2'h1 ? _GEN_1419 : _GEN_1988; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2136 = _GEN_734[7:6] == 2'h1 ? _GEN_1420 : _GEN_1989; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2137 = _GEN_734[7:6] == 2'h1 ? _GEN_1421 : _GEN_1990; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2138 = _GEN_734[7:6] == 2'h1 ? _GEN_1422 : _GEN_1991; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2139 = _GEN_734[7:6] == 2'h1 ? _GEN_1423 : _GEN_1992; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2140 = _GEN_734[7:6] == 2'h1 ? _GEN_1424 : _GEN_1993; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2141 = _GEN_734[7:6] == 2'h1 ? _GEN_1425 : _GEN_1994; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2142 = _GEN_734[7:6] == 2'h1 ? _GEN_1426 : _GEN_1995; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2143 = _GEN_734[7:6] == 2'h1 ? _GEN_1427 : _GEN_1996; // @[d_cache.scala 210:52]
  wire [7:0] _GEN_2144 = _GEN_734[7:6] == 2'h1 ? _GEN_1428 : _GEN_1997; // @[d_cache.scala 210:52]
  wire [511:0] _GEN_2145 = _GEN_734[7:6] == 2'h1 ? ram_2_0 : _GEN_1917; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2146 = _GEN_734[7:6] == 2'h1 ? ram_2_1 : _GEN_1918; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2147 = _GEN_734[7:6] == 2'h1 ? ram_2_2 : _GEN_1919; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2148 = _GEN_734[7:6] == 2'h1 ? ram_2_3 : _GEN_1920; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2149 = _GEN_734[7:6] == 2'h1 ? ram_2_4 : _GEN_1921; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2150 = _GEN_734[7:6] == 2'h1 ? ram_2_5 : _GEN_1922; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2151 = _GEN_734[7:6] == 2'h1 ? ram_2_6 : _GEN_1923; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2152 = _GEN_734[7:6] == 2'h1 ? ram_2_7 : _GEN_1924; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2153 = _GEN_734[7:6] == 2'h1 ? ram_2_8 : _GEN_1925; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2154 = _GEN_734[7:6] == 2'h1 ? ram_2_9 : _GEN_1926; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2155 = _GEN_734[7:6] == 2'h1 ? ram_2_10 : _GEN_1927; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2156 = _GEN_734[7:6] == 2'h1 ? ram_2_11 : _GEN_1928; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2157 = _GEN_734[7:6] == 2'h1 ? ram_2_12 : _GEN_1929; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2158 = _GEN_734[7:6] == 2'h1 ? ram_2_13 : _GEN_1930; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2159 = _GEN_734[7:6] == 2'h1 ? ram_2_14 : _GEN_1931; // @[d_cache.scala 21:24 210:52]
  wire [511:0] _GEN_2160 = _GEN_734[7:6] == 2'h1 ? ram_2_15 : _GEN_1932; // @[d_cache.scala 21:24 210:52]
  wire [31:0] _GEN_2161 = _GEN_734[7:6] == 2'h1 ? tag_2_0 : _GEN_1933; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2162 = _GEN_734[7:6] == 2'h1 ? tag_2_1 : _GEN_1934; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2163 = _GEN_734[7:6] == 2'h1 ? tag_2_2 : _GEN_1935; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2164 = _GEN_734[7:6] == 2'h1 ? tag_2_3 : _GEN_1936; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2165 = _GEN_734[7:6] == 2'h1 ? tag_2_4 : _GEN_1937; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2166 = _GEN_734[7:6] == 2'h1 ? tag_2_5 : _GEN_1938; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2167 = _GEN_734[7:6] == 2'h1 ? tag_2_6 : _GEN_1939; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2168 = _GEN_734[7:6] == 2'h1 ? tag_2_7 : _GEN_1940; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2169 = _GEN_734[7:6] == 2'h1 ? tag_2_8 : _GEN_1941; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2170 = _GEN_734[7:6] == 2'h1 ? tag_2_9 : _GEN_1942; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2171 = _GEN_734[7:6] == 2'h1 ? tag_2_10 : _GEN_1943; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2172 = _GEN_734[7:6] == 2'h1 ? tag_2_11 : _GEN_1944; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2173 = _GEN_734[7:6] == 2'h1 ? tag_2_12 : _GEN_1945; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2174 = _GEN_734[7:6] == 2'h1 ? tag_2_13 : _GEN_1946; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2175 = _GEN_734[7:6] == 2'h1 ? tag_2_14 : _GEN_1947; // @[d_cache.scala 210:52 26:24]
  wire [31:0] _GEN_2176 = _GEN_734[7:6] == 2'h1 ? tag_2_15 : _GEN_1948; // @[d_cache.scala 210:52 26:24]
  wire  _GEN_2177 = _GEN_734[7:6] == 2'h1 ? dirty_2_0 : _GEN_1949; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2178 = _GEN_734[7:6] == 2'h1 ? dirty_2_1 : _GEN_1950; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2179 = _GEN_734[7:6] == 2'h1 ? dirty_2_2 : _GEN_1951; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2180 = _GEN_734[7:6] == 2'h1 ? dirty_2_3 : _GEN_1952; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2181 = _GEN_734[7:6] == 2'h1 ? dirty_2_4 : _GEN_1953; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2182 = _GEN_734[7:6] == 2'h1 ? dirty_2_5 : _GEN_1954; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2183 = _GEN_734[7:6] == 2'h1 ? dirty_2_6 : _GEN_1955; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2184 = _GEN_734[7:6] == 2'h1 ? dirty_2_7 : _GEN_1956; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2185 = _GEN_734[7:6] == 2'h1 ? dirty_2_8 : _GEN_1957; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2186 = _GEN_734[7:6] == 2'h1 ? dirty_2_9 : _GEN_1958; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2187 = _GEN_734[7:6] == 2'h1 ? dirty_2_10 : _GEN_1959; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2188 = _GEN_734[7:6] == 2'h1 ? dirty_2_11 : _GEN_1960; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2189 = _GEN_734[7:6] == 2'h1 ? dirty_2_12 : _GEN_1961; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2190 = _GEN_734[7:6] == 2'h1 ? dirty_2_13 : _GEN_1962; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2191 = _GEN_734[7:6] == 2'h1 ? dirty_2_14 : _GEN_1963; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2192 = _GEN_734[7:6] == 2'h1 ? dirty_2_15 : _GEN_1964; // @[d_cache.scala 210:52 36:26]
  wire  _GEN_2193 = _GEN_734[7:6] == 2'h1 ? valid_2_0 : _GEN_1965; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2194 = _GEN_734[7:6] == 2'h1 ? valid_2_1 : _GEN_1966; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2195 = _GEN_734[7:6] == 2'h1 ? valid_2_2 : _GEN_1967; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2196 = _GEN_734[7:6] == 2'h1 ? valid_2_3 : _GEN_1968; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2197 = _GEN_734[7:6] == 2'h1 ? valid_2_4 : _GEN_1969; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2198 = _GEN_734[7:6] == 2'h1 ? valid_2_5 : _GEN_1970; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2199 = _GEN_734[7:6] == 2'h1 ? valid_2_6 : _GEN_1971; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2200 = _GEN_734[7:6] == 2'h1 ? valid_2_7 : _GEN_1972; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2201 = _GEN_734[7:6] == 2'h1 ? valid_2_8 : _GEN_1973; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2202 = _GEN_734[7:6] == 2'h1 ? valid_2_9 : _GEN_1974; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2203 = _GEN_734[7:6] == 2'h1 ? valid_2_10 : _GEN_1975; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2204 = _GEN_734[7:6] == 2'h1 ? valid_2_11 : _GEN_1976; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2205 = _GEN_734[7:6] == 2'h1 ? valid_2_12 : _GEN_1977; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2206 = _GEN_734[7:6] == 2'h1 ? valid_2_13 : _GEN_1978; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2207 = _GEN_734[7:6] == 2'h1 ? valid_2_14 : _GEN_1979; // @[d_cache.scala 210:52 31:26]
  wire  _GEN_2208 = _GEN_734[7:6] == 2'h1 ? valid_2_15 : _GEN_1980; // @[d_cache.scala 210:52 31:26]
  wire [511:0] _GEN_2209 = _GEN_734[7:6] == 2'h1 ? ram_3_0 : _GEN_1998; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2210 = _GEN_734[7:6] == 2'h1 ? ram_3_1 : _GEN_1999; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2211 = _GEN_734[7:6] == 2'h1 ? ram_3_2 : _GEN_2000; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2212 = _GEN_734[7:6] == 2'h1 ? ram_3_3 : _GEN_2001; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2213 = _GEN_734[7:6] == 2'h1 ? ram_3_4 : _GEN_2002; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2214 = _GEN_734[7:6] == 2'h1 ? ram_3_5 : _GEN_2003; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2215 = _GEN_734[7:6] == 2'h1 ? ram_3_6 : _GEN_2004; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2216 = _GEN_734[7:6] == 2'h1 ? ram_3_7 : _GEN_2005; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2217 = _GEN_734[7:6] == 2'h1 ? ram_3_8 : _GEN_2006; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2218 = _GEN_734[7:6] == 2'h1 ? ram_3_9 : _GEN_2007; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2219 = _GEN_734[7:6] == 2'h1 ? ram_3_10 : _GEN_2008; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2220 = _GEN_734[7:6] == 2'h1 ? ram_3_11 : _GEN_2009; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2221 = _GEN_734[7:6] == 2'h1 ? ram_3_12 : _GEN_2010; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2222 = _GEN_734[7:6] == 2'h1 ? ram_3_13 : _GEN_2011; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2223 = _GEN_734[7:6] == 2'h1 ? ram_3_14 : _GEN_2012; // @[d_cache.scala 210:52 22:24]
  wire [511:0] _GEN_2224 = _GEN_734[7:6] == 2'h1 ? ram_3_15 : _GEN_2013; // @[d_cache.scala 210:52 22:24]
  wire [31:0] _GEN_2225 = _GEN_734[7:6] == 2'h1 ? tag_3_0 : _GEN_2014; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2226 = _GEN_734[7:6] == 2'h1 ? tag_3_1 : _GEN_2015; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2227 = _GEN_734[7:6] == 2'h1 ? tag_3_2 : _GEN_2016; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2228 = _GEN_734[7:6] == 2'h1 ? tag_3_3 : _GEN_2017; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2229 = _GEN_734[7:6] == 2'h1 ? tag_3_4 : _GEN_2018; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2230 = _GEN_734[7:6] == 2'h1 ? tag_3_5 : _GEN_2019; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2231 = _GEN_734[7:6] == 2'h1 ? tag_3_6 : _GEN_2020; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2232 = _GEN_734[7:6] == 2'h1 ? tag_3_7 : _GEN_2021; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2233 = _GEN_734[7:6] == 2'h1 ? tag_3_8 : _GEN_2022; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2234 = _GEN_734[7:6] == 2'h1 ? tag_3_9 : _GEN_2023; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2235 = _GEN_734[7:6] == 2'h1 ? tag_3_10 : _GEN_2024; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2236 = _GEN_734[7:6] == 2'h1 ? tag_3_11 : _GEN_2025; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2237 = _GEN_734[7:6] == 2'h1 ? tag_3_12 : _GEN_2026; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2238 = _GEN_734[7:6] == 2'h1 ? tag_3_13 : _GEN_2027; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2239 = _GEN_734[7:6] == 2'h1 ? tag_3_14 : _GEN_2028; // @[d_cache.scala 210:52 27:24]
  wire [31:0] _GEN_2240 = _GEN_734[7:6] == 2'h1 ? tag_3_15 : _GEN_2029; // @[d_cache.scala 210:52 27:24]
  wire  _GEN_2241 = _GEN_734[7:6] == 2'h1 ? dirty_3_0 : _GEN_2030; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2242 = _GEN_734[7:6] == 2'h1 ? dirty_3_1 : _GEN_2031; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2243 = _GEN_734[7:6] == 2'h1 ? dirty_3_2 : _GEN_2032; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2244 = _GEN_734[7:6] == 2'h1 ? dirty_3_3 : _GEN_2033; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2245 = _GEN_734[7:6] == 2'h1 ? dirty_3_4 : _GEN_2034; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2246 = _GEN_734[7:6] == 2'h1 ? dirty_3_5 : _GEN_2035; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2247 = _GEN_734[7:6] == 2'h1 ? dirty_3_6 : _GEN_2036; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2248 = _GEN_734[7:6] == 2'h1 ? dirty_3_7 : _GEN_2037; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2249 = _GEN_734[7:6] == 2'h1 ? dirty_3_8 : _GEN_2038; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2250 = _GEN_734[7:6] == 2'h1 ? dirty_3_9 : _GEN_2039; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2251 = _GEN_734[7:6] == 2'h1 ? dirty_3_10 : _GEN_2040; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2252 = _GEN_734[7:6] == 2'h1 ? dirty_3_11 : _GEN_2041; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2253 = _GEN_734[7:6] == 2'h1 ? dirty_3_12 : _GEN_2042; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2254 = _GEN_734[7:6] == 2'h1 ? dirty_3_13 : _GEN_2043; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2255 = _GEN_734[7:6] == 2'h1 ? dirty_3_14 : _GEN_2044; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2256 = _GEN_734[7:6] == 2'h1 ? dirty_3_15 : _GEN_2045; // @[d_cache.scala 210:52 37:26]
  wire  _GEN_2257 = _GEN_734[7:6] == 2'h1 ? valid_3_0 : _GEN_2046; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2258 = _GEN_734[7:6] == 2'h1 ? valid_3_1 : _GEN_2047; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2259 = _GEN_734[7:6] == 2'h1 ? valid_3_2 : _GEN_2048; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2260 = _GEN_734[7:6] == 2'h1 ? valid_3_3 : _GEN_2049; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2261 = _GEN_734[7:6] == 2'h1 ? valid_3_4 : _GEN_2050; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2262 = _GEN_734[7:6] == 2'h1 ? valid_3_5 : _GEN_2051; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2263 = _GEN_734[7:6] == 2'h1 ? valid_3_6 : _GEN_2052; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2264 = _GEN_734[7:6] == 2'h1 ? valid_3_7 : _GEN_2053; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2265 = _GEN_734[7:6] == 2'h1 ? valid_3_8 : _GEN_2054; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2266 = _GEN_734[7:6] == 2'h1 ? valid_3_9 : _GEN_2055; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2267 = _GEN_734[7:6] == 2'h1 ? valid_3_10 : _GEN_2056; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2268 = _GEN_734[7:6] == 2'h1 ? valid_3_11 : _GEN_2057; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2269 = _GEN_734[7:6] == 2'h1 ? valid_3_12 : _GEN_2058; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2270 = _GEN_734[7:6] == 2'h1 ? valid_3_13 : _GEN_2059; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2271 = _GEN_734[7:6] == 2'h1 ? valid_3_14 : _GEN_2060; // @[d_cache.scala 210:52 32:26]
  wire  _GEN_2272 = _GEN_734[7:6] == 2'h1 ? valid_3_15 : _GEN_2061; // @[d_cache.scala 210:52 32:26]
  wire [511:0] _GEN_2273 = _GEN_734[7:6] == 2'h0 ? _GEN_1103 : _GEN_2062; // @[d_cache.scala 193:46]
  wire [41:0] _GEN_2274 = _GEN_734[7:6] == 2'h0 ? _GEN_1104 : _GEN_2063; // @[d_cache.scala 193:46]
  wire [511:0] _GEN_2275 = _GEN_734[7:6] == 2'h0 ? _GEN_1105 : ram_0_0; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2276 = _GEN_734[7:6] == 2'h0 ? _GEN_1106 : ram_0_1; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2277 = _GEN_734[7:6] == 2'h0 ? _GEN_1107 : ram_0_2; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2278 = _GEN_734[7:6] == 2'h0 ? _GEN_1108 : ram_0_3; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2279 = _GEN_734[7:6] == 2'h0 ? _GEN_1109 : ram_0_4; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2280 = _GEN_734[7:6] == 2'h0 ? _GEN_1110 : ram_0_5; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2281 = _GEN_734[7:6] == 2'h0 ? _GEN_1111 : ram_0_6; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2282 = _GEN_734[7:6] == 2'h0 ? _GEN_1112 : ram_0_7; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2283 = _GEN_734[7:6] == 2'h0 ? _GEN_1113 : ram_0_8; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2284 = _GEN_734[7:6] == 2'h0 ? _GEN_1114 : ram_0_9; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2285 = _GEN_734[7:6] == 2'h0 ? _GEN_1115 : ram_0_10; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2286 = _GEN_734[7:6] == 2'h0 ? _GEN_1116 : ram_0_11; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2287 = _GEN_734[7:6] == 2'h0 ? _GEN_1117 : ram_0_12; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2288 = _GEN_734[7:6] == 2'h0 ? _GEN_1118 : ram_0_13; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2289 = _GEN_734[7:6] == 2'h0 ? _GEN_1119 : ram_0_14; // @[d_cache.scala 19:24 193:46]
  wire [511:0] _GEN_2290 = _GEN_734[7:6] == 2'h0 ? _GEN_1120 : ram_0_15; // @[d_cache.scala 19:24 193:46]
  wire [31:0] _GEN_2291 = _GEN_734[7:6] == 2'h0 ? _GEN_1121 : tag_0_0; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2292 = _GEN_734[7:6] == 2'h0 ? _GEN_1122 : tag_0_1; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2293 = _GEN_734[7:6] == 2'h0 ? _GEN_1123 : tag_0_2; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2294 = _GEN_734[7:6] == 2'h0 ? _GEN_1124 : tag_0_3; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2295 = _GEN_734[7:6] == 2'h0 ? _GEN_1125 : tag_0_4; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2296 = _GEN_734[7:6] == 2'h0 ? _GEN_1126 : tag_0_5; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2297 = _GEN_734[7:6] == 2'h0 ? _GEN_1127 : tag_0_6; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2298 = _GEN_734[7:6] == 2'h0 ? _GEN_1128 : tag_0_7; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2299 = _GEN_734[7:6] == 2'h0 ? _GEN_1129 : tag_0_8; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2300 = _GEN_734[7:6] == 2'h0 ? _GEN_1130 : tag_0_9; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2301 = _GEN_734[7:6] == 2'h0 ? _GEN_1131 : tag_0_10; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2302 = _GEN_734[7:6] == 2'h0 ? _GEN_1132 : tag_0_11; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2303 = _GEN_734[7:6] == 2'h0 ? _GEN_1133 : tag_0_12; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2304 = _GEN_734[7:6] == 2'h0 ? _GEN_1134 : tag_0_13; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2305 = _GEN_734[7:6] == 2'h0 ? _GEN_1135 : tag_0_14; // @[d_cache.scala 193:46 24:24]
  wire [31:0] _GEN_2306 = _GEN_734[7:6] == 2'h0 ? _GEN_1136 : tag_0_15; // @[d_cache.scala 193:46 24:24]
  wire  _GEN_2307 = _GEN_734[7:6] == 2'h0 ? _GEN_1137 : dirty_0_0; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2308 = _GEN_734[7:6] == 2'h0 ? _GEN_1138 : dirty_0_1; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2309 = _GEN_734[7:6] == 2'h0 ? _GEN_1139 : dirty_0_2; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2310 = _GEN_734[7:6] == 2'h0 ? _GEN_1140 : dirty_0_3; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2311 = _GEN_734[7:6] == 2'h0 ? _GEN_1141 : dirty_0_4; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2312 = _GEN_734[7:6] == 2'h0 ? _GEN_1142 : dirty_0_5; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2313 = _GEN_734[7:6] == 2'h0 ? _GEN_1143 : dirty_0_6; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2314 = _GEN_734[7:6] == 2'h0 ? _GEN_1144 : dirty_0_7; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2315 = _GEN_734[7:6] == 2'h0 ? _GEN_1145 : dirty_0_8; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2316 = _GEN_734[7:6] == 2'h0 ? _GEN_1146 : dirty_0_9; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2317 = _GEN_734[7:6] == 2'h0 ? _GEN_1147 : dirty_0_10; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2318 = _GEN_734[7:6] == 2'h0 ? _GEN_1148 : dirty_0_11; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2319 = _GEN_734[7:6] == 2'h0 ? _GEN_1149 : dirty_0_12; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2320 = _GEN_734[7:6] == 2'h0 ? _GEN_1150 : dirty_0_13; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2321 = _GEN_734[7:6] == 2'h0 ? _GEN_1151 : dirty_0_14; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2322 = _GEN_734[7:6] == 2'h0 ? _GEN_1152 : dirty_0_15; // @[d_cache.scala 193:46 34:26]
  wire  _GEN_2323 = _GEN_734[7:6] == 2'h0 ? _GEN_1153 : valid_0_0; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2324 = _GEN_734[7:6] == 2'h0 ? _GEN_1154 : valid_0_1; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2325 = _GEN_734[7:6] == 2'h0 ? _GEN_1155 : valid_0_2; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2326 = _GEN_734[7:6] == 2'h0 ? _GEN_1156 : valid_0_3; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2327 = _GEN_734[7:6] == 2'h0 ? _GEN_1157 : valid_0_4; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2328 = _GEN_734[7:6] == 2'h0 ? _GEN_1158 : valid_0_5; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2329 = _GEN_734[7:6] == 2'h0 ? _GEN_1159 : valid_0_6; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2330 = _GEN_734[7:6] == 2'h0 ? _GEN_1160 : valid_0_7; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2331 = _GEN_734[7:6] == 2'h0 ? _GEN_1161 : valid_0_8; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2332 = _GEN_734[7:6] == 2'h0 ? _GEN_1162 : valid_0_9; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2333 = _GEN_734[7:6] == 2'h0 ? _GEN_1163 : valid_0_10; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2334 = _GEN_734[7:6] == 2'h0 ? _GEN_1164 : valid_0_11; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2335 = _GEN_734[7:6] == 2'h0 ? _GEN_1165 : valid_0_12; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2336 = _GEN_734[7:6] == 2'h0 ? _GEN_1166 : valid_0_13; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2337 = _GEN_734[7:6] == 2'h0 ? _GEN_1167 : valid_0_14; // @[d_cache.scala 193:46 29:26]
  wire  _GEN_2338 = _GEN_734[7:6] == 2'h0 ? _GEN_1168 : valid_0_15; // @[d_cache.scala 193:46 29:26]
  wire [3:0] _GEN_2339 = _GEN_734[7:6] == 2'h0 ? _GEN_1169 : _GEN_2128; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2340 = _GEN_734[7:6] == 2'h0 ? _GEN_1170 : _GEN_2129; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2341 = _GEN_734[7:6] == 2'h0 ? _GEN_1171 : _GEN_2130; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2342 = _GEN_734[7:6] == 2'h0 ? _GEN_1172 : _GEN_2131; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2343 = _GEN_734[7:6] == 2'h0 ? _GEN_1173 : _GEN_2132; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2344 = _GEN_734[7:6] == 2'h0 ? _GEN_1174 : _GEN_2133; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2345 = _GEN_734[7:6] == 2'h0 ? _GEN_1175 : _GEN_2134; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2346 = _GEN_734[7:6] == 2'h0 ? _GEN_1176 : _GEN_2135; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2347 = _GEN_734[7:6] == 2'h0 ? _GEN_1177 : _GEN_2136; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2348 = _GEN_734[7:6] == 2'h0 ? _GEN_1178 : _GEN_2137; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2349 = _GEN_734[7:6] == 2'h0 ? _GEN_1179 : _GEN_2138; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2350 = _GEN_734[7:6] == 2'h0 ? _GEN_1180 : _GEN_2139; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2351 = _GEN_734[7:6] == 2'h0 ? _GEN_1181 : _GEN_2140; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2352 = _GEN_734[7:6] == 2'h0 ? _GEN_1182 : _GEN_2141; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2353 = _GEN_734[7:6] == 2'h0 ? _GEN_1183 : _GEN_2142; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2354 = _GEN_734[7:6] == 2'h0 ? _GEN_1184 : _GEN_2143; // @[d_cache.scala 193:46]
  wire [7:0] _GEN_2355 = _GEN_734[7:6] == 2'h0 ? _GEN_1185 : _GEN_2144; // @[d_cache.scala 193:46]
  wire [511:0] _GEN_2356 = _GEN_734[7:6] == 2'h0 ? ram_1_0 : _GEN_2064; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2357 = _GEN_734[7:6] == 2'h0 ? ram_1_1 : _GEN_2065; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2358 = _GEN_734[7:6] == 2'h0 ? ram_1_2 : _GEN_2066; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2359 = _GEN_734[7:6] == 2'h0 ? ram_1_3 : _GEN_2067; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2360 = _GEN_734[7:6] == 2'h0 ? ram_1_4 : _GEN_2068; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2361 = _GEN_734[7:6] == 2'h0 ? ram_1_5 : _GEN_2069; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2362 = _GEN_734[7:6] == 2'h0 ? ram_1_6 : _GEN_2070; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2363 = _GEN_734[7:6] == 2'h0 ? ram_1_7 : _GEN_2071; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2364 = _GEN_734[7:6] == 2'h0 ? ram_1_8 : _GEN_2072; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2365 = _GEN_734[7:6] == 2'h0 ? ram_1_9 : _GEN_2073; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2366 = _GEN_734[7:6] == 2'h0 ? ram_1_10 : _GEN_2074; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2367 = _GEN_734[7:6] == 2'h0 ? ram_1_11 : _GEN_2075; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2368 = _GEN_734[7:6] == 2'h0 ? ram_1_12 : _GEN_2076; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2369 = _GEN_734[7:6] == 2'h0 ? ram_1_13 : _GEN_2077; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2370 = _GEN_734[7:6] == 2'h0 ? ram_1_14 : _GEN_2078; // @[d_cache.scala 193:46 20:24]
  wire [511:0] _GEN_2371 = _GEN_734[7:6] == 2'h0 ? ram_1_15 : _GEN_2079; // @[d_cache.scala 193:46 20:24]
  wire [31:0] _GEN_2372 = _GEN_734[7:6] == 2'h0 ? tag_1_0 : _GEN_2080; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2373 = _GEN_734[7:6] == 2'h0 ? tag_1_1 : _GEN_2081; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2374 = _GEN_734[7:6] == 2'h0 ? tag_1_2 : _GEN_2082; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2375 = _GEN_734[7:6] == 2'h0 ? tag_1_3 : _GEN_2083; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2376 = _GEN_734[7:6] == 2'h0 ? tag_1_4 : _GEN_2084; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2377 = _GEN_734[7:6] == 2'h0 ? tag_1_5 : _GEN_2085; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2378 = _GEN_734[7:6] == 2'h0 ? tag_1_6 : _GEN_2086; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2379 = _GEN_734[7:6] == 2'h0 ? tag_1_7 : _GEN_2087; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2380 = _GEN_734[7:6] == 2'h0 ? tag_1_8 : _GEN_2088; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2381 = _GEN_734[7:6] == 2'h0 ? tag_1_9 : _GEN_2089; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2382 = _GEN_734[7:6] == 2'h0 ? tag_1_10 : _GEN_2090; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2383 = _GEN_734[7:6] == 2'h0 ? tag_1_11 : _GEN_2091; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2384 = _GEN_734[7:6] == 2'h0 ? tag_1_12 : _GEN_2092; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2385 = _GEN_734[7:6] == 2'h0 ? tag_1_13 : _GEN_2093; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2386 = _GEN_734[7:6] == 2'h0 ? tag_1_14 : _GEN_2094; // @[d_cache.scala 193:46 25:24]
  wire [31:0] _GEN_2387 = _GEN_734[7:6] == 2'h0 ? tag_1_15 : _GEN_2095; // @[d_cache.scala 193:46 25:24]
  wire  _GEN_2388 = _GEN_734[7:6] == 2'h0 ? dirty_1_0 : _GEN_2096; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2389 = _GEN_734[7:6] == 2'h0 ? dirty_1_1 : _GEN_2097; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2390 = _GEN_734[7:6] == 2'h0 ? dirty_1_2 : _GEN_2098; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2391 = _GEN_734[7:6] == 2'h0 ? dirty_1_3 : _GEN_2099; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2392 = _GEN_734[7:6] == 2'h0 ? dirty_1_4 : _GEN_2100; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2393 = _GEN_734[7:6] == 2'h0 ? dirty_1_5 : _GEN_2101; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2394 = _GEN_734[7:6] == 2'h0 ? dirty_1_6 : _GEN_2102; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2395 = _GEN_734[7:6] == 2'h0 ? dirty_1_7 : _GEN_2103; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2396 = _GEN_734[7:6] == 2'h0 ? dirty_1_8 : _GEN_2104; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2397 = _GEN_734[7:6] == 2'h0 ? dirty_1_9 : _GEN_2105; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2398 = _GEN_734[7:6] == 2'h0 ? dirty_1_10 : _GEN_2106; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2399 = _GEN_734[7:6] == 2'h0 ? dirty_1_11 : _GEN_2107; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2400 = _GEN_734[7:6] == 2'h0 ? dirty_1_12 : _GEN_2108; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2401 = _GEN_734[7:6] == 2'h0 ? dirty_1_13 : _GEN_2109; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2402 = _GEN_734[7:6] == 2'h0 ? dirty_1_14 : _GEN_2110; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2403 = _GEN_734[7:6] == 2'h0 ? dirty_1_15 : _GEN_2111; // @[d_cache.scala 193:46 35:26]
  wire  _GEN_2404 = _GEN_734[7:6] == 2'h0 ? valid_1_0 : _GEN_2112; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2405 = _GEN_734[7:6] == 2'h0 ? valid_1_1 : _GEN_2113; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2406 = _GEN_734[7:6] == 2'h0 ? valid_1_2 : _GEN_2114; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2407 = _GEN_734[7:6] == 2'h0 ? valid_1_3 : _GEN_2115; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2408 = _GEN_734[7:6] == 2'h0 ? valid_1_4 : _GEN_2116; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2409 = _GEN_734[7:6] == 2'h0 ? valid_1_5 : _GEN_2117; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2410 = _GEN_734[7:6] == 2'h0 ? valid_1_6 : _GEN_2118; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2411 = _GEN_734[7:6] == 2'h0 ? valid_1_7 : _GEN_2119; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2412 = _GEN_734[7:6] == 2'h0 ? valid_1_8 : _GEN_2120; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2413 = _GEN_734[7:6] == 2'h0 ? valid_1_9 : _GEN_2121; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2414 = _GEN_734[7:6] == 2'h0 ? valid_1_10 : _GEN_2122; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2415 = _GEN_734[7:6] == 2'h0 ? valid_1_11 : _GEN_2123; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2416 = _GEN_734[7:6] == 2'h0 ? valid_1_12 : _GEN_2124; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2417 = _GEN_734[7:6] == 2'h0 ? valid_1_13 : _GEN_2125; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2418 = _GEN_734[7:6] == 2'h0 ? valid_1_14 : _GEN_2126; // @[d_cache.scala 193:46 30:26]
  wire  _GEN_2419 = _GEN_734[7:6] == 2'h0 ? valid_1_15 : _GEN_2127; // @[d_cache.scala 193:46 30:26]
  wire [511:0] _GEN_2420 = _GEN_734[7:6] == 2'h0 ? ram_2_0 : _GEN_2145; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2421 = _GEN_734[7:6] == 2'h0 ? ram_2_1 : _GEN_2146; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2422 = _GEN_734[7:6] == 2'h0 ? ram_2_2 : _GEN_2147; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2423 = _GEN_734[7:6] == 2'h0 ? ram_2_3 : _GEN_2148; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2424 = _GEN_734[7:6] == 2'h0 ? ram_2_4 : _GEN_2149; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2425 = _GEN_734[7:6] == 2'h0 ? ram_2_5 : _GEN_2150; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2426 = _GEN_734[7:6] == 2'h0 ? ram_2_6 : _GEN_2151; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2427 = _GEN_734[7:6] == 2'h0 ? ram_2_7 : _GEN_2152; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2428 = _GEN_734[7:6] == 2'h0 ? ram_2_8 : _GEN_2153; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2429 = _GEN_734[7:6] == 2'h0 ? ram_2_9 : _GEN_2154; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2430 = _GEN_734[7:6] == 2'h0 ? ram_2_10 : _GEN_2155; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2431 = _GEN_734[7:6] == 2'h0 ? ram_2_11 : _GEN_2156; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2432 = _GEN_734[7:6] == 2'h0 ? ram_2_12 : _GEN_2157; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2433 = _GEN_734[7:6] == 2'h0 ? ram_2_13 : _GEN_2158; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2434 = _GEN_734[7:6] == 2'h0 ? ram_2_14 : _GEN_2159; // @[d_cache.scala 193:46 21:24]
  wire [511:0] _GEN_2435 = _GEN_734[7:6] == 2'h0 ? ram_2_15 : _GEN_2160; // @[d_cache.scala 193:46 21:24]
  wire [31:0] _GEN_2436 = _GEN_734[7:6] == 2'h0 ? tag_2_0 : _GEN_2161; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2437 = _GEN_734[7:6] == 2'h0 ? tag_2_1 : _GEN_2162; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2438 = _GEN_734[7:6] == 2'h0 ? tag_2_2 : _GEN_2163; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2439 = _GEN_734[7:6] == 2'h0 ? tag_2_3 : _GEN_2164; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2440 = _GEN_734[7:6] == 2'h0 ? tag_2_4 : _GEN_2165; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2441 = _GEN_734[7:6] == 2'h0 ? tag_2_5 : _GEN_2166; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2442 = _GEN_734[7:6] == 2'h0 ? tag_2_6 : _GEN_2167; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2443 = _GEN_734[7:6] == 2'h0 ? tag_2_7 : _GEN_2168; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2444 = _GEN_734[7:6] == 2'h0 ? tag_2_8 : _GEN_2169; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2445 = _GEN_734[7:6] == 2'h0 ? tag_2_9 : _GEN_2170; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2446 = _GEN_734[7:6] == 2'h0 ? tag_2_10 : _GEN_2171; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2447 = _GEN_734[7:6] == 2'h0 ? tag_2_11 : _GEN_2172; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2448 = _GEN_734[7:6] == 2'h0 ? tag_2_12 : _GEN_2173; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2449 = _GEN_734[7:6] == 2'h0 ? tag_2_13 : _GEN_2174; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2450 = _GEN_734[7:6] == 2'h0 ? tag_2_14 : _GEN_2175; // @[d_cache.scala 193:46 26:24]
  wire [31:0] _GEN_2451 = _GEN_734[7:6] == 2'h0 ? tag_2_15 : _GEN_2176; // @[d_cache.scala 193:46 26:24]
  wire  _GEN_2452 = _GEN_734[7:6] == 2'h0 ? dirty_2_0 : _GEN_2177; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2453 = _GEN_734[7:6] == 2'h0 ? dirty_2_1 : _GEN_2178; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2454 = _GEN_734[7:6] == 2'h0 ? dirty_2_2 : _GEN_2179; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2455 = _GEN_734[7:6] == 2'h0 ? dirty_2_3 : _GEN_2180; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2456 = _GEN_734[7:6] == 2'h0 ? dirty_2_4 : _GEN_2181; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2457 = _GEN_734[7:6] == 2'h0 ? dirty_2_5 : _GEN_2182; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2458 = _GEN_734[7:6] == 2'h0 ? dirty_2_6 : _GEN_2183; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2459 = _GEN_734[7:6] == 2'h0 ? dirty_2_7 : _GEN_2184; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2460 = _GEN_734[7:6] == 2'h0 ? dirty_2_8 : _GEN_2185; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2461 = _GEN_734[7:6] == 2'h0 ? dirty_2_9 : _GEN_2186; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2462 = _GEN_734[7:6] == 2'h0 ? dirty_2_10 : _GEN_2187; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2463 = _GEN_734[7:6] == 2'h0 ? dirty_2_11 : _GEN_2188; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2464 = _GEN_734[7:6] == 2'h0 ? dirty_2_12 : _GEN_2189; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2465 = _GEN_734[7:6] == 2'h0 ? dirty_2_13 : _GEN_2190; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2466 = _GEN_734[7:6] == 2'h0 ? dirty_2_14 : _GEN_2191; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2467 = _GEN_734[7:6] == 2'h0 ? dirty_2_15 : _GEN_2192; // @[d_cache.scala 193:46 36:26]
  wire  _GEN_2468 = _GEN_734[7:6] == 2'h0 ? valid_2_0 : _GEN_2193; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2469 = _GEN_734[7:6] == 2'h0 ? valid_2_1 : _GEN_2194; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2470 = _GEN_734[7:6] == 2'h0 ? valid_2_2 : _GEN_2195; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2471 = _GEN_734[7:6] == 2'h0 ? valid_2_3 : _GEN_2196; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2472 = _GEN_734[7:6] == 2'h0 ? valid_2_4 : _GEN_2197; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2473 = _GEN_734[7:6] == 2'h0 ? valid_2_5 : _GEN_2198; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2474 = _GEN_734[7:6] == 2'h0 ? valid_2_6 : _GEN_2199; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2475 = _GEN_734[7:6] == 2'h0 ? valid_2_7 : _GEN_2200; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2476 = _GEN_734[7:6] == 2'h0 ? valid_2_8 : _GEN_2201; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2477 = _GEN_734[7:6] == 2'h0 ? valid_2_9 : _GEN_2202; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2478 = _GEN_734[7:6] == 2'h0 ? valid_2_10 : _GEN_2203; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2479 = _GEN_734[7:6] == 2'h0 ? valid_2_11 : _GEN_2204; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2480 = _GEN_734[7:6] == 2'h0 ? valid_2_12 : _GEN_2205; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2481 = _GEN_734[7:6] == 2'h0 ? valid_2_13 : _GEN_2206; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2482 = _GEN_734[7:6] == 2'h0 ? valid_2_14 : _GEN_2207; // @[d_cache.scala 193:46 31:26]
  wire  _GEN_2483 = _GEN_734[7:6] == 2'h0 ? valid_2_15 : _GEN_2208; // @[d_cache.scala 193:46 31:26]
  wire [511:0] _GEN_2484 = _GEN_734[7:6] == 2'h0 ? ram_3_0 : _GEN_2209; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2485 = _GEN_734[7:6] == 2'h0 ? ram_3_1 : _GEN_2210; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2486 = _GEN_734[7:6] == 2'h0 ? ram_3_2 : _GEN_2211; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2487 = _GEN_734[7:6] == 2'h0 ? ram_3_3 : _GEN_2212; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2488 = _GEN_734[7:6] == 2'h0 ? ram_3_4 : _GEN_2213; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2489 = _GEN_734[7:6] == 2'h0 ? ram_3_5 : _GEN_2214; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2490 = _GEN_734[7:6] == 2'h0 ? ram_3_6 : _GEN_2215; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2491 = _GEN_734[7:6] == 2'h0 ? ram_3_7 : _GEN_2216; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2492 = _GEN_734[7:6] == 2'h0 ? ram_3_8 : _GEN_2217; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2493 = _GEN_734[7:6] == 2'h0 ? ram_3_9 : _GEN_2218; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2494 = _GEN_734[7:6] == 2'h0 ? ram_3_10 : _GEN_2219; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2495 = _GEN_734[7:6] == 2'h0 ? ram_3_11 : _GEN_2220; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2496 = _GEN_734[7:6] == 2'h0 ? ram_3_12 : _GEN_2221; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2497 = _GEN_734[7:6] == 2'h0 ? ram_3_13 : _GEN_2222; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2498 = _GEN_734[7:6] == 2'h0 ? ram_3_14 : _GEN_2223; // @[d_cache.scala 193:46 22:24]
  wire [511:0] _GEN_2499 = _GEN_734[7:6] == 2'h0 ? ram_3_15 : _GEN_2224; // @[d_cache.scala 193:46 22:24]
  wire [31:0] _GEN_2500 = _GEN_734[7:6] == 2'h0 ? tag_3_0 : _GEN_2225; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2501 = _GEN_734[7:6] == 2'h0 ? tag_3_1 : _GEN_2226; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2502 = _GEN_734[7:6] == 2'h0 ? tag_3_2 : _GEN_2227; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2503 = _GEN_734[7:6] == 2'h0 ? tag_3_3 : _GEN_2228; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2504 = _GEN_734[7:6] == 2'h0 ? tag_3_4 : _GEN_2229; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2505 = _GEN_734[7:6] == 2'h0 ? tag_3_5 : _GEN_2230; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2506 = _GEN_734[7:6] == 2'h0 ? tag_3_6 : _GEN_2231; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2507 = _GEN_734[7:6] == 2'h0 ? tag_3_7 : _GEN_2232; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2508 = _GEN_734[7:6] == 2'h0 ? tag_3_8 : _GEN_2233; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2509 = _GEN_734[7:6] == 2'h0 ? tag_3_9 : _GEN_2234; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2510 = _GEN_734[7:6] == 2'h0 ? tag_3_10 : _GEN_2235; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2511 = _GEN_734[7:6] == 2'h0 ? tag_3_11 : _GEN_2236; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2512 = _GEN_734[7:6] == 2'h0 ? tag_3_12 : _GEN_2237; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2513 = _GEN_734[7:6] == 2'h0 ? tag_3_13 : _GEN_2238; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2514 = _GEN_734[7:6] == 2'h0 ? tag_3_14 : _GEN_2239; // @[d_cache.scala 193:46 27:24]
  wire [31:0] _GEN_2515 = _GEN_734[7:6] == 2'h0 ? tag_3_15 : _GEN_2240; // @[d_cache.scala 193:46 27:24]
  wire  _GEN_2516 = _GEN_734[7:6] == 2'h0 ? dirty_3_0 : _GEN_2241; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2517 = _GEN_734[7:6] == 2'h0 ? dirty_3_1 : _GEN_2242; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2518 = _GEN_734[7:6] == 2'h0 ? dirty_3_2 : _GEN_2243; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2519 = _GEN_734[7:6] == 2'h0 ? dirty_3_3 : _GEN_2244; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2520 = _GEN_734[7:6] == 2'h0 ? dirty_3_4 : _GEN_2245; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2521 = _GEN_734[7:6] == 2'h0 ? dirty_3_5 : _GEN_2246; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2522 = _GEN_734[7:6] == 2'h0 ? dirty_3_6 : _GEN_2247; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2523 = _GEN_734[7:6] == 2'h0 ? dirty_3_7 : _GEN_2248; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2524 = _GEN_734[7:6] == 2'h0 ? dirty_3_8 : _GEN_2249; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2525 = _GEN_734[7:6] == 2'h0 ? dirty_3_9 : _GEN_2250; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2526 = _GEN_734[7:6] == 2'h0 ? dirty_3_10 : _GEN_2251; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2527 = _GEN_734[7:6] == 2'h0 ? dirty_3_11 : _GEN_2252; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2528 = _GEN_734[7:6] == 2'h0 ? dirty_3_12 : _GEN_2253; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2529 = _GEN_734[7:6] == 2'h0 ? dirty_3_13 : _GEN_2254; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2530 = _GEN_734[7:6] == 2'h0 ? dirty_3_14 : _GEN_2255; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2531 = _GEN_734[7:6] == 2'h0 ? dirty_3_15 : _GEN_2256; // @[d_cache.scala 193:46 37:26]
  wire  _GEN_2532 = _GEN_734[7:6] == 2'h0 ? valid_3_0 : _GEN_2257; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2533 = _GEN_734[7:6] == 2'h0 ? valid_3_1 : _GEN_2258; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2534 = _GEN_734[7:6] == 2'h0 ? valid_3_2 : _GEN_2259; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2535 = _GEN_734[7:6] == 2'h0 ? valid_3_3 : _GEN_2260; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2536 = _GEN_734[7:6] == 2'h0 ? valid_3_4 : _GEN_2261; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2537 = _GEN_734[7:6] == 2'h0 ? valid_3_5 : _GEN_2262; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2538 = _GEN_734[7:6] == 2'h0 ? valid_3_6 : _GEN_2263; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2539 = _GEN_734[7:6] == 2'h0 ? valid_3_7 : _GEN_2264; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2540 = _GEN_734[7:6] == 2'h0 ? valid_3_8 : _GEN_2265; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2541 = _GEN_734[7:6] == 2'h0 ? valid_3_9 : _GEN_2266; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2542 = _GEN_734[7:6] == 2'h0 ? valid_3_10 : _GEN_2267; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2543 = _GEN_734[7:6] == 2'h0 ? valid_3_11 : _GEN_2268; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2544 = _GEN_734[7:6] == 2'h0 ? valid_3_12 : _GEN_2269; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2545 = _GEN_734[7:6] == 2'h0 ? valid_3_13 : _GEN_2270; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2546 = _GEN_734[7:6] == 2'h0 ? valid_3_14 : _GEN_2271; // @[d_cache.scala 193:46 32:26]
  wire  _GEN_2547 = _GEN_734[7:6] == 2'h0 ? valid_3_15 : _GEN_2272; // @[d_cache.scala 193:46 32:26]
  wire [3:0] _GEN_2548 = unuse_way == 3'h4 ? 4'h1 : _GEN_2339; // @[d_cache.scala 186:40 187:23]
  wire [511:0] _GEN_2549 = unuse_way == 3'h4 ? _GEN_879 : _GEN_2484; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2550 = unuse_way == 3'h4 ? _GEN_880 : _GEN_2485; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2551 = unuse_way == 3'h4 ? _GEN_881 : _GEN_2486; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2552 = unuse_way == 3'h4 ? _GEN_882 : _GEN_2487; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2553 = unuse_way == 3'h4 ? _GEN_883 : _GEN_2488; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2554 = unuse_way == 3'h4 ? _GEN_884 : _GEN_2489; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2555 = unuse_way == 3'h4 ? _GEN_885 : _GEN_2490; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2556 = unuse_way == 3'h4 ? _GEN_886 : _GEN_2491; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2557 = unuse_way == 3'h4 ? _GEN_887 : _GEN_2492; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2558 = unuse_way == 3'h4 ? _GEN_888 : _GEN_2493; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2559 = unuse_way == 3'h4 ? _GEN_889 : _GEN_2494; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2560 = unuse_way == 3'h4 ? _GEN_890 : _GEN_2495; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2561 = unuse_way == 3'h4 ? _GEN_891 : _GEN_2496; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2562 = unuse_way == 3'h4 ? _GEN_892 : _GEN_2497; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2563 = unuse_way == 3'h4 ? _GEN_893 : _GEN_2498; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2564 = unuse_way == 3'h4 ? _GEN_894 : _GEN_2499; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2565 = unuse_way == 3'h4 ? _GEN_895 : _GEN_2500; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2566 = unuse_way == 3'h4 ? _GEN_896 : _GEN_2501; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2567 = unuse_way == 3'h4 ? _GEN_897 : _GEN_2502; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2568 = unuse_way == 3'h4 ? _GEN_898 : _GEN_2503; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2569 = unuse_way == 3'h4 ? _GEN_899 : _GEN_2504; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2570 = unuse_way == 3'h4 ? _GEN_900 : _GEN_2505; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2571 = unuse_way == 3'h4 ? _GEN_901 : _GEN_2506; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2572 = unuse_way == 3'h4 ? _GEN_902 : _GEN_2507; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2573 = unuse_way == 3'h4 ? _GEN_903 : _GEN_2508; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2574 = unuse_way == 3'h4 ? _GEN_904 : _GEN_2509; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2575 = unuse_way == 3'h4 ? _GEN_905 : _GEN_2510; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2576 = unuse_way == 3'h4 ? _GEN_906 : _GEN_2511; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2577 = unuse_way == 3'h4 ? _GEN_907 : _GEN_2512; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2578 = unuse_way == 3'h4 ? _GEN_908 : _GEN_2513; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2579 = unuse_way == 3'h4 ? _GEN_909 : _GEN_2514; // @[d_cache.scala 186:40]
  wire [31:0] _GEN_2580 = unuse_way == 3'h4 ? _GEN_910 : _GEN_2515; // @[d_cache.scala 186:40]
  wire  _GEN_2581 = unuse_way == 3'h4 ? _GEN_911 : _GEN_2532; // @[d_cache.scala 186:40]
  wire  _GEN_2582 = unuse_way == 3'h4 ? _GEN_912 : _GEN_2533; // @[d_cache.scala 186:40]
  wire  _GEN_2583 = unuse_way == 3'h4 ? _GEN_913 : _GEN_2534; // @[d_cache.scala 186:40]
  wire  _GEN_2584 = unuse_way == 3'h4 ? _GEN_914 : _GEN_2535; // @[d_cache.scala 186:40]
  wire  _GEN_2585 = unuse_way == 3'h4 ? _GEN_915 : _GEN_2536; // @[d_cache.scala 186:40]
  wire  _GEN_2586 = unuse_way == 3'h4 ? _GEN_916 : _GEN_2537; // @[d_cache.scala 186:40]
  wire  _GEN_2587 = unuse_way == 3'h4 ? _GEN_917 : _GEN_2538; // @[d_cache.scala 186:40]
  wire  _GEN_2588 = unuse_way == 3'h4 ? _GEN_918 : _GEN_2539; // @[d_cache.scala 186:40]
  wire  _GEN_2589 = unuse_way == 3'h4 ? _GEN_919 : _GEN_2540; // @[d_cache.scala 186:40]
  wire  _GEN_2590 = unuse_way == 3'h4 ? _GEN_920 : _GEN_2541; // @[d_cache.scala 186:40]
  wire  _GEN_2591 = unuse_way == 3'h4 ? _GEN_921 : _GEN_2542; // @[d_cache.scala 186:40]
  wire  _GEN_2592 = unuse_way == 3'h4 ? _GEN_922 : _GEN_2543; // @[d_cache.scala 186:40]
  wire  _GEN_2593 = unuse_way == 3'h4 ? _GEN_923 : _GEN_2544; // @[d_cache.scala 186:40]
  wire  _GEN_2594 = unuse_way == 3'h4 ? _GEN_924 : _GEN_2545; // @[d_cache.scala 186:40]
  wire  _GEN_2595 = unuse_way == 3'h4 ? _GEN_925 : _GEN_2546; // @[d_cache.scala 186:40]
  wire  _GEN_2596 = unuse_way == 3'h4 ? _GEN_926 : _GEN_2547; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2597 = unuse_way == 3'h4 ? _GEN_927 : _GEN_2340; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2598 = unuse_way == 3'h4 ? _GEN_928 : _GEN_2341; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2599 = unuse_way == 3'h4 ? _GEN_929 : _GEN_2342; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2600 = unuse_way == 3'h4 ? _GEN_930 : _GEN_2343; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2601 = unuse_way == 3'h4 ? _GEN_931 : _GEN_2344; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2602 = unuse_way == 3'h4 ? _GEN_932 : _GEN_2345; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2603 = unuse_way == 3'h4 ? _GEN_933 : _GEN_2346; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2604 = unuse_way == 3'h4 ? _GEN_934 : _GEN_2347; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2605 = unuse_way == 3'h4 ? _GEN_935 : _GEN_2348; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2606 = unuse_way == 3'h4 ? _GEN_936 : _GEN_2349; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2607 = unuse_way == 3'h4 ? _GEN_937 : _GEN_2350; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2608 = unuse_way == 3'h4 ? _GEN_938 : _GEN_2351; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2609 = unuse_way == 3'h4 ? _GEN_939 : _GEN_2352; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2610 = unuse_way == 3'h4 ? _GEN_940 : _GEN_2353; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2611 = unuse_way == 3'h4 ? _GEN_941 : _GEN_2354; // @[d_cache.scala 186:40]
  wire [7:0] _GEN_2612 = unuse_way == 3'h4 ? _GEN_942 : _GEN_2355; // @[d_cache.scala 186:40]
  wire [511:0] _GEN_2613 = unuse_way == 3'h4 ? write_back_data : _GEN_2273; // @[d_cache.scala 186:40 44:34]
  wire [41:0] _GEN_2614 = unuse_way == 3'h4 ? {{10'd0}, write_back_addr} : _GEN_2274; // @[d_cache.scala 186:40 45:34]
  wire [511:0] _GEN_2615 = unuse_way == 3'h4 ? ram_0_0 : _GEN_2275; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2616 = unuse_way == 3'h4 ? ram_0_1 : _GEN_2276; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2617 = unuse_way == 3'h4 ? ram_0_2 : _GEN_2277; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2618 = unuse_way == 3'h4 ? ram_0_3 : _GEN_2278; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2619 = unuse_way == 3'h4 ? ram_0_4 : _GEN_2279; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2620 = unuse_way == 3'h4 ? ram_0_5 : _GEN_2280; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2621 = unuse_way == 3'h4 ? ram_0_6 : _GEN_2281; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2622 = unuse_way == 3'h4 ? ram_0_7 : _GEN_2282; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2623 = unuse_way == 3'h4 ? ram_0_8 : _GEN_2283; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2624 = unuse_way == 3'h4 ? ram_0_9 : _GEN_2284; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2625 = unuse_way == 3'h4 ? ram_0_10 : _GEN_2285; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2626 = unuse_way == 3'h4 ? ram_0_11 : _GEN_2286; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2627 = unuse_way == 3'h4 ? ram_0_12 : _GEN_2287; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2628 = unuse_way == 3'h4 ? ram_0_13 : _GEN_2288; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2629 = unuse_way == 3'h4 ? ram_0_14 : _GEN_2289; // @[d_cache.scala 186:40 19:24]
  wire [511:0] _GEN_2630 = unuse_way == 3'h4 ? ram_0_15 : _GEN_2290; // @[d_cache.scala 186:40 19:24]
  wire [31:0] _GEN_2631 = unuse_way == 3'h4 ? tag_0_0 : _GEN_2291; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2632 = unuse_way == 3'h4 ? tag_0_1 : _GEN_2292; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2633 = unuse_way == 3'h4 ? tag_0_2 : _GEN_2293; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2634 = unuse_way == 3'h4 ? tag_0_3 : _GEN_2294; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2635 = unuse_way == 3'h4 ? tag_0_4 : _GEN_2295; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2636 = unuse_way == 3'h4 ? tag_0_5 : _GEN_2296; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2637 = unuse_way == 3'h4 ? tag_0_6 : _GEN_2297; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2638 = unuse_way == 3'h4 ? tag_0_7 : _GEN_2298; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2639 = unuse_way == 3'h4 ? tag_0_8 : _GEN_2299; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2640 = unuse_way == 3'h4 ? tag_0_9 : _GEN_2300; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2641 = unuse_way == 3'h4 ? tag_0_10 : _GEN_2301; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2642 = unuse_way == 3'h4 ? tag_0_11 : _GEN_2302; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2643 = unuse_way == 3'h4 ? tag_0_12 : _GEN_2303; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2644 = unuse_way == 3'h4 ? tag_0_13 : _GEN_2304; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2645 = unuse_way == 3'h4 ? tag_0_14 : _GEN_2305; // @[d_cache.scala 186:40 24:24]
  wire [31:0] _GEN_2646 = unuse_way == 3'h4 ? tag_0_15 : _GEN_2306; // @[d_cache.scala 186:40 24:24]
  wire  _GEN_2647 = unuse_way == 3'h4 ? dirty_0_0 : _GEN_2307; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2648 = unuse_way == 3'h4 ? dirty_0_1 : _GEN_2308; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2649 = unuse_way == 3'h4 ? dirty_0_2 : _GEN_2309; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2650 = unuse_way == 3'h4 ? dirty_0_3 : _GEN_2310; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2651 = unuse_way == 3'h4 ? dirty_0_4 : _GEN_2311; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2652 = unuse_way == 3'h4 ? dirty_0_5 : _GEN_2312; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2653 = unuse_way == 3'h4 ? dirty_0_6 : _GEN_2313; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2654 = unuse_way == 3'h4 ? dirty_0_7 : _GEN_2314; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2655 = unuse_way == 3'h4 ? dirty_0_8 : _GEN_2315; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2656 = unuse_way == 3'h4 ? dirty_0_9 : _GEN_2316; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2657 = unuse_way == 3'h4 ? dirty_0_10 : _GEN_2317; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2658 = unuse_way == 3'h4 ? dirty_0_11 : _GEN_2318; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2659 = unuse_way == 3'h4 ? dirty_0_12 : _GEN_2319; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2660 = unuse_way == 3'h4 ? dirty_0_13 : _GEN_2320; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2661 = unuse_way == 3'h4 ? dirty_0_14 : _GEN_2321; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2662 = unuse_way == 3'h4 ? dirty_0_15 : _GEN_2322; // @[d_cache.scala 186:40 34:26]
  wire  _GEN_2663 = unuse_way == 3'h4 ? valid_0_0 : _GEN_2323; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2664 = unuse_way == 3'h4 ? valid_0_1 : _GEN_2324; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2665 = unuse_way == 3'h4 ? valid_0_2 : _GEN_2325; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2666 = unuse_way == 3'h4 ? valid_0_3 : _GEN_2326; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2667 = unuse_way == 3'h4 ? valid_0_4 : _GEN_2327; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2668 = unuse_way == 3'h4 ? valid_0_5 : _GEN_2328; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2669 = unuse_way == 3'h4 ? valid_0_6 : _GEN_2329; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2670 = unuse_way == 3'h4 ? valid_0_7 : _GEN_2330; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2671 = unuse_way == 3'h4 ? valid_0_8 : _GEN_2331; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2672 = unuse_way == 3'h4 ? valid_0_9 : _GEN_2332; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2673 = unuse_way == 3'h4 ? valid_0_10 : _GEN_2333; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2674 = unuse_way == 3'h4 ? valid_0_11 : _GEN_2334; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2675 = unuse_way == 3'h4 ? valid_0_12 : _GEN_2335; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2676 = unuse_way == 3'h4 ? valid_0_13 : _GEN_2336; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2677 = unuse_way == 3'h4 ? valid_0_14 : _GEN_2337; // @[d_cache.scala 186:40 29:26]
  wire  _GEN_2678 = unuse_way == 3'h4 ? valid_0_15 : _GEN_2338; // @[d_cache.scala 186:40 29:26]
  wire [511:0] _GEN_2679 = unuse_way == 3'h4 ? ram_1_0 : _GEN_2356; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2680 = unuse_way == 3'h4 ? ram_1_1 : _GEN_2357; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2681 = unuse_way == 3'h4 ? ram_1_2 : _GEN_2358; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2682 = unuse_way == 3'h4 ? ram_1_3 : _GEN_2359; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2683 = unuse_way == 3'h4 ? ram_1_4 : _GEN_2360; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2684 = unuse_way == 3'h4 ? ram_1_5 : _GEN_2361; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2685 = unuse_way == 3'h4 ? ram_1_6 : _GEN_2362; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2686 = unuse_way == 3'h4 ? ram_1_7 : _GEN_2363; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2687 = unuse_way == 3'h4 ? ram_1_8 : _GEN_2364; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2688 = unuse_way == 3'h4 ? ram_1_9 : _GEN_2365; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2689 = unuse_way == 3'h4 ? ram_1_10 : _GEN_2366; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2690 = unuse_way == 3'h4 ? ram_1_11 : _GEN_2367; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2691 = unuse_way == 3'h4 ? ram_1_12 : _GEN_2368; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2692 = unuse_way == 3'h4 ? ram_1_13 : _GEN_2369; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2693 = unuse_way == 3'h4 ? ram_1_14 : _GEN_2370; // @[d_cache.scala 186:40 20:24]
  wire [511:0] _GEN_2694 = unuse_way == 3'h4 ? ram_1_15 : _GEN_2371; // @[d_cache.scala 186:40 20:24]
  wire [31:0] _GEN_2695 = unuse_way == 3'h4 ? tag_1_0 : _GEN_2372; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2696 = unuse_way == 3'h4 ? tag_1_1 : _GEN_2373; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2697 = unuse_way == 3'h4 ? tag_1_2 : _GEN_2374; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2698 = unuse_way == 3'h4 ? tag_1_3 : _GEN_2375; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2699 = unuse_way == 3'h4 ? tag_1_4 : _GEN_2376; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2700 = unuse_way == 3'h4 ? tag_1_5 : _GEN_2377; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2701 = unuse_way == 3'h4 ? tag_1_6 : _GEN_2378; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2702 = unuse_way == 3'h4 ? tag_1_7 : _GEN_2379; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2703 = unuse_way == 3'h4 ? tag_1_8 : _GEN_2380; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2704 = unuse_way == 3'h4 ? tag_1_9 : _GEN_2381; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2705 = unuse_way == 3'h4 ? tag_1_10 : _GEN_2382; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2706 = unuse_way == 3'h4 ? tag_1_11 : _GEN_2383; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2707 = unuse_way == 3'h4 ? tag_1_12 : _GEN_2384; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2708 = unuse_way == 3'h4 ? tag_1_13 : _GEN_2385; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2709 = unuse_way == 3'h4 ? tag_1_14 : _GEN_2386; // @[d_cache.scala 186:40 25:24]
  wire [31:0] _GEN_2710 = unuse_way == 3'h4 ? tag_1_15 : _GEN_2387; // @[d_cache.scala 186:40 25:24]
  wire  _GEN_2711 = unuse_way == 3'h4 ? dirty_1_0 : _GEN_2388; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2712 = unuse_way == 3'h4 ? dirty_1_1 : _GEN_2389; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2713 = unuse_way == 3'h4 ? dirty_1_2 : _GEN_2390; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2714 = unuse_way == 3'h4 ? dirty_1_3 : _GEN_2391; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2715 = unuse_way == 3'h4 ? dirty_1_4 : _GEN_2392; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2716 = unuse_way == 3'h4 ? dirty_1_5 : _GEN_2393; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2717 = unuse_way == 3'h4 ? dirty_1_6 : _GEN_2394; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2718 = unuse_way == 3'h4 ? dirty_1_7 : _GEN_2395; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2719 = unuse_way == 3'h4 ? dirty_1_8 : _GEN_2396; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2720 = unuse_way == 3'h4 ? dirty_1_9 : _GEN_2397; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2721 = unuse_way == 3'h4 ? dirty_1_10 : _GEN_2398; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2722 = unuse_way == 3'h4 ? dirty_1_11 : _GEN_2399; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2723 = unuse_way == 3'h4 ? dirty_1_12 : _GEN_2400; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2724 = unuse_way == 3'h4 ? dirty_1_13 : _GEN_2401; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2725 = unuse_way == 3'h4 ? dirty_1_14 : _GEN_2402; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2726 = unuse_way == 3'h4 ? dirty_1_15 : _GEN_2403; // @[d_cache.scala 186:40 35:26]
  wire  _GEN_2727 = unuse_way == 3'h4 ? valid_1_0 : _GEN_2404; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2728 = unuse_way == 3'h4 ? valid_1_1 : _GEN_2405; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2729 = unuse_way == 3'h4 ? valid_1_2 : _GEN_2406; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2730 = unuse_way == 3'h4 ? valid_1_3 : _GEN_2407; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2731 = unuse_way == 3'h4 ? valid_1_4 : _GEN_2408; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2732 = unuse_way == 3'h4 ? valid_1_5 : _GEN_2409; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2733 = unuse_way == 3'h4 ? valid_1_6 : _GEN_2410; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2734 = unuse_way == 3'h4 ? valid_1_7 : _GEN_2411; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2735 = unuse_way == 3'h4 ? valid_1_8 : _GEN_2412; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2736 = unuse_way == 3'h4 ? valid_1_9 : _GEN_2413; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2737 = unuse_way == 3'h4 ? valid_1_10 : _GEN_2414; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2738 = unuse_way == 3'h4 ? valid_1_11 : _GEN_2415; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2739 = unuse_way == 3'h4 ? valid_1_12 : _GEN_2416; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2740 = unuse_way == 3'h4 ? valid_1_13 : _GEN_2417; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2741 = unuse_way == 3'h4 ? valid_1_14 : _GEN_2418; // @[d_cache.scala 186:40 30:26]
  wire  _GEN_2742 = unuse_way == 3'h4 ? valid_1_15 : _GEN_2419; // @[d_cache.scala 186:40 30:26]
  wire [511:0] _GEN_2743 = unuse_way == 3'h4 ? ram_2_0 : _GEN_2420; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2744 = unuse_way == 3'h4 ? ram_2_1 : _GEN_2421; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2745 = unuse_way == 3'h4 ? ram_2_2 : _GEN_2422; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2746 = unuse_way == 3'h4 ? ram_2_3 : _GEN_2423; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2747 = unuse_way == 3'h4 ? ram_2_4 : _GEN_2424; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2748 = unuse_way == 3'h4 ? ram_2_5 : _GEN_2425; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2749 = unuse_way == 3'h4 ? ram_2_6 : _GEN_2426; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2750 = unuse_way == 3'h4 ? ram_2_7 : _GEN_2427; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2751 = unuse_way == 3'h4 ? ram_2_8 : _GEN_2428; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2752 = unuse_way == 3'h4 ? ram_2_9 : _GEN_2429; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2753 = unuse_way == 3'h4 ? ram_2_10 : _GEN_2430; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2754 = unuse_way == 3'h4 ? ram_2_11 : _GEN_2431; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2755 = unuse_way == 3'h4 ? ram_2_12 : _GEN_2432; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2756 = unuse_way == 3'h4 ? ram_2_13 : _GEN_2433; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2757 = unuse_way == 3'h4 ? ram_2_14 : _GEN_2434; // @[d_cache.scala 186:40 21:24]
  wire [511:0] _GEN_2758 = unuse_way == 3'h4 ? ram_2_15 : _GEN_2435; // @[d_cache.scala 186:40 21:24]
  wire [31:0] _GEN_2759 = unuse_way == 3'h4 ? tag_2_0 : _GEN_2436; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2760 = unuse_way == 3'h4 ? tag_2_1 : _GEN_2437; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2761 = unuse_way == 3'h4 ? tag_2_2 : _GEN_2438; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2762 = unuse_way == 3'h4 ? tag_2_3 : _GEN_2439; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2763 = unuse_way == 3'h4 ? tag_2_4 : _GEN_2440; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2764 = unuse_way == 3'h4 ? tag_2_5 : _GEN_2441; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2765 = unuse_way == 3'h4 ? tag_2_6 : _GEN_2442; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2766 = unuse_way == 3'h4 ? tag_2_7 : _GEN_2443; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2767 = unuse_way == 3'h4 ? tag_2_8 : _GEN_2444; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2768 = unuse_way == 3'h4 ? tag_2_9 : _GEN_2445; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2769 = unuse_way == 3'h4 ? tag_2_10 : _GEN_2446; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2770 = unuse_way == 3'h4 ? tag_2_11 : _GEN_2447; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2771 = unuse_way == 3'h4 ? tag_2_12 : _GEN_2448; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2772 = unuse_way == 3'h4 ? tag_2_13 : _GEN_2449; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2773 = unuse_way == 3'h4 ? tag_2_14 : _GEN_2450; // @[d_cache.scala 186:40 26:24]
  wire [31:0] _GEN_2774 = unuse_way == 3'h4 ? tag_2_15 : _GEN_2451; // @[d_cache.scala 186:40 26:24]
  wire  _GEN_2775 = unuse_way == 3'h4 ? dirty_2_0 : _GEN_2452; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2776 = unuse_way == 3'h4 ? dirty_2_1 : _GEN_2453; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2777 = unuse_way == 3'h4 ? dirty_2_2 : _GEN_2454; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2778 = unuse_way == 3'h4 ? dirty_2_3 : _GEN_2455; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2779 = unuse_way == 3'h4 ? dirty_2_4 : _GEN_2456; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2780 = unuse_way == 3'h4 ? dirty_2_5 : _GEN_2457; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2781 = unuse_way == 3'h4 ? dirty_2_6 : _GEN_2458; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2782 = unuse_way == 3'h4 ? dirty_2_7 : _GEN_2459; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2783 = unuse_way == 3'h4 ? dirty_2_8 : _GEN_2460; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2784 = unuse_way == 3'h4 ? dirty_2_9 : _GEN_2461; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2785 = unuse_way == 3'h4 ? dirty_2_10 : _GEN_2462; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2786 = unuse_way == 3'h4 ? dirty_2_11 : _GEN_2463; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2787 = unuse_way == 3'h4 ? dirty_2_12 : _GEN_2464; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2788 = unuse_way == 3'h4 ? dirty_2_13 : _GEN_2465; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2789 = unuse_way == 3'h4 ? dirty_2_14 : _GEN_2466; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2790 = unuse_way == 3'h4 ? dirty_2_15 : _GEN_2467; // @[d_cache.scala 186:40 36:26]
  wire  _GEN_2791 = unuse_way == 3'h4 ? valid_2_0 : _GEN_2468; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2792 = unuse_way == 3'h4 ? valid_2_1 : _GEN_2469; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2793 = unuse_way == 3'h4 ? valid_2_2 : _GEN_2470; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2794 = unuse_way == 3'h4 ? valid_2_3 : _GEN_2471; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2795 = unuse_way == 3'h4 ? valid_2_4 : _GEN_2472; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2796 = unuse_way == 3'h4 ? valid_2_5 : _GEN_2473; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2797 = unuse_way == 3'h4 ? valid_2_6 : _GEN_2474; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2798 = unuse_way == 3'h4 ? valid_2_7 : _GEN_2475; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2799 = unuse_way == 3'h4 ? valid_2_8 : _GEN_2476; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2800 = unuse_way == 3'h4 ? valid_2_9 : _GEN_2477; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2801 = unuse_way == 3'h4 ? valid_2_10 : _GEN_2478; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2802 = unuse_way == 3'h4 ? valid_2_11 : _GEN_2479; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2803 = unuse_way == 3'h4 ? valid_2_12 : _GEN_2480; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2804 = unuse_way == 3'h4 ? valid_2_13 : _GEN_2481; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2805 = unuse_way == 3'h4 ? valid_2_14 : _GEN_2482; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2806 = unuse_way == 3'h4 ? valid_2_15 : _GEN_2483; // @[d_cache.scala 186:40 31:26]
  wire  _GEN_2807 = unuse_way == 3'h4 ? dirty_3_0 : _GEN_2516; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2808 = unuse_way == 3'h4 ? dirty_3_1 : _GEN_2517; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2809 = unuse_way == 3'h4 ? dirty_3_2 : _GEN_2518; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2810 = unuse_way == 3'h4 ? dirty_3_3 : _GEN_2519; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2811 = unuse_way == 3'h4 ? dirty_3_4 : _GEN_2520; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2812 = unuse_way == 3'h4 ? dirty_3_5 : _GEN_2521; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2813 = unuse_way == 3'h4 ? dirty_3_6 : _GEN_2522; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2814 = unuse_way == 3'h4 ? dirty_3_7 : _GEN_2523; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2815 = unuse_way == 3'h4 ? dirty_3_8 : _GEN_2524; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2816 = unuse_way == 3'h4 ? dirty_3_9 : _GEN_2525; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2817 = unuse_way == 3'h4 ? dirty_3_10 : _GEN_2526; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2818 = unuse_way == 3'h4 ? dirty_3_11 : _GEN_2527; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2819 = unuse_way == 3'h4 ? dirty_3_12 : _GEN_2528; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2820 = unuse_way == 3'h4 ? dirty_3_13 : _GEN_2529; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2821 = unuse_way == 3'h4 ? dirty_3_14 : _GEN_2530; // @[d_cache.scala 186:40 37:26]
  wire  _GEN_2822 = unuse_way == 3'h4 ? dirty_3_15 : _GEN_2531; // @[d_cache.scala 186:40 37:26]
  wire [3:0] _GEN_2823 = unuse_way == 3'h3 ? 4'h1 : _GEN_2548; // @[d_cache.scala 180:40 181:23]
  wire [511:0] _GEN_2824 = unuse_way == 3'h3 ? _GEN_815 : _GEN_2743; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2825 = unuse_way == 3'h3 ? _GEN_816 : _GEN_2744; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2826 = unuse_way == 3'h3 ? _GEN_817 : _GEN_2745; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2827 = unuse_way == 3'h3 ? _GEN_818 : _GEN_2746; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2828 = unuse_way == 3'h3 ? _GEN_819 : _GEN_2747; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2829 = unuse_way == 3'h3 ? _GEN_820 : _GEN_2748; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2830 = unuse_way == 3'h3 ? _GEN_821 : _GEN_2749; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2831 = unuse_way == 3'h3 ? _GEN_822 : _GEN_2750; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2832 = unuse_way == 3'h3 ? _GEN_823 : _GEN_2751; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2833 = unuse_way == 3'h3 ? _GEN_824 : _GEN_2752; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2834 = unuse_way == 3'h3 ? _GEN_825 : _GEN_2753; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2835 = unuse_way == 3'h3 ? _GEN_826 : _GEN_2754; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2836 = unuse_way == 3'h3 ? _GEN_827 : _GEN_2755; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2837 = unuse_way == 3'h3 ? _GEN_828 : _GEN_2756; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2838 = unuse_way == 3'h3 ? _GEN_829 : _GEN_2757; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2839 = unuse_way == 3'h3 ? _GEN_830 : _GEN_2758; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2840 = unuse_way == 3'h3 ? _GEN_831 : _GEN_2759; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2841 = unuse_way == 3'h3 ? _GEN_832 : _GEN_2760; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2842 = unuse_way == 3'h3 ? _GEN_833 : _GEN_2761; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2843 = unuse_way == 3'h3 ? _GEN_834 : _GEN_2762; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2844 = unuse_way == 3'h3 ? _GEN_835 : _GEN_2763; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2845 = unuse_way == 3'h3 ? _GEN_836 : _GEN_2764; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2846 = unuse_way == 3'h3 ? _GEN_837 : _GEN_2765; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2847 = unuse_way == 3'h3 ? _GEN_838 : _GEN_2766; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2848 = unuse_way == 3'h3 ? _GEN_839 : _GEN_2767; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2849 = unuse_way == 3'h3 ? _GEN_840 : _GEN_2768; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2850 = unuse_way == 3'h3 ? _GEN_841 : _GEN_2769; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2851 = unuse_way == 3'h3 ? _GEN_842 : _GEN_2770; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2852 = unuse_way == 3'h3 ? _GEN_843 : _GEN_2771; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2853 = unuse_way == 3'h3 ? _GEN_844 : _GEN_2772; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2854 = unuse_way == 3'h3 ? _GEN_845 : _GEN_2773; // @[d_cache.scala 180:40]
  wire [31:0] _GEN_2855 = unuse_way == 3'h3 ? _GEN_846 : _GEN_2774; // @[d_cache.scala 180:40]
  wire  _GEN_2856 = unuse_way == 3'h3 ? _GEN_847 : _GEN_2791; // @[d_cache.scala 180:40]
  wire  _GEN_2857 = unuse_way == 3'h3 ? _GEN_848 : _GEN_2792; // @[d_cache.scala 180:40]
  wire  _GEN_2858 = unuse_way == 3'h3 ? _GEN_849 : _GEN_2793; // @[d_cache.scala 180:40]
  wire  _GEN_2859 = unuse_way == 3'h3 ? _GEN_850 : _GEN_2794; // @[d_cache.scala 180:40]
  wire  _GEN_2860 = unuse_way == 3'h3 ? _GEN_851 : _GEN_2795; // @[d_cache.scala 180:40]
  wire  _GEN_2861 = unuse_way == 3'h3 ? _GEN_852 : _GEN_2796; // @[d_cache.scala 180:40]
  wire  _GEN_2862 = unuse_way == 3'h3 ? _GEN_853 : _GEN_2797; // @[d_cache.scala 180:40]
  wire  _GEN_2863 = unuse_way == 3'h3 ? _GEN_854 : _GEN_2798; // @[d_cache.scala 180:40]
  wire  _GEN_2864 = unuse_way == 3'h3 ? _GEN_855 : _GEN_2799; // @[d_cache.scala 180:40]
  wire  _GEN_2865 = unuse_way == 3'h3 ? _GEN_856 : _GEN_2800; // @[d_cache.scala 180:40]
  wire  _GEN_2866 = unuse_way == 3'h3 ? _GEN_857 : _GEN_2801; // @[d_cache.scala 180:40]
  wire  _GEN_2867 = unuse_way == 3'h3 ? _GEN_858 : _GEN_2802; // @[d_cache.scala 180:40]
  wire  _GEN_2868 = unuse_way == 3'h3 ? _GEN_859 : _GEN_2803; // @[d_cache.scala 180:40]
  wire  _GEN_2869 = unuse_way == 3'h3 ? _GEN_860 : _GEN_2804; // @[d_cache.scala 180:40]
  wire  _GEN_2870 = unuse_way == 3'h3 ? _GEN_861 : _GEN_2805; // @[d_cache.scala 180:40]
  wire  _GEN_2871 = unuse_way == 3'h3 ? _GEN_862 : _GEN_2806; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2872 = unuse_way == 3'h3 ? _GEN_863 : _GEN_2597; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2873 = unuse_way == 3'h3 ? _GEN_864 : _GEN_2598; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2874 = unuse_way == 3'h3 ? _GEN_865 : _GEN_2599; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2875 = unuse_way == 3'h3 ? _GEN_866 : _GEN_2600; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2876 = unuse_way == 3'h3 ? _GEN_867 : _GEN_2601; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2877 = unuse_way == 3'h3 ? _GEN_868 : _GEN_2602; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2878 = unuse_way == 3'h3 ? _GEN_869 : _GEN_2603; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2879 = unuse_way == 3'h3 ? _GEN_870 : _GEN_2604; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2880 = unuse_way == 3'h3 ? _GEN_871 : _GEN_2605; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2881 = unuse_way == 3'h3 ? _GEN_872 : _GEN_2606; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2882 = unuse_way == 3'h3 ? _GEN_873 : _GEN_2607; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2883 = unuse_way == 3'h3 ? _GEN_874 : _GEN_2608; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2884 = unuse_way == 3'h3 ? _GEN_875 : _GEN_2609; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2885 = unuse_way == 3'h3 ? _GEN_876 : _GEN_2610; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2886 = unuse_way == 3'h3 ? _GEN_877 : _GEN_2611; // @[d_cache.scala 180:40]
  wire [7:0] _GEN_2887 = unuse_way == 3'h3 ? _GEN_878 : _GEN_2612; // @[d_cache.scala 180:40]
  wire [511:0] _GEN_2888 = unuse_way == 3'h3 ? ram_3_0 : _GEN_2549; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2889 = unuse_way == 3'h3 ? ram_3_1 : _GEN_2550; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2890 = unuse_way == 3'h3 ? ram_3_2 : _GEN_2551; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2891 = unuse_way == 3'h3 ? ram_3_3 : _GEN_2552; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2892 = unuse_way == 3'h3 ? ram_3_4 : _GEN_2553; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2893 = unuse_way == 3'h3 ? ram_3_5 : _GEN_2554; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2894 = unuse_way == 3'h3 ? ram_3_6 : _GEN_2555; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2895 = unuse_way == 3'h3 ? ram_3_7 : _GEN_2556; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2896 = unuse_way == 3'h3 ? ram_3_8 : _GEN_2557; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2897 = unuse_way == 3'h3 ? ram_3_9 : _GEN_2558; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2898 = unuse_way == 3'h3 ? ram_3_10 : _GEN_2559; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2899 = unuse_way == 3'h3 ? ram_3_11 : _GEN_2560; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2900 = unuse_way == 3'h3 ? ram_3_12 : _GEN_2561; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2901 = unuse_way == 3'h3 ? ram_3_13 : _GEN_2562; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2902 = unuse_way == 3'h3 ? ram_3_14 : _GEN_2563; // @[d_cache.scala 180:40 22:24]
  wire [511:0] _GEN_2903 = unuse_way == 3'h3 ? ram_3_15 : _GEN_2564; // @[d_cache.scala 180:40 22:24]
  wire [31:0] _GEN_2904 = unuse_way == 3'h3 ? tag_3_0 : _GEN_2565; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2905 = unuse_way == 3'h3 ? tag_3_1 : _GEN_2566; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2906 = unuse_way == 3'h3 ? tag_3_2 : _GEN_2567; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2907 = unuse_way == 3'h3 ? tag_3_3 : _GEN_2568; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2908 = unuse_way == 3'h3 ? tag_3_4 : _GEN_2569; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2909 = unuse_way == 3'h3 ? tag_3_5 : _GEN_2570; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2910 = unuse_way == 3'h3 ? tag_3_6 : _GEN_2571; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2911 = unuse_way == 3'h3 ? tag_3_7 : _GEN_2572; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2912 = unuse_way == 3'h3 ? tag_3_8 : _GEN_2573; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2913 = unuse_way == 3'h3 ? tag_3_9 : _GEN_2574; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2914 = unuse_way == 3'h3 ? tag_3_10 : _GEN_2575; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2915 = unuse_way == 3'h3 ? tag_3_11 : _GEN_2576; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2916 = unuse_way == 3'h3 ? tag_3_12 : _GEN_2577; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2917 = unuse_way == 3'h3 ? tag_3_13 : _GEN_2578; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2918 = unuse_way == 3'h3 ? tag_3_14 : _GEN_2579; // @[d_cache.scala 180:40 27:24]
  wire [31:0] _GEN_2919 = unuse_way == 3'h3 ? tag_3_15 : _GEN_2580; // @[d_cache.scala 180:40 27:24]
  wire  _GEN_2920 = unuse_way == 3'h3 ? valid_3_0 : _GEN_2581; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2921 = unuse_way == 3'h3 ? valid_3_1 : _GEN_2582; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2922 = unuse_way == 3'h3 ? valid_3_2 : _GEN_2583; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2923 = unuse_way == 3'h3 ? valid_3_3 : _GEN_2584; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2924 = unuse_way == 3'h3 ? valid_3_4 : _GEN_2585; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2925 = unuse_way == 3'h3 ? valid_3_5 : _GEN_2586; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2926 = unuse_way == 3'h3 ? valid_3_6 : _GEN_2587; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2927 = unuse_way == 3'h3 ? valid_3_7 : _GEN_2588; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2928 = unuse_way == 3'h3 ? valid_3_8 : _GEN_2589; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2929 = unuse_way == 3'h3 ? valid_3_9 : _GEN_2590; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2930 = unuse_way == 3'h3 ? valid_3_10 : _GEN_2591; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2931 = unuse_way == 3'h3 ? valid_3_11 : _GEN_2592; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2932 = unuse_way == 3'h3 ? valid_3_12 : _GEN_2593; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2933 = unuse_way == 3'h3 ? valid_3_13 : _GEN_2594; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2934 = unuse_way == 3'h3 ? valid_3_14 : _GEN_2595; // @[d_cache.scala 180:40 32:26]
  wire  _GEN_2935 = unuse_way == 3'h3 ? valid_3_15 : _GEN_2596; // @[d_cache.scala 180:40 32:26]
  wire [511:0] _GEN_2936 = unuse_way == 3'h3 ? write_back_data : _GEN_2613; // @[d_cache.scala 180:40 44:34]
  wire [41:0] _GEN_2937 = unuse_way == 3'h3 ? {{10'd0}, write_back_addr} : _GEN_2614; // @[d_cache.scala 180:40 45:34]
  wire [511:0] _GEN_2938 = unuse_way == 3'h3 ? ram_0_0 : _GEN_2615; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2939 = unuse_way == 3'h3 ? ram_0_1 : _GEN_2616; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2940 = unuse_way == 3'h3 ? ram_0_2 : _GEN_2617; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2941 = unuse_way == 3'h3 ? ram_0_3 : _GEN_2618; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2942 = unuse_way == 3'h3 ? ram_0_4 : _GEN_2619; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2943 = unuse_way == 3'h3 ? ram_0_5 : _GEN_2620; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2944 = unuse_way == 3'h3 ? ram_0_6 : _GEN_2621; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2945 = unuse_way == 3'h3 ? ram_0_7 : _GEN_2622; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2946 = unuse_way == 3'h3 ? ram_0_8 : _GEN_2623; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2947 = unuse_way == 3'h3 ? ram_0_9 : _GEN_2624; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2948 = unuse_way == 3'h3 ? ram_0_10 : _GEN_2625; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2949 = unuse_way == 3'h3 ? ram_0_11 : _GEN_2626; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2950 = unuse_way == 3'h3 ? ram_0_12 : _GEN_2627; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2951 = unuse_way == 3'h3 ? ram_0_13 : _GEN_2628; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2952 = unuse_way == 3'h3 ? ram_0_14 : _GEN_2629; // @[d_cache.scala 180:40 19:24]
  wire [511:0] _GEN_2953 = unuse_way == 3'h3 ? ram_0_15 : _GEN_2630; // @[d_cache.scala 180:40 19:24]
  wire [31:0] _GEN_2954 = unuse_way == 3'h3 ? tag_0_0 : _GEN_2631; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2955 = unuse_way == 3'h3 ? tag_0_1 : _GEN_2632; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2956 = unuse_way == 3'h3 ? tag_0_2 : _GEN_2633; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2957 = unuse_way == 3'h3 ? tag_0_3 : _GEN_2634; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2958 = unuse_way == 3'h3 ? tag_0_4 : _GEN_2635; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2959 = unuse_way == 3'h3 ? tag_0_5 : _GEN_2636; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2960 = unuse_way == 3'h3 ? tag_0_6 : _GEN_2637; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2961 = unuse_way == 3'h3 ? tag_0_7 : _GEN_2638; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2962 = unuse_way == 3'h3 ? tag_0_8 : _GEN_2639; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2963 = unuse_way == 3'h3 ? tag_0_9 : _GEN_2640; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2964 = unuse_way == 3'h3 ? tag_0_10 : _GEN_2641; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2965 = unuse_way == 3'h3 ? tag_0_11 : _GEN_2642; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2966 = unuse_way == 3'h3 ? tag_0_12 : _GEN_2643; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2967 = unuse_way == 3'h3 ? tag_0_13 : _GEN_2644; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2968 = unuse_way == 3'h3 ? tag_0_14 : _GEN_2645; // @[d_cache.scala 180:40 24:24]
  wire [31:0] _GEN_2969 = unuse_way == 3'h3 ? tag_0_15 : _GEN_2646; // @[d_cache.scala 180:40 24:24]
  wire  _GEN_2970 = unuse_way == 3'h3 ? dirty_0_0 : _GEN_2647; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2971 = unuse_way == 3'h3 ? dirty_0_1 : _GEN_2648; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2972 = unuse_way == 3'h3 ? dirty_0_2 : _GEN_2649; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2973 = unuse_way == 3'h3 ? dirty_0_3 : _GEN_2650; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2974 = unuse_way == 3'h3 ? dirty_0_4 : _GEN_2651; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2975 = unuse_way == 3'h3 ? dirty_0_5 : _GEN_2652; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2976 = unuse_way == 3'h3 ? dirty_0_6 : _GEN_2653; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2977 = unuse_way == 3'h3 ? dirty_0_7 : _GEN_2654; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2978 = unuse_way == 3'h3 ? dirty_0_8 : _GEN_2655; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2979 = unuse_way == 3'h3 ? dirty_0_9 : _GEN_2656; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2980 = unuse_way == 3'h3 ? dirty_0_10 : _GEN_2657; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2981 = unuse_way == 3'h3 ? dirty_0_11 : _GEN_2658; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2982 = unuse_way == 3'h3 ? dirty_0_12 : _GEN_2659; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2983 = unuse_way == 3'h3 ? dirty_0_13 : _GEN_2660; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2984 = unuse_way == 3'h3 ? dirty_0_14 : _GEN_2661; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2985 = unuse_way == 3'h3 ? dirty_0_15 : _GEN_2662; // @[d_cache.scala 180:40 34:26]
  wire  _GEN_2986 = unuse_way == 3'h3 ? valid_0_0 : _GEN_2663; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2987 = unuse_way == 3'h3 ? valid_0_1 : _GEN_2664; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2988 = unuse_way == 3'h3 ? valid_0_2 : _GEN_2665; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2989 = unuse_way == 3'h3 ? valid_0_3 : _GEN_2666; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2990 = unuse_way == 3'h3 ? valid_0_4 : _GEN_2667; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2991 = unuse_way == 3'h3 ? valid_0_5 : _GEN_2668; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2992 = unuse_way == 3'h3 ? valid_0_6 : _GEN_2669; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2993 = unuse_way == 3'h3 ? valid_0_7 : _GEN_2670; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2994 = unuse_way == 3'h3 ? valid_0_8 : _GEN_2671; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2995 = unuse_way == 3'h3 ? valid_0_9 : _GEN_2672; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2996 = unuse_way == 3'h3 ? valid_0_10 : _GEN_2673; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2997 = unuse_way == 3'h3 ? valid_0_11 : _GEN_2674; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2998 = unuse_way == 3'h3 ? valid_0_12 : _GEN_2675; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_2999 = unuse_way == 3'h3 ? valid_0_13 : _GEN_2676; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_3000 = unuse_way == 3'h3 ? valid_0_14 : _GEN_2677; // @[d_cache.scala 180:40 29:26]
  wire  _GEN_3001 = unuse_way == 3'h3 ? valid_0_15 : _GEN_2678; // @[d_cache.scala 180:40 29:26]
  wire [511:0] _GEN_3002 = unuse_way == 3'h3 ? ram_1_0 : _GEN_2679; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3003 = unuse_way == 3'h3 ? ram_1_1 : _GEN_2680; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3004 = unuse_way == 3'h3 ? ram_1_2 : _GEN_2681; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3005 = unuse_way == 3'h3 ? ram_1_3 : _GEN_2682; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3006 = unuse_way == 3'h3 ? ram_1_4 : _GEN_2683; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3007 = unuse_way == 3'h3 ? ram_1_5 : _GEN_2684; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3008 = unuse_way == 3'h3 ? ram_1_6 : _GEN_2685; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3009 = unuse_way == 3'h3 ? ram_1_7 : _GEN_2686; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3010 = unuse_way == 3'h3 ? ram_1_8 : _GEN_2687; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3011 = unuse_way == 3'h3 ? ram_1_9 : _GEN_2688; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3012 = unuse_way == 3'h3 ? ram_1_10 : _GEN_2689; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3013 = unuse_way == 3'h3 ? ram_1_11 : _GEN_2690; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3014 = unuse_way == 3'h3 ? ram_1_12 : _GEN_2691; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3015 = unuse_way == 3'h3 ? ram_1_13 : _GEN_2692; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3016 = unuse_way == 3'h3 ? ram_1_14 : _GEN_2693; // @[d_cache.scala 180:40 20:24]
  wire [511:0] _GEN_3017 = unuse_way == 3'h3 ? ram_1_15 : _GEN_2694; // @[d_cache.scala 180:40 20:24]
  wire [31:0] _GEN_3018 = unuse_way == 3'h3 ? tag_1_0 : _GEN_2695; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3019 = unuse_way == 3'h3 ? tag_1_1 : _GEN_2696; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3020 = unuse_way == 3'h3 ? tag_1_2 : _GEN_2697; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3021 = unuse_way == 3'h3 ? tag_1_3 : _GEN_2698; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3022 = unuse_way == 3'h3 ? tag_1_4 : _GEN_2699; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3023 = unuse_way == 3'h3 ? tag_1_5 : _GEN_2700; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3024 = unuse_way == 3'h3 ? tag_1_6 : _GEN_2701; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3025 = unuse_way == 3'h3 ? tag_1_7 : _GEN_2702; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3026 = unuse_way == 3'h3 ? tag_1_8 : _GEN_2703; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3027 = unuse_way == 3'h3 ? tag_1_9 : _GEN_2704; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3028 = unuse_way == 3'h3 ? tag_1_10 : _GEN_2705; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3029 = unuse_way == 3'h3 ? tag_1_11 : _GEN_2706; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3030 = unuse_way == 3'h3 ? tag_1_12 : _GEN_2707; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3031 = unuse_way == 3'h3 ? tag_1_13 : _GEN_2708; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3032 = unuse_way == 3'h3 ? tag_1_14 : _GEN_2709; // @[d_cache.scala 180:40 25:24]
  wire [31:0] _GEN_3033 = unuse_way == 3'h3 ? tag_1_15 : _GEN_2710; // @[d_cache.scala 180:40 25:24]
  wire  _GEN_3034 = unuse_way == 3'h3 ? dirty_1_0 : _GEN_2711; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3035 = unuse_way == 3'h3 ? dirty_1_1 : _GEN_2712; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3036 = unuse_way == 3'h3 ? dirty_1_2 : _GEN_2713; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3037 = unuse_way == 3'h3 ? dirty_1_3 : _GEN_2714; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3038 = unuse_way == 3'h3 ? dirty_1_4 : _GEN_2715; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3039 = unuse_way == 3'h3 ? dirty_1_5 : _GEN_2716; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3040 = unuse_way == 3'h3 ? dirty_1_6 : _GEN_2717; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3041 = unuse_way == 3'h3 ? dirty_1_7 : _GEN_2718; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3042 = unuse_way == 3'h3 ? dirty_1_8 : _GEN_2719; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3043 = unuse_way == 3'h3 ? dirty_1_9 : _GEN_2720; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3044 = unuse_way == 3'h3 ? dirty_1_10 : _GEN_2721; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3045 = unuse_way == 3'h3 ? dirty_1_11 : _GEN_2722; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3046 = unuse_way == 3'h3 ? dirty_1_12 : _GEN_2723; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3047 = unuse_way == 3'h3 ? dirty_1_13 : _GEN_2724; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3048 = unuse_way == 3'h3 ? dirty_1_14 : _GEN_2725; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3049 = unuse_way == 3'h3 ? dirty_1_15 : _GEN_2726; // @[d_cache.scala 180:40 35:26]
  wire  _GEN_3050 = unuse_way == 3'h3 ? valid_1_0 : _GEN_2727; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3051 = unuse_way == 3'h3 ? valid_1_1 : _GEN_2728; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3052 = unuse_way == 3'h3 ? valid_1_2 : _GEN_2729; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3053 = unuse_way == 3'h3 ? valid_1_3 : _GEN_2730; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3054 = unuse_way == 3'h3 ? valid_1_4 : _GEN_2731; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3055 = unuse_way == 3'h3 ? valid_1_5 : _GEN_2732; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3056 = unuse_way == 3'h3 ? valid_1_6 : _GEN_2733; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3057 = unuse_way == 3'h3 ? valid_1_7 : _GEN_2734; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3058 = unuse_way == 3'h3 ? valid_1_8 : _GEN_2735; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3059 = unuse_way == 3'h3 ? valid_1_9 : _GEN_2736; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3060 = unuse_way == 3'h3 ? valid_1_10 : _GEN_2737; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3061 = unuse_way == 3'h3 ? valid_1_11 : _GEN_2738; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3062 = unuse_way == 3'h3 ? valid_1_12 : _GEN_2739; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3063 = unuse_way == 3'h3 ? valid_1_13 : _GEN_2740; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3064 = unuse_way == 3'h3 ? valid_1_14 : _GEN_2741; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3065 = unuse_way == 3'h3 ? valid_1_15 : _GEN_2742; // @[d_cache.scala 180:40 30:26]
  wire  _GEN_3066 = unuse_way == 3'h3 ? dirty_2_0 : _GEN_2775; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3067 = unuse_way == 3'h3 ? dirty_2_1 : _GEN_2776; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3068 = unuse_way == 3'h3 ? dirty_2_2 : _GEN_2777; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3069 = unuse_way == 3'h3 ? dirty_2_3 : _GEN_2778; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3070 = unuse_way == 3'h3 ? dirty_2_4 : _GEN_2779; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3071 = unuse_way == 3'h3 ? dirty_2_5 : _GEN_2780; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3072 = unuse_way == 3'h3 ? dirty_2_6 : _GEN_2781; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3073 = unuse_way == 3'h3 ? dirty_2_7 : _GEN_2782; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3074 = unuse_way == 3'h3 ? dirty_2_8 : _GEN_2783; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3075 = unuse_way == 3'h3 ? dirty_2_9 : _GEN_2784; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3076 = unuse_way == 3'h3 ? dirty_2_10 : _GEN_2785; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3077 = unuse_way == 3'h3 ? dirty_2_11 : _GEN_2786; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3078 = unuse_way == 3'h3 ? dirty_2_12 : _GEN_2787; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3079 = unuse_way == 3'h3 ? dirty_2_13 : _GEN_2788; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3080 = unuse_way == 3'h3 ? dirty_2_14 : _GEN_2789; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3081 = unuse_way == 3'h3 ? dirty_2_15 : _GEN_2790; // @[d_cache.scala 180:40 36:26]
  wire  _GEN_3082 = unuse_way == 3'h3 ? dirty_3_0 : _GEN_2807; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3083 = unuse_way == 3'h3 ? dirty_3_1 : _GEN_2808; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3084 = unuse_way == 3'h3 ? dirty_3_2 : _GEN_2809; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3085 = unuse_way == 3'h3 ? dirty_3_3 : _GEN_2810; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3086 = unuse_way == 3'h3 ? dirty_3_4 : _GEN_2811; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3087 = unuse_way == 3'h3 ? dirty_3_5 : _GEN_2812; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3088 = unuse_way == 3'h3 ? dirty_3_6 : _GEN_2813; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3089 = unuse_way == 3'h3 ? dirty_3_7 : _GEN_2814; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3090 = unuse_way == 3'h3 ? dirty_3_8 : _GEN_2815; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3091 = unuse_way == 3'h3 ? dirty_3_9 : _GEN_2816; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3092 = unuse_way == 3'h3 ? dirty_3_10 : _GEN_2817; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3093 = unuse_way == 3'h3 ? dirty_3_11 : _GEN_2818; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3094 = unuse_way == 3'h3 ? dirty_3_12 : _GEN_2819; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3095 = unuse_way == 3'h3 ? dirty_3_13 : _GEN_2820; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3096 = unuse_way == 3'h3 ? dirty_3_14 : _GEN_2821; // @[d_cache.scala 180:40 37:26]
  wire  _GEN_3097 = unuse_way == 3'h3 ? dirty_3_15 : _GEN_2822; // @[d_cache.scala 180:40 37:26]
  wire [3:0] _GEN_3098 = unuse_way == 3'h2 ? 4'h1 : _GEN_2823; // @[d_cache.scala 174:40 175:23]
  wire [511:0] _GEN_3099 = unuse_way == 3'h2 ? _GEN_751 : _GEN_3002; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3100 = unuse_way == 3'h2 ? _GEN_752 : _GEN_3003; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3101 = unuse_way == 3'h2 ? _GEN_753 : _GEN_3004; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3102 = unuse_way == 3'h2 ? _GEN_754 : _GEN_3005; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3103 = unuse_way == 3'h2 ? _GEN_755 : _GEN_3006; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3104 = unuse_way == 3'h2 ? _GEN_756 : _GEN_3007; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3105 = unuse_way == 3'h2 ? _GEN_757 : _GEN_3008; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3106 = unuse_way == 3'h2 ? _GEN_758 : _GEN_3009; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3107 = unuse_way == 3'h2 ? _GEN_759 : _GEN_3010; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3108 = unuse_way == 3'h2 ? _GEN_760 : _GEN_3011; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3109 = unuse_way == 3'h2 ? _GEN_761 : _GEN_3012; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3110 = unuse_way == 3'h2 ? _GEN_762 : _GEN_3013; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3111 = unuse_way == 3'h2 ? _GEN_763 : _GEN_3014; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3112 = unuse_way == 3'h2 ? _GEN_764 : _GEN_3015; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3113 = unuse_way == 3'h2 ? _GEN_765 : _GEN_3016; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3114 = unuse_way == 3'h2 ? _GEN_766 : _GEN_3017; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3115 = unuse_way == 3'h2 ? _GEN_767 : _GEN_3018; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3116 = unuse_way == 3'h2 ? _GEN_768 : _GEN_3019; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3117 = unuse_way == 3'h2 ? _GEN_769 : _GEN_3020; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3118 = unuse_way == 3'h2 ? _GEN_770 : _GEN_3021; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3119 = unuse_way == 3'h2 ? _GEN_771 : _GEN_3022; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3120 = unuse_way == 3'h2 ? _GEN_772 : _GEN_3023; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3121 = unuse_way == 3'h2 ? _GEN_773 : _GEN_3024; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3122 = unuse_way == 3'h2 ? _GEN_774 : _GEN_3025; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3123 = unuse_way == 3'h2 ? _GEN_775 : _GEN_3026; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3124 = unuse_way == 3'h2 ? _GEN_776 : _GEN_3027; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3125 = unuse_way == 3'h2 ? _GEN_777 : _GEN_3028; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3126 = unuse_way == 3'h2 ? _GEN_778 : _GEN_3029; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3127 = unuse_way == 3'h2 ? _GEN_779 : _GEN_3030; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3128 = unuse_way == 3'h2 ? _GEN_780 : _GEN_3031; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3129 = unuse_way == 3'h2 ? _GEN_781 : _GEN_3032; // @[d_cache.scala 174:40]
  wire [31:0] _GEN_3130 = unuse_way == 3'h2 ? _GEN_782 : _GEN_3033; // @[d_cache.scala 174:40]
  wire  _GEN_3131 = unuse_way == 3'h2 ? _GEN_783 : _GEN_3050; // @[d_cache.scala 174:40]
  wire  _GEN_3132 = unuse_way == 3'h2 ? _GEN_784 : _GEN_3051; // @[d_cache.scala 174:40]
  wire  _GEN_3133 = unuse_way == 3'h2 ? _GEN_785 : _GEN_3052; // @[d_cache.scala 174:40]
  wire  _GEN_3134 = unuse_way == 3'h2 ? _GEN_786 : _GEN_3053; // @[d_cache.scala 174:40]
  wire  _GEN_3135 = unuse_way == 3'h2 ? _GEN_787 : _GEN_3054; // @[d_cache.scala 174:40]
  wire  _GEN_3136 = unuse_way == 3'h2 ? _GEN_788 : _GEN_3055; // @[d_cache.scala 174:40]
  wire  _GEN_3137 = unuse_way == 3'h2 ? _GEN_789 : _GEN_3056; // @[d_cache.scala 174:40]
  wire  _GEN_3138 = unuse_way == 3'h2 ? _GEN_790 : _GEN_3057; // @[d_cache.scala 174:40]
  wire  _GEN_3139 = unuse_way == 3'h2 ? _GEN_791 : _GEN_3058; // @[d_cache.scala 174:40]
  wire  _GEN_3140 = unuse_way == 3'h2 ? _GEN_792 : _GEN_3059; // @[d_cache.scala 174:40]
  wire  _GEN_3141 = unuse_way == 3'h2 ? _GEN_793 : _GEN_3060; // @[d_cache.scala 174:40]
  wire  _GEN_3142 = unuse_way == 3'h2 ? _GEN_794 : _GEN_3061; // @[d_cache.scala 174:40]
  wire  _GEN_3143 = unuse_way == 3'h2 ? _GEN_795 : _GEN_3062; // @[d_cache.scala 174:40]
  wire  _GEN_3144 = unuse_way == 3'h2 ? _GEN_796 : _GEN_3063; // @[d_cache.scala 174:40]
  wire  _GEN_3145 = unuse_way == 3'h2 ? _GEN_797 : _GEN_3064; // @[d_cache.scala 174:40]
  wire  _GEN_3146 = unuse_way == 3'h2 ? _GEN_798 : _GEN_3065; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3147 = unuse_way == 3'h2 ? _GEN_799 : _GEN_2872; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3148 = unuse_way == 3'h2 ? _GEN_800 : _GEN_2873; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3149 = unuse_way == 3'h2 ? _GEN_801 : _GEN_2874; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3150 = unuse_way == 3'h2 ? _GEN_802 : _GEN_2875; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3151 = unuse_way == 3'h2 ? _GEN_803 : _GEN_2876; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3152 = unuse_way == 3'h2 ? _GEN_804 : _GEN_2877; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3153 = unuse_way == 3'h2 ? _GEN_805 : _GEN_2878; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3154 = unuse_way == 3'h2 ? _GEN_806 : _GEN_2879; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3155 = unuse_way == 3'h2 ? _GEN_807 : _GEN_2880; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3156 = unuse_way == 3'h2 ? _GEN_808 : _GEN_2881; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3157 = unuse_way == 3'h2 ? _GEN_809 : _GEN_2882; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3158 = unuse_way == 3'h2 ? _GEN_810 : _GEN_2883; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3159 = unuse_way == 3'h2 ? _GEN_811 : _GEN_2884; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3160 = unuse_way == 3'h2 ? _GEN_812 : _GEN_2885; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3161 = unuse_way == 3'h2 ? _GEN_813 : _GEN_2886; // @[d_cache.scala 174:40]
  wire [7:0] _GEN_3162 = unuse_way == 3'h2 ? _GEN_814 : _GEN_2887; // @[d_cache.scala 174:40]
  wire [511:0] _GEN_3163 = unuse_way == 3'h2 ? ram_2_0 : _GEN_2824; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3164 = unuse_way == 3'h2 ? ram_2_1 : _GEN_2825; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3165 = unuse_way == 3'h2 ? ram_2_2 : _GEN_2826; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3166 = unuse_way == 3'h2 ? ram_2_3 : _GEN_2827; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3167 = unuse_way == 3'h2 ? ram_2_4 : _GEN_2828; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3168 = unuse_way == 3'h2 ? ram_2_5 : _GEN_2829; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3169 = unuse_way == 3'h2 ? ram_2_6 : _GEN_2830; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3170 = unuse_way == 3'h2 ? ram_2_7 : _GEN_2831; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3171 = unuse_way == 3'h2 ? ram_2_8 : _GEN_2832; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3172 = unuse_way == 3'h2 ? ram_2_9 : _GEN_2833; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3173 = unuse_way == 3'h2 ? ram_2_10 : _GEN_2834; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3174 = unuse_way == 3'h2 ? ram_2_11 : _GEN_2835; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3175 = unuse_way == 3'h2 ? ram_2_12 : _GEN_2836; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3176 = unuse_way == 3'h2 ? ram_2_13 : _GEN_2837; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3177 = unuse_way == 3'h2 ? ram_2_14 : _GEN_2838; // @[d_cache.scala 174:40 21:24]
  wire [511:0] _GEN_3178 = unuse_way == 3'h2 ? ram_2_15 : _GEN_2839; // @[d_cache.scala 174:40 21:24]
  wire [31:0] _GEN_3179 = unuse_way == 3'h2 ? tag_2_0 : _GEN_2840; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3180 = unuse_way == 3'h2 ? tag_2_1 : _GEN_2841; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3181 = unuse_way == 3'h2 ? tag_2_2 : _GEN_2842; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3182 = unuse_way == 3'h2 ? tag_2_3 : _GEN_2843; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3183 = unuse_way == 3'h2 ? tag_2_4 : _GEN_2844; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3184 = unuse_way == 3'h2 ? tag_2_5 : _GEN_2845; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3185 = unuse_way == 3'h2 ? tag_2_6 : _GEN_2846; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3186 = unuse_way == 3'h2 ? tag_2_7 : _GEN_2847; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3187 = unuse_way == 3'h2 ? tag_2_8 : _GEN_2848; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3188 = unuse_way == 3'h2 ? tag_2_9 : _GEN_2849; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3189 = unuse_way == 3'h2 ? tag_2_10 : _GEN_2850; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3190 = unuse_way == 3'h2 ? tag_2_11 : _GEN_2851; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3191 = unuse_way == 3'h2 ? tag_2_12 : _GEN_2852; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3192 = unuse_way == 3'h2 ? tag_2_13 : _GEN_2853; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3193 = unuse_way == 3'h2 ? tag_2_14 : _GEN_2854; // @[d_cache.scala 174:40 26:24]
  wire [31:0] _GEN_3194 = unuse_way == 3'h2 ? tag_2_15 : _GEN_2855; // @[d_cache.scala 174:40 26:24]
  wire  _GEN_3195 = unuse_way == 3'h2 ? valid_2_0 : _GEN_2856; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3196 = unuse_way == 3'h2 ? valid_2_1 : _GEN_2857; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3197 = unuse_way == 3'h2 ? valid_2_2 : _GEN_2858; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3198 = unuse_way == 3'h2 ? valid_2_3 : _GEN_2859; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3199 = unuse_way == 3'h2 ? valid_2_4 : _GEN_2860; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3200 = unuse_way == 3'h2 ? valid_2_5 : _GEN_2861; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3201 = unuse_way == 3'h2 ? valid_2_6 : _GEN_2862; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3202 = unuse_way == 3'h2 ? valid_2_7 : _GEN_2863; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3203 = unuse_way == 3'h2 ? valid_2_8 : _GEN_2864; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3204 = unuse_way == 3'h2 ? valid_2_9 : _GEN_2865; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3205 = unuse_way == 3'h2 ? valid_2_10 : _GEN_2866; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3206 = unuse_way == 3'h2 ? valid_2_11 : _GEN_2867; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3207 = unuse_way == 3'h2 ? valid_2_12 : _GEN_2868; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3208 = unuse_way == 3'h2 ? valid_2_13 : _GEN_2869; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3209 = unuse_way == 3'h2 ? valid_2_14 : _GEN_2870; // @[d_cache.scala 174:40 31:26]
  wire  _GEN_3210 = unuse_way == 3'h2 ? valid_2_15 : _GEN_2871; // @[d_cache.scala 174:40 31:26]
  wire [511:0] _GEN_3211 = unuse_way == 3'h2 ? ram_3_0 : _GEN_2888; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3212 = unuse_way == 3'h2 ? ram_3_1 : _GEN_2889; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3213 = unuse_way == 3'h2 ? ram_3_2 : _GEN_2890; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3214 = unuse_way == 3'h2 ? ram_3_3 : _GEN_2891; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3215 = unuse_way == 3'h2 ? ram_3_4 : _GEN_2892; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3216 = unuse_way == 3'h2 ? ram_3_5 : _GEN_2893; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3217 = unuse_way == 3'h2 ? ram_3_6 : _GEN_2894; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3218 = unuse_way == 3'h2 ? ram_3_7 : _GEN_2895; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3219 = unuse_way == 3'h2 ? ram_3_8 : _GEN_2896; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3220 = unuse_way == 3'h2 ? ram_3_9 : _GEN_2897; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3221 = unuse_way == 3'h2 ? ram_3_10 : _GEN_2898; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3222 = unuse_way == 3'h2 ? ram_3_11 : _GEN_2899; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3223 = unuse_way == 3'h2 ? ram_3_12 : _GEN_2900; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3224 = unuse_way == 3'h2 ? ram_3_13 : _GEN_2901; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3225 = unuse_way == 3'h2 ? ram_3_14 : _GEN_2902; // @[d_cache.scala 174:40 22:24]
  wire [511:0] _GEN_3226 = unuse_way == 3'h2 ? ram_3_15 : _GEN_2903; // @[d_cache.scala 174:40 22:24]
  wire [31:0] _GEN_3227 = unuse_way == 3'h2 ? tag_3_0 : _GEN_2904; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3228 = unuse_way == 3'h2 ? tag_3_1 : _GEN_2905; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3229 = unuse_way == 3'h2 ? tag_3_2 : _GEN_2906; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3230 = unuse_way == 3'h2 ? tag_3_3 : _GEN_2907; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3231 = unuse_way == 3'h2 ? tag_3_4 : _GEN_2908; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3232 = unuse_way == 3'h2 ? tag_3_5 : _GEN_2909; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3233 = unuse_way == 3'h2 ? tag_3_6 : _GEN_2910; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3234 = unuse_way == 3'h2 ? tag_3_7 : _GEN_2911; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3235 = unuse_way == 3'h2 ? tag_3_8 : _GEN_2912; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3236 = unuse_way == 3'h2 ? tag_3_9 : _GEN_2913; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3237 = unuse_way == 3'h2 ? tag_3_10 : _GEN_2914; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3238 = unuse_way == 3'h2 ? tag_3_11 : _GEN_2915; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3239 = unuse_way == 3'h2 ? tag_3_12 : _GEN_2916; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3240 = unuse_way == 3'h2 ? tag_3_13 : _GEN_2917; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3241 = unuse_way == 3'h2 ? tag_3_14 : _GEN_2918; // @[d_cache.scala 174:40 27:24]
  wire [31:0] _GEN_3242 = unuse_way == 3'h2 ? tag_3_15 : _GEN_2919; // @[d_cache.scala 174:40 27:24]
  wire  _GEN_3243 = unuse_way == 3'h2 ? valid_3_0 : _GEN_2920; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3244 = unuse_way == 3'h2 ? valid_3_1 : _GEN_2921; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3245 = unuse_way == 3'h2 ? valid_3_2 : _GEN_2922; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3246 = unuse_way == 3'h2 ? valid_3_3 : _GEN_2923; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3247 = unuse_way == 3'h2 ? valid_3_4 : _GEN_2924; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3248 = unuse_way == 3'h2 ? valid_3_5 : _GEN_2925; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3249 = unuse_way == 3'h2 ? valid_3_6 : _GEN_2926; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3250 = unuse_way == 3'h2 ? valid_3_7 : _GEN_2927; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3251 = unuse_way == 3'h2 ? valid_3_8 : _GEN_2928; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3252 = unuse_way == 3'h2 ? valid_3_9 : _GEN_2929; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3253 = unuse_way == 3'h2 ? valid_3_10 : _GEN_2930; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3254 = unuse_way == 3'h2 ? valid_3_11 : _GEN_2931; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3255 = unuse_way == 3'h2 ? valid_3_12 : _GEN_2932; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3256 = unuse_way == 3'h2 ? valid_3_13 : _GEN_2933; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3257 = unuse_way == 3'h2 ? valid_3_14 : _GEN_2934; // @[d_cache.scala 174:40 32:26]
  wire  _GEN_3258 = unuse_way == 3'h2 ? valid_3_15 : _GEN_2935; // @[d_cache.scala 174:40 32:26]
  wire [511:0] _GEN_3259 = unuse_way == 3'h2 ? write_back_data : _GEN_2936; // @[d_cache.scala 174:40 44:34]
  wire [41:0] _GEN_3260 = unuse_way == 3'h2 ? {{10'd0}, write_back_addr} : _GEN_2937; // @[d_cache.scala 174:40 45:34]
  wire [511:0] _GEN_3261 = unuse_way == 3'h2 ? ram_0_0 : _GEN_2938; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3262 = unuse_way == 3'h2 ? ram_0_1 : _GEN_2939; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3263 = unuse_way == 3'h2 ? ram_0_2 : _GEN_2940; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3264 = unuse_way == 3'h2 ? ram_0_3 : _GEN_2941; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3265 = unuse_way == 3'h2 ? ram_0_4 : _GEN_2942; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3266 = unuse_way == 3'h2 ? ram_0_5 : _GEN_2943; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3267 = unuse_way == 3'h2 ? ram_0_6 : _GEN_2944; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3268 = unuse_way == 3'h2 ? ram_0_7 : _GEN_2945; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3269 = unuse_way == 3'h2 ? ram_0_8 : _GEN_2946; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3270 = unuse_way == 3'h2 ? ram_0_9 : _GEN_2947; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3271 = unuse_way == 3'h2 ? ram_0_10 : _GEN_2948; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3272 = unuse_way == 3'h2 ? ram_0_11 : _GEN_2949; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3273 = unuse_way == 3'h2 ? ram_0_12 : _GEN_2950; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3274 = unuse_way == 3'h2 ? ram_0_13 : _GEN_2951; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3275 = unuse_way == 3'h2 ? ram_0_14 : _GEN_2952; // @[d_cache.scala 174:40 19:24]
  wire [511:0] _GEN_3276 = unuse_way == 3'h2 ? ram_0_15 : _GEN_2953; // @[d_cache.scala 174:40 19:24]
  wire [31:0] _GEN_3277 = unuse_way == 3'h2 ? tag_0_0 : _GEN_2954; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3278 = unuse_way == 3'h2 ? tag_0_1 : _GEN_2955; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3279 = unuse_way == 3'h2 ? tag_0_2 : _GEN_2956; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3280 = unuse_way == 3'h2 ? tag_0_3 : _GEN_2957; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3281 = unuse_way == 3'h2 ? tag_0_4 : _GEN_2958; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3282 = unuse_way == 3'h2 ? tag_0_5 : _GEN_2959; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3283 = unuse_way == 3'h2 ? tag_0_6 : _GEN_2960; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3284 = unuse_way == 3'h2 ? tag_0_7 : _GEN_2961; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3285 = unuse_way == 3'h2 ? tag_0_8 : _GEN_2962; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3286 = unuse_way == 3'h2 ? tag_0_9 : _GEN_2963; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3287 = unuse_way == 3'h2 ? tag_0_10 : _GEN_2964; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3288 = unuse_way == 3'h2 ? tag_0_11 : _GEN_2965; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3289 = unuse_way == 3'h2 ? tag_0_12 : _GEN_2966; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3290 = unuse_way == 3'h2 ? tag_0_13 : _GEN_2967; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3291 = unuse_way == 3'h2 ? tag_0_14 : _GEN_2968; // @[d_cache.scala 174:40 24:24]
  wire [31:0] _GEN_3292 = unuse_way == 3'h2 ? tag_0_15 : _GEN_2969; // @[d_cache.scala 174:40 24:24]
  wire  _GEN_3293 = unuse_way == 3'h2 ? dirty_0_0 : _GEN_2970; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3294 = unuse_way == 3'h2 ? dirty_0_1 : _GEN_2971; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3295 = unuse_way == 3'h2 ? dirty_0_2 : _GEN_2972; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3296 = unuse_way == 3'h2 ? dirty_0_3 : _GEN_2973; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3297 = unuse_way == 3'h2 ? dirty_0_4 : _GEN_2974; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3298 = unuse_way == 3'h2 ? dirty_0_5 : _GEN_2975; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3299 = unuse_way == 3'h2 ? dirty_0_6 : _GEN_2976; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3300 = unuse_way == 3'h2 ? dirty_0_7 : _GEN_2977; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3301 = unuse_way == 3'h2 ? dirty_0_8 : _GEN_2978; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3302 = unuse_way == 3'h2 ? dirty_0_9 : _GEN_2979; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3303 = unuse_way == 3'h2 ? dirty_0_10 : _GEN_2980; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3304 = unuse_way == 3'h2 ? dirty_0_11 : _GEN_2981; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3305 = unuse_way == 3'h2 ? dirty_0_12 : _GEN_2982; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3306 = unuse_way == 3'h2 ? dirty_0_13 : _GEN_2983; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3307 = unuse_way == 3'h2 ? dirty_0_14 : _GEN_2984; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3308 = unuse_way == 3'h2 ? dirty_0_15 : _GEN_2985; // @[d_cache.scala 174:40 34:26]
  wire  _GEN_3309 = unuse_way == 3'h2 ? valid_0_0 : _GEN_2986; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3310 = unuse_way == 3'h2 ? valid_0_1 : _GEN_2987; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3311 = unuse_way == 3'h2 ? valid_0_2 : _GEN_2988; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3312 = unuse_way == 3'h2 ? valid_0_3 : _GEN_2989; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3313 = unuse_way == 3'h2 ? valid_0_4 : _GEN_2990; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3314 = unuse_way == 3'h2 ? valid_0_5 : _GEN_2991; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3315 = unuse_way == 3'h2 ? valid_0_6 : _GEN_2992; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3316 = unuse_way == 3'h2 ? valid_0_7 : _GEN_2993; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3317 = unuse_way == 3'h2 ? valid_0_8 : _GEN_2994; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3318 = unuse_way == 3'h2 ? valid_0_9 : _GEN_2995; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3319 = unuse_way == 3'h2 ? valid_0_10 : _GEN_2996; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3320 = unuse_way == 3'h2 ? valid_0_11 : _GEN_2997; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3321 = unuse_way == 3'h2 ? valid_0_12 : _GEN_2998; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3322 = unuse_way == 3'h2 ? valid_0_13 : _GEN_2999; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3323 = unuse_way == 3'h2 ? valid_0_14 : _GEN_3000; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3324 = unuse_way == 3'h2 ? valid_0_15 : _GEN_3001; // @[d_cache.scala 174:40 29:26]
  wire  _GEN_3325 = unuse_way == 3'h2 ? dirty_1_0 : _GEN_3034; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3326 = unuse_way == 3'h2 ? dirty_1_1 : _GEN_3035; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3327 = unuse_way == 3'h2 ? dirty_1_2 : _GEN_3036; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3328 = unuse_way == 3'h2 ? dirty_1_3 : _GEN_3037; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3329 = unuse_way == 3'h2 ? dirty_1_4 : _GEN_3038; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3330 = unuse_way == 3'h2 ? dirty_1_5 : _GEN_3039; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3331 = unuse_way == 3'h2 ? dirty_1_6 : _GEN_3040; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3332 = unuse_way == 3'h2 ? dirty_1_7 : _GEN_3041; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3333 = unuse_way == 3'h2 ? dirty_1_8 : _GEN_3042; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3334 = unuse_way == 3'h2 ? dirty_1_9 : _GEN_3043; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3335 = unuse_way == 3'h2 ? dirty_1_10 : _GEN_3044; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3336 = unuse_way == 3'h2 ? dirty_1_11 : _GEN_3045; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3337 = unuse_way == 3'h2 ? dirty_1_12 : _GEN_3046; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3338 = unuse_way == 3'h2 ? dirty_1_13 : _GEN_3047; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3339 = unuse_way == 3'h2 ? dirty_1_14 : _GEN_3048; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3340 = unuse_way == 3'h2 ? dirty_1_15 : _GEN_3049; // @[d_cache.scala 174:40 35:26]
  wire  _GEN_3341 = unuse_way == 3'h2 ? dirty_2_0 : _GEN_3066; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3342 = unuse_way == 3'h2 ? dirty_2_1 : _GEN_3067; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3343 = unuse_way == 3'h2 ? dirty_2_2 : _GEN_3068; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3344 = unuse_way == 3'h2 ? dirty_2_3 : _GEN_3069; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3345 = unuse_way == 3'h2 ? dirty_2_4 : _GEN_3070; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3346 = unuse_way == 3'h2 ? dirty_2_5 : _GEN_3071; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3347 = unuse_way == 3'h2 ? dirty_2_6 : _GEN_3072; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3348 = unuse_way == 3'h2 ? dirty_2_7 : _GEN_3073; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3349 = unuse_way == 3'h2 ? dirty_2_8 : _GEN_3074; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3350 = unuse_way == 3'h2 ? dirty_2_9 : _GEN_3075; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3351 = unuse_way == 3'h2 ? dirty_2_10 : _GEN_3076; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3352 = unuse_way == 3'h2 ? dirty_2_11 : _GEN_3077; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3353 = unuse_way == 3'h2 ? dirty_2_12 : _GEN_3078; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3354 = unuse_way == 3'h2 ? dirty_2_13 : _GEN_3079; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3355 = unuse_way == 3'h2 ? dirty_2_14 : _GEN_3080; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3356 = unuse_way == 3'h2 ? dirty_2_15 : _GEN_3081; // @[d_cache.scala 174:40 36:26]
  wire  _GEN_3357 = unuse_way == 3'h2 ? dirty_3_0 : _GEN_3082; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3358 = unuse_way == 3'h2 ? dirty_3_1 : _GEN_3083; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3359 = unuse_way == 3'h2 ? dirty_3_2 : _GEN_3084; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3360 = unuse_way == 3'h2 ? dirty_3_3 : _GEN_3085; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3361 = unuse_way == 3'h2 ? dirty_3_4 : _GEN_3086; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3362 = unuse_way == 3'h2 ? dirty_3_5 : _GEN_3087; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3363 = unuse_way == 3'h2 ? dirty_3_6 : _GEN_3088; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3364 = unuse_way == 3'h2 ? dirty_3_7 : _GEN_3089; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3365 = unuse_way == 3'h2 ? dirty_3_8 : _GEN_3090; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3366 = unuse_way == 3'h2 ? dirty_3_9 : _GEN_3091; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3367 = unuse_way == 3'h2 ? dirty_3_10 : _GEN_3092; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3368 = unuse_way == 3'h2 ? dirty_3_11 : _GEN_3093; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3369 = unuse_way == 3'h2 ? dirty_3_12 : _GEN_3094; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3370 = unuse_way == 3'h2 ? dirty_3_13 : _GEN_3095; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3371 = unuse_way == 3'h2 ? dirty_3_14 : _GEN_3096; // @[d_cache.scala 174:40 37:26]
  wire  _GEN_3372 = unuse_way == 3'h2 ? dirty_3_15 : _GEN_3097; // @[d_cache.scala 174:40 37:26]
  wire [3:0] _GEN_3373 = unuse_way == 3'h1 ? 4'h1 : _GEN_3098; // @[d_cache.scala 168:34 169:23]
  wire [511:0] _GEN_3374 = unuse_way == 3'h1 ? _GEN_671 : _GEN_3261; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3375 = unuse_way == 3'h1 ? _GEN_672 : _GEN_3262; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3376 = unuse_way == 3'h1 ? _GEN_673 : _GEN_3263; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3377 = unuse_way == 3'h1 ? _GEN_674 : _GEN_3264; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3378 = unuse_way == 3'h1 ? _GEN_675 : _GEN_3265; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3379 = unuse_way == 3'h1 ? _GEN_676 : _GEN_3266; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3380 = unuse_way == 3'h1 ? _GEN_677 : _GEN_3267; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3381 = unuse_way == 3'h1 ? _GEN_678 : _GEN_3268; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3382 = unuse_way == 3'h1 ? _GEN_679 : _GEN_3269; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3383 = unuse_way == 3'h1 ? _GEN_680 : _GEN_3270; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3384 = unuse_way == 3'h1 ? _GEN_681 : _GEN_3271; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3385 = unuse_way == 3'h1 ? _GEN_682 : _GEN_3272; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3386 = unuse_way == 3'h1 ? _GEN_683 : _GEN_3273; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3387 = unuse_way == 3'h1 ? _GEN_684 : _GEN_3274; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3388 = unuse_way == 3'h1 ? _GEN_685 : _GEN_3275; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3389 = unuse_way == 3'h1 ? _GEN_686 : _GEN_3276; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3390 = unuse_way == 3'h1 ? _GEN_687 : _GEN_3277; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3391 = unuse_way == 3'h1 ? _GEN_688 : _GEN_3278; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3392 = unuse_way == 3'h1 ? _GEN_689 : _GEN_3279; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3393 = unuse_way == 3'h1 ? _GEN_690 : _GEN_3280; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3394 = unuse_way == 3'h1 ? _GEN_691 : _GEN_3281; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3395 = unuse_way == 3'h1 ? _GEN_692 : _GEN_3282; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3396 = unuse_way == 3'h1 ? _GEN_693 : _GEN_3283; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3397 = unuse_way == 3'h1 ? _GEN_694 : _GEN_3284; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3398 = unuse_way == 3'h1 ? _GEN_695 : _GEN_3285; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3399 = unuse_way == 3'h1 ? _GEN_696 : _GEN_3286; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3400 = unuse_way == 3'h1 ? _GEN_697 : _GEN_3287; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3401 = unuse_way == 3'h1 ? _GEN_698 : _GEN_3288; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3402 = unuse_way == 3'h1 ? _GEN_699 : _GEN_3289; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3403 = unuse_way == 3'h1 ? _GEN_700 : _GEN_3290; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3404 = unuse_way == 3'h1 ? _GEN_701 : _GEN_3291; // @[d_cache.scala 168:34]
  wire [31:0] _GEN_3405 = unuse_way == 3'h1 ? _GEN_702 : _GEN_3292; // @[d_cache.scala 168:34]
  wire  _GEN_3406 = unuse_way == 3'h1 ? _GEN_703 : _GEN_3309; // @[d_cache.scala 168:34]
  wire  _GEN_3407 = unuse_way == 3'h1 ? _GEN_704 : _GEN_3310; // @[d_cache.scala 168:34]
  wire  _GEN_3408 = unuse_way == 3'h1 ? _GEN_705 : _GEN_3311; // @[d_cache.scala 168:34]
  wire  _GEN_3409 = unuse_way == 3'h1 ? _GEN_706 : _GEN_3312; // @[d_cache.scala 168:34]
  wire  _GEN_3410 = unuse_way == 3'h1 ? _GEN_707 : _GEN_3313; // @[d_cache.scala 168:34]
  wire  _GEN_3411 = unuse_way == 3'h1 ? _GEN_708 : _GEN_3314; // @[d_cache.scala 168:34]
  wire  _GEN_3412 = unuse_way == 3'h1 ? _GEN_709 : _GEN_3315; // @[d_cache.scala 168:34]
  wire  _GEN_3413 = unuse_way == 3'h1 ? _GEN_710 : _GEN_3316; // @[d_cache.scala 168:34]
  wire  _GEN_3414 = unuse_way == 3'h1 ? _GEN_711 : _GEN_3317; // @[d_cache.scala 168:34]
  wire  _GEN_3415 = unuse_way == 3'h1 ? _GEN_712 : _GEN_3318; // @[d_cache.scala 168:34]
  wire  _GEN_3416 = unuse_way == 3'h1 ? _GEN_713 : _GEN_3319; // @[d_cache.scala 168:34]
  wire  _GEN_3417 = unuse_way == 3'h1 ? _GEN_714 : _GEN_3320; // @[d_cache.scala 168:34]
  wire  _GEN_3418 = unuse_way == 3'h1 ? _GEN_715 : _GEN_3321; // @[d_cache.scala 168:34]
  wire  _GEN_3419 = unuse_way == 3'h1 ? _GEN_716 : _GEN_3322; // @[d_cache.scala 168:34]
  wire  _GEN_3420 = unuse_way == 3'h1 ? _GEN_717 : _GEN_3323; // @[d_cache.scala 168:34]
  wire  _GEN_3421 = unuse_way == 3'h1 ? _GEN_718 : _GEN_3324; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3422 = unuse_way == 3'h1 ? _GEN_735 : _GEN_3147; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3423 = unuse_way == 3'h1 ? _GEN_736 : _GEN_3148; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3424 = unuse_way == 3'h1 ? _GEN_737 : _GEN_3149; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3425 = unuse_way == 3'h1 ? _GEN_738 : _GEN_3150; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3426 = unuse_way == 3'h1 ? _GEN_739 : _GEN_3151; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3427 = unuse_way == 3'h1 ? _GEN_740 : _GEN_3152; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3428 = unuse_way == 3'h1 ? _GEN_741 : _GEN_3153; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3429 = unuse_way == 3'h1 ? _GEN_742 : _GEN_3154; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3430 = unuse_way == 3'h1 ? _GEN_743 : _GEN_3155; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3431 = unuse_way == 3'h1 ? _GEN_744 : _GEN_3156; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3432 = unuse_way == 3'h1 ? _GEN_745 : _GEN_3157; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3433 = unuse_way == 3'h1 ? _GEN_746 : _GEN_3158; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3434 = unuse_way == 3'h1 ? _GEN_747 : _GEN_3159; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3435 = unuse_way == 3'h1 ? _GEN_748 : _GEN_3160; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3436 = unuse_way == 3'h1 ? _GEN_749 : _GEN_3161; // @[d_cache.scala 168:34]
  wire [7:0] _GEN_3437 = unuse_way == 3'h1 ? _GEN_750 : _GEN_3162; // @[d_cache.scala 168:34]
  wire [511:0] _GEN_3438 = unuse_way == 3'h1 ? ram_1_0 : _GEN_3099; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3439 = unuse_way == 3'h1 ? ram_1_1 : _GEN_3100; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3440 = unuse_way == 3'h1 ? ram_1_2 : _GEN_3101; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3441 = unuse_way == 3'h1 ? ram_1_3 : _GEN_3102; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3442 = unuse_way == 3'h1 ? ram_1_4 : _GEN_3103; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3443 = unuse_way == 3'h1 ? ram_1_5 : _GEN_3104; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3444 = unuse_way == 3'h1 ? ram_1_6 : _GEN_3105; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3445 = unuse_way == 3'h1 ? ram_1_7 : _GEN_3106; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3446 = unuse_way == 3'h1 ? ram_1_8 : _GEN_3107; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3447 = unuse_way == 3'h1 ? ram_1_9 : _GEN_3108; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3448 = unuse_way == 3'h1 ? ram_1_10 : _GEN_3109; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3449 = unuse_way == 3'h1 ? ram_1_11 : _GEN_3110; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3450 = unuse_way == 3'h1 ? ram_1_12 : _GEN_3111; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3451 = unuse_way == 3'h1 ? ram_1_13 : _GEN_3112; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3452 = unuse_way == 3'h1 ? ram_1_14 : _GEN_3113; // @[d_cache.scala 168:34 20:24]
  wire [511:0] _GEN_3453 = unuse_way == 3'h1 ? ram_1_15 : _GEN_3114; // @[d_cache.scala 168:34 20:24]
  wire [31:0] _GEN_3454 = unuse_way == 3'h1 ? tag_1_0 : _GEN_3115; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3455 = unuse_way == 3'h1 ? tag_1_1 : _GEN_3116; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3456 = unuse_way == 3'h1 ? tag_1_2 : _GEN_3117; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3457 = unuse_way == 3'h1 ? tag_1_3 : _GEN_3118; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3458 = unuse_way == 3'h1 ? tag_1_4 : _GEN_3119; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3459 = unuse_way == 3'h1 ? tag_1_5 : _GEN_3120; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3460 = unuse_way == 3'h1 ? tag_1_6 : _GEN_3121; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3461 = unuse_way == 3'h1 ? tag_1_7 : _GEN_3122; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3462 = unuse_way == 3'h1 ? tag_1_8 : _GEN_3123; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3463 = unuse_way == 3'h1 ? tag_1_9 : _GEN_3124; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3464 = unuse_way == 3'h1 ? tag_1_10 : _GEN_3125; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3465 = unuse_way == 3'h1 ? tag_1_11 : _GEN_3126; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3466 = unuse_way == 3'h1 ? tag_1_12 : _GEN_3127; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3467 = unuse_way == 3'h1 ? tag_1_13 : _GEN_3128; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3468 = unuse_way == 3'h1 ? tag_1_14 : _GEN_3129; // @[d_cache.scala 168:34 25:24]
  wire [31:0] _GEN_3469 = unuse_way == 3'h1 ? tag_1_15 : _GEN_3130; // @[d_cache.scala 168:34 25:24]
  wire  _GEN_3470 = unuse_way == 3'h1 ? valid_1_0 : _GEN_3131; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3471 = unuse_way == 3'h1 ? valid_1_1 : _GEN_3132; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3472 = unuse_way == 3'h1 ? valid_1_2 : _GEN_3133; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3473 = unuse_way == 3'h1 ? valid_1_3 : _GEN_3134; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3474 = unuse_way == 3'h1 ? valid_1_4 : _GEN_3135; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3475 = unuse_way == 3'h1 ? valid_1_5 : _GEN_3136; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3476 = unuse_way == 3'h1 ? valid_1_6 : _GEN_3137; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3477 = unuse_way == 3'h1 ? valid_1_7 : _GEN_3138; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3478 = unuse_way == 3'h1 ? valid_1_8 : _GEN_3139; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3479 = unuse_way == 3'h1 ? valid_1_9 : _GEN_3140; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3480 = unuse_way == 3'h1 ? valid_1_10 : _GEN_3141; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3481 = unuse_way == 3'h1 ? valid_1_11 : _GEN_3142; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3482 = unuse_way == 3'h1 ? valid_1_12 : _GEN_3143; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3483 = unuse_way == 3'h1 ? valid_1_13 : _GEN_3144; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3484 = unuse_way == 3'h1 ? valid_1_14 : _GEN_3145; // @[d_cache.scala 168:34 30:26]
  wire  _GEN_3485 = unuse_way == 3'h1 ? valid_1_15 : _GEN_3146; // @[d_cache.scala 168:34 30:26]
  wire [511:0] _GEN_3486 = unuse_way == 3'h1 ? ram_2_0 : _GEN_3163; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3487 = unuse_way == 3'h1 ? ram_2_1 : _GEN_3164; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3488 = unuse_way == 3'h1 ? ram_2_2 : _GEN_3165; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3489 = unuse_way == 3'h1 ? ram_2_3 : _GEN_3166; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3490 = unuse_way == 3'h1 ? ram_2_4 : _GEN_3167; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3491 = unuse_way == 3'h1 ? ram_2_5 : _GEN_3168; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3492 = unuse_way == 3'h1 ? ram_2_6 : _GEN_3169; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3493 = unuse_way == 3'h1 ? ram_2_7 : _GEN_3170; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3494 = unuse_way == 3'h1 ? ram_2_8 : _GEN_3171; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3495 = unuse_way == 3'h1 ? ram_2_9 : _GEN_3172; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3496 = unuse_way == 3'h1 ? ram_2_10 : _GEN_3173; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3497 = unuse_way == 3'h1 ? ram_2_11 : _GEN_3174; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3498 = unuse_way == 3'h1 ? ram_2_12 : _GEN_3175; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3499 = unuse_way == 3'h1 ? ram_2_13 : _GEN_3176; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3500 = unuse_way == 3'h1 ? ram_2_14 : _GEN_3177; // @[d_cache.scala 168:34 21:24]
  wire [511:0] _GEN_3501 = unuse_way == 3'h1 ? ram_2_15 : _GEN_3178; // @[d_cache.scala 168:34 21:24]
  wire [31:0] _GEN_3502 = unuse_way == 3'h1 ? tag_2_0 : _GEN_3179; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3503 = unuse_way == 3'h1 ? tag_2_1 : _GEN_3180; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3504 = unuse_way == 3'h1 ? tag_2_2 : _GEN_3181; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3505 = unuse_way == 3'h1 ? tag_2_3 : _GEN_3182; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3506 = unuse_way == 3'h1 ? tag_2_4 : _GEN_3183; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3507 = unuse_way == 3'h1 ? tag_2_5 : _GEN_3184; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3508 = unuse_way == 3'h1 ? tag_2_6 : _GEN_3185; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3509 = unuse_way == 3'h1 ? tag_2_7 : _GEN_3186; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3510 = unuse_way == 3'h1 ? tag_2_8 : _GEN_3187; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3511 = unuse_way == 3'h1 ? tag_2_9 : _GEN_3188; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3512 = unuse_way == 3'h1 ? tag_2_10 : _GEN_3189; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3513 = unuse_way == 3'h1 ? tag_2_11 : _GEN_3190; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3514 = unuse_way == 3'h1 ? tag_2_12 : _GEN_3191; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3515 = unuse_way == 3'h1 ? tag_2_13 : _GEN_3192; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3516 = unuse_way == 3'h1 ? tag_2_14 : _GEN_3193; // @[d_cache.scala 168:34 26:24]
  wire [31:0] _GEN_3517 = unuse_way == 3'h1 ? tag_2_15 : _GEN_3194; // @[d_cache.scala 168:34 26:24]
  wire  _GEN_3518 = unuse_way == 3'h1 ? valid_2_0 : _GEN_3195; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3519 = unuse_way == 3'h1 ? valid_2_1 : _GEN_3196; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3520 = unuse_way == 3'h1 ? valid_2_2 : _GEN_3197; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3521 = unuse_way == 3'h1 ? valid_2_3 : _GEN_3198; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3522 = unuse_way == 3'h1 ? valid_2_4 : _GEN_3199; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3523 = unuse_way == 3'h1 ? valid_2_5 : _GEN_3200; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3524 = unuse_way == 3'h1 ? valid_2_6 : _GEN_3201; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3525 = unuse_way == 3'h1 ? valid_2_7 : _GEN_3202; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3526 = unuse_way == 3'h1 ? valid_2_8 : _GEN_3203; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3527 = unuse_way == 3'h1 ? valid_2_9 : _GEN_3204; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3528 = unuse_way == 3'h1 ? valid_2_10 : _GEN_3205; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3529 = unuse_way == 3'h1 ? valid_2_11 : _GEN_3206; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3530 = unuse_way == 3'h1 ? valid_2_12 : _GEN_3207; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3531 = unuse_way == 3'h1 ? valid_2_13 : _GEN_3208; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3532 = unuse_way == 3'h1 ? valid_2_14 : _GEN_3209; // @[d_cache.scala 168:34 31:26]
  wire  _GEN_3533 = unuse_way == 3'h1 ? valid_2_15 : _GEN_3210; // @[d_cache.scala 168:34 31:26]
  wire [511:0] _GEN_3534 = unuse_way == 3'h1 ? ram_3_0 : _GEN_3211; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3535 = unuse_way == 3'h1 ? ram_3_1 : _GEN_3212; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3536 = unuse_way == 3'h1 ? ram_3_2 : _GEN_3213; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3537 = unuse_way == 3'h1 ? ram_3_3 : _GEN_3214; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3538 = unuse_way == 3'h1 ? ram_3_4 : _GEN_3215; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3539 = unuse_way == 3'h1 ? ram_3_5 : _GEN_3216; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3540 = unuse_way == 3'h1 ? ram_3_6 : _GEN_3217; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3541 = unuse_way == 3'h1 ? ram_3_7 : _GEN_3218; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3542 = unuse_way == 3'h1 ? ram_3_8 : _GEN_3219; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3543 = unuse_way == 3'h1 ? ram_3_9 : _GEN_3220; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3544 = unuse_way == 3'h1 ? ram_3_10 : _GEN_3221; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3545 = unuse_way == 3'h1 ? ram_3_11 : _GEN_3222; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3546 = unuse_way == 3'h1 ? ram_3_12 : _GEN_3223; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3547 = unuse_way == 3'h1 ? ram_3_13 : _GEN_3224; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3548 = unuse_way == 3'h1 ? ram_3_14 : _GEN_3225; // @[d_cache.scala 168:34 22:24]
  wire [511:0] _GEN_3549 = unuse_way == 3'h1 ? ram_3_15 : _GEN_3226; // @[d_cache.scala 168:34 22:24]
  wire [31:0] _GEN_3550 = unuse_way == 3'h1 ? tag_3_0 : _GEN_3227; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3551 = unuse_way == 3'h1 ? tag_3_1 : _GEN_3228; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3552 = unuse_way == 3'h1 ? tag_3_2 : _GEN_3229; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3553 = unuse_way == 3'h1 ? tag_3_3 : _GEN_3230; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3554 = unuse_way == 3'h1 ? tag_3_4 : _GEN_3231; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3555 = unuse_way == 3'h1 ? tag_3_5 : _GEN_3232; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3556 = unuse_way == 3'h1 ? tag_3_6 : _GEN_3233; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3557 = unuse_way == 3'h1 ? tag_3_7 : _GEN_3234; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3558 = unuse_way == 3'h1 ? tag_3_8 : _GEN_3235; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3559 = unuse_way == 3'h1 ? tag_3_9 : _GEN_3236; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3560 = unuse_way == 3'h1 ? tag_3_10 : _GEN_3237; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3561 = unuse_way == 3'h1 ? tag_3_11 : _GEN_3238; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3562 = unuse_way == 3'h1 ? tag_3_12 : _GEN_3239; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3563 = unuse_way == 3'h1 ? tag_3_13 : _GEN_3240; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3564 = unuse_way == 3'h1 ? tag_3_14 : _GEN_3241; // @[d_cache.scala 168:34 27:24]
  wire [31:0] _GEN_3565 = unuse_way == 3'h1 ? tag_3_15 : _GEN_3242; // @[d_cache.scala 168:34 27:24]
  wire  _GEN_3566 = unuse_way == 3'h1 ? valid_3_0 : _GEN_3243; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3567 = unuse_way == 3'h1 ? valid_3_1 : _GEN_3244; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3568 = unuse_way == 3'h1 ? valid_3_2 : _GEN_3245; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3569 = unuse_way == 3'h1 ? valid_3_3 : _GEN_3246; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3570 = unuse_way == 3'h1 ? valid_3_4 : _GEN_3247; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3571 = unuse_way == 3'h1 ? valid_3_5 : _GEN_3248; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3572 = unuse_way == 3'h1 ? valid_3_6 : _GEN_3249; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3573 = unuse_way == 3'h1 ? valid_3_7 : _GEN_3250; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3574 = unuse_way == 3'h1 ? valid_3_8 : _GEN_3251; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3575 = unuse_way == 3'h1 ? valid_3_9 : _GEN_3252; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3576 = unuse_way == 3'h1 ? valid_3_10 : _GEN_3253; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3577 = unuse_way == 3'h1 ? valid_3_11 : _GEN_3254; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3578 = unuse_way == 3'h1 ? valid_3_12 : _GEN_3255; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3579 = unuse_way == 3'h1 ? valid_3_13 : _GEN_3256; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3580 = unuse_way == 3'h1 ? valid_3_14 : _GEN_3257; // @[d_cache.scala 168:34 32:26]
  wire  _GEN_3581 = unuse_way == 3'h1 ? valid_3_15 : _GEN_3258; // @[d_cache.scala 168:34 32:26]
  wire [511:0] _GEN_3582 = unuse_way == 3'h1 ? write_back_data : _GEN_3259; // @[d_cache.scala 168:34 44:34]
  wire [41:0] _GEN_3583 = unuse_way == 3'h1 ? {{10'd0}, write_back_addr} : _GEN_3260; // @[d_cache.scala 168:34 45:34]
  wire  _GEN_3584 = unuse_way == 3'h1 ? dirty_0_0 : _GEN_3293; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3585 = unuse_way == 3'h1 ? dirty_0_1 : _GEN_3294; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3586 = unuse_way == 3'h1 ? dirty_0_2 : _GEN_3295; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3587 = unuse_way == 3'h1 ? dirty_0_3 : _GEN_3296; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3588 = unuse_way == 3'h1 ? dirty_0_4 : _GEN_3297; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3589 = unuse_way == 3'h1 ? dirty_0_5 : _GEN_3298; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3590 = unuse_way == 3'h1 ? dirty_0_6 : _GEN_3299; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3591 = unuse_way == 3'h1 ? dirty_0_7 : _GEN_3300; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3592 = unuse_way == 3'h1 ? dirty_0_8 : _GEN_3301; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3593 = unuse_way == 3'h1 ? dirty_0_9 : _GEN_3302; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3594 = unuse_way == 3'h1 ? dirty_0_10 : _GEN_3303; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3595 = unuse_way == 3'h1 ? dirty_0_11 : _GEN_3304; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3596 = unuse_way == 3'h1 ? dirty_0_12 : _GEN_3305; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3597 = unuse_way == 3'h1 ? dirty_0_13 : _GEN_3306; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3598 = unuse_way == 3'h1 ? dirty_0_14 : _GEN_3307; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3599 = unuse_way == 3'h1 ? dirty_0_15 : _GEN_3308; // @[d_cache.scala 168:34 34:26]
  wire  _GEN_3600 = unuse_way == 3'h1 ? dirty_1_0 : _GEN_3325; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3601 = unuse_way == 3'h1 ? dirty_1_1 : _GEN_3326; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3602 = unuse_way == 3'h1 ? dirty_1_2 : _GEN_3327; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3603 = unuse_way == 3'h1 ? dirty_1_3 : _GEN_3328; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3604 = unuse_way == 3'h1 ? dirty_1_4 : _GEN_3329; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3605 = unuse_way == 3'h1 ? dirty_1_5 : _GEN_3330; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3606 = unuse_way == 3'h1 ? dirty_1_6 : _GEN_3331; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3607 = unuse_way == 3'h1 ? dirty_1_7 : _GEN_3332; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3608 = unuse_way == 3'h1 ? dirty_1_8 : _GEN_3333; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3609 = unuse_way == 3'h1 ? dirty_1_9 : _GEN_3334; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3610 = unuse_way == 3'h1 ? dirty_1_10 : _GEN_3335; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3611 = unuse_way == 3'h1 ? dirty_1_11 : _GEN_3336; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3612 = unuse_way == 3'h1 ? dirty_1_12 : _GEN_3337; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3613 = unuse_way == 3'h1 ? dirty_1_13 : _GEN_3338; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3614 = unuse_way == 3'h1 ? dirty_1_14 : _GEN_3339; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3615 = unuse_way == 3'h1 ? dirty_1_15 : _GEN_3340; // @[d_cache.scala 168:34 35:26]
  wire  _GEN_3616 = unuse_way == 3'h1 ? dirty_2_0 : _GEN_3341; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3617 = unuse_way == 3'h1 ? dirty_2_1 : _GEN_3342; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3618 = unuse_way == 3'h1 ? dirty_2_2 : _GEN_3343; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3619 = unuse_way == 3'h1 ? dirty_2_3 : _GEN_3344; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3620 = unuse_way == 3'h1 ? dirty_2_4 : _GEN_3345; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3621 = unuse_way == 3'h1 ? dirty_2_5 : _GEN_3346; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3622 = unuse_way == 3'h1 ? dirty_2_6 : _GEN_3347; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3623 = unuse_way == 3'h1 ? dirty_2_7 : _GEN_3348; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3624 = unuse_way == 3'h1 ? dirty_2_8 : _GEN_3349; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3625 = unuse_way == 3'h1 ? dirty_2_9 : _GEN_3350; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3626 = unuse_way == 3'h1 ? dirty_2_10 : _GEN_3351; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3627 = unuse_way == 3'h1 ? dirty_2_11 : _GEN_3352; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3628 = unuse_way == 3'h1 ? dirty_2_12 : _GEN_3353; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3629 = unuse_way == 3'h1 ? dirty_2_13 : _GEN_3354; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3630 = unuse_way == 3'h1 ? dirty_2_14 : _GEN_3355; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3631 = unuse_way == 3'h1 ? dirty_2_15 : _GEN_3356; // @[d_cache.scala 168:34 36:26]
  wire  _GEN_3632 = unuse_way == 3'h1 ? dirty_3_0 : _GEN_3357; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3633 = unuse_way == 3'h1 ? dirty_3_1 : _GEN_3358; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3634 = unuse_way == 3'h1 ? dirty_3_2 : _GEN_3359; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3635 = unuse_way == 3'h1 ? dirty_3_3 : _GEN_3360; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3636 = unuse_way == 3'h1 ? dirty_3_4 : _GEN_3361; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3637 = unuse_way == 3'h1 ? dirty_3_5 : _GEN_3362; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3638 = unuse_way == 3'h1 ? dirty_3_6 : _GEN_3363; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3639 = unuse_way == 3'h1 ? dirty_3_7 : _GEN_3364; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3640 = unuse_way == 3'h1 ? dirty_3_8 : _GEN_3365; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3641 = unuse_way == 3'h1 ? dirty_3_9 : _GEN_3366; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3642 = unuse_way == 3'h1 ? dirty_3_10 : _GEN_3367; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3643 = unuse_way == 3'h1 ? dirty_3_11 : _GEN_3368; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3644 = unuse_way == 3'h1 ? dirty_3_12 : _GEN_3369; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3645 = unuse_way == 3'h1 ? dirty_3_13 : _GEN_3370; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3646 = unuse_way == 3'h1 ? dirty_3_14 : _GEN_3371; // @[d_cache.scala 168:34 37:26]
  wire  _GEN_3647 = unuse_way == 3'h1 ? dirty_3_15 : _GEN_3372; // @[d_cache.scala 168:34 37:26]
  wire [511:0] _write_back_data_T = {{64'd0}, write_back_data[511:64]}; // @[d_cache.scala 266:52]
  wire [511:0] _GEN_3648 = io_from_axi_wready ? _write_back_data_T : write_back_data; // @[d_cache.scala 265:37 266:33 44:34]
  wire [3:0] _GEN_3649 = io_from_axi_bvalid ? 4'h1 : state; // @[d_cache.scala 268:37 269:23 100:24]
  wire [3:0] _GEN_3650 = io_from_axi_rvalid ? 4'h0 : state; // @[d_cache.scala 273:37 274:23 100:24]
  wire [3:0] _GEN_3651 = 4'h8 == state ? _GEN_670 : state; // @[d_cache.scala 105:18 100:24]
  wire [3:0] _GEN_3652 = 4'h7 == state ? _GEN_3650 : _GEN_3651; // @[d_cache.scala 105:18]
  wire [511:0] _GEN_3653 = 4'h6 == state ? _GEN_3648 : write_back_data; // @[d_cache.scala 105:18 44:34]
  wire [3:0] _GEN_3654 = 4'h6 == state ? _GEN_3649 : _GEN_3652; // @[d_cache.scala 105:18]
  wire [3:0] _GEN_3655 = 4'h5 == state ? _GEN_3373 : _GEN_3654; // @[d_cache.scala 105:18]
  wire [511:0] _GEN_3656 = 4'h5 == state ? _GEN_3374 : ram_0_0; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3657 = 4'h5 == state ? _GEN_3375 : ram_0_1; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3658 = 4'h5 == state ? _GEN_3376 : ram_0_2; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3659 = 4'h5 == state ? _GEN_3377 : ram_0_3; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3660 = 4'h5 == state ? _GEN_3378 : ram_0_4; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3661 = 4'h5 == state ? _GEN_3379 : ram_0_5; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3662 = 4'h5 == state ? _GEN_3380 : ram_0_6; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3663 = 4'h5 == state ? _GEN_3381 : ram_0_7; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3664 = 4'h5 == state ? _GEN_3382 : ram_0_8; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3665 = 4'h5 == state ? _GEN_3383 : ram_0_9; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3666 = 4'h5 == state ? _GEN_3384 : ram_0_10; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3667 = 4'h5 == state ? _GEN_3385 : ram_0_11; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3668 = 4'h5 == state ? _GEN_3386 : ram_0_12; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3669 = 4'h5 == state ? _GEN_3387 : ram_0_13; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3670 = 4'h5 == state ? _GEN_3388 : ram_0_14; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3671 = 4'h5 == state ? _GEN_3389 : ram_0_15; // @[d_cache.scala 105:18 19:24]
  wire [31:0] _GEN_3672 = 4'h5 == state ? _GEN_3390 : tag_0_0; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3673 = 4'h5 == state ? _GEN_3391 : tag_0_1; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3674 = 4'h5 == state ? _GEN_3392 : tag_0_2; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3675 = 4'h5 == state ? _GEN_3393 : tag_0_3; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3676 = 4'h5 == state ? _GEN_3394 : tag_0_4; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3677 = 4'h5 == state ? _GEN_3395 : tag_0_5; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3678 = 4'h5 == state ? _GEN_3396 : tag_0_6; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3679 = 4'h5 == state ? _GEN_3397 : tag_0_7; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3680 = 4'h5 == state ? _GEN_3398 : tag_0_8; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3681 = 4'h5 == state ? _GEN_3399 : tag_0_9; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3682 = 4'h5 == state ? _GEN_3400 : tag_0_10; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3683 = 4'h5 == state ? _GEN_3401 : tag_0_11; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3684 = 4'h5 == state ? _GEN_3402 : tag_0_12; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3685 = 4'h5 == state ? _GEN_3403 : tag_0_13; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3686 = 4'h5 == state ? _GEN_3404 : tag_0_14; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3687 = 4'h5 == state ? _GEN_3405 : tag_0_15; // @[d_cache.scala 105:18 24:24]
  wire  _GEN_3688 = 4'h5 == state ? _GEN_3406 : valid_0_0; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3689 = 4'h5 == state ? _GEN_3407 : valid_0_1; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3690 = 4'h5 == state ? _GEN_3408 : valid_0_2; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3691 = 4'h5 == state ? _GEN_3409 : valid_0_3; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3692 = 4'h5 == state ? _GEN_3410 : valid_0_4; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3693 = 4'h5 == state ? _GEN_3411 : valid_0_5; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3694 = 4'h5 == state ? _GEN_3412 : valid_0_6; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3695 = 4'h5 == state ? _GEN_3413 : valid_0_7; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3696 = 4'h5 == state ? _GEN_3414 : valid_0_8; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3697 = 4'h5 == state ? _GEN_3415 : valid_0_9; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3698 = 4'h5 == state ? _GEN_3416 : valid_0_10; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3699 = 4'h5 == state ? _GEN_3417 : valid_0_11; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3700 = 4'h5 == state ? _GEN_3418 : valid_0_12; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3701 = 4'h5 == state ? _GEN_3419 : valid_0_13; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3702 = 4'h5 == state ? _GEN_3420 : valid_0_14; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3703 = 4'h5 == state ? _GEN_3421 : valid_0_15; // @[d_cache.scala 105:18 29:26]
  wire [7:0] _GEN_3704 = 4'h5 == state ? _GEN_3422 : quene_0; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3705 = 4'h5 == state ? _GEN_3423 : quene_1; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3706 = 4'h5 == state ? _GEN_3424 : quene_2; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3707 = 4'h5 == state ? _GEN_3425 : quene_3; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3708 = 4'h5 == state ? _GEN_3426 : quene_4; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3709 = 4'h5 == state ? _GEN_3427 : quene_5; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3710 = 4'h5 == state ? _GEN_3428 : quene_6; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3711 = 4'h5 == state ? _GEN_3429 : quene_7; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3712 = 4'h5 == state ? _GEN_3430 : quene_8; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3713 = 4'h5 == state ? _GEN_3431 : quene_9; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3714 = 4'h5 == state ? _GEN_3432 : quene_10; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3715 = 4'h5 == state ? _GEN_3433 : quene_11; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3716 = 4'h5 == state ? _GEN_3434 : quene_12; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3717 = 4'h5 == state ? _GEN_3435 : quene_13; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3718 = 4'h5 == state ? _GEN_3436 : quene_14; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3719 = 4'h5 == state ? _GEN_3437 : quene_15; // @[d_cache.scala 105:18 52:24]
  wire [511:0] _GEN_3720 = 4'h5 == state ? _GEN_3438 : ram_1_0; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3721 = 4'h5 == state ? _GEN_3439 : ram_1_1; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3722 = 4'h5 == state ? _GEN_3440 : ram_1_2; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3723 = 4'h5 == state ? _GEN_3441 : ram_1_3; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3724 = 4'h5 == state ? _GEN_3442 : ram_1_4; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3725 = 4'h5 == state ? _GEN_3443 : ram_1_5; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3726 = 4'h5 == state ? _GEN_3444 : ram_1_6; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3727 = 4'h5 == state ? _GEN_3445 : ram_1_7; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3728 = 4'h5 == state ? _GEN_3446 : ram_1_8; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3729 = 4'h5 == state ? _GEN_3447 : ram_1_9; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3730 = 4'h5 == state ? _GEN_3448 : ram_1_10; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3731 = 4'h5 == state ? _GEN_3449 : ram_1_11; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3732 = 4'h5 == state ? _GEN_3450 : ram_1_12; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3733 = 4'h5 == state ? _GEN_3451 : ram_1_13; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3734 = 4'h5 == state ? _GEN_3452 : ram_1_14; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3735 = 4'h5 == state ? _GEN_3453 : ram_1_15; // @[d_cache.scala 105:18 20:24]
  wire [31:0] _GEN_3736 = 4'h5 == state ? _GEN_3454 : tag_1_0; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3737 = 4'h5 == state ? _GEN_3455 : tag_1_1; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3738 = 4'h5 == state ? _GEN_3456 : tag_1_2; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3739 = 4'h5 == state ? _GEN_3457 : tag_1_3; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3740 = 4'h5 == state ? _GEN_3458 : tag_1_4; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3741 = 4'h5 == state ? _GEN_3459 : tag_1_5; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3742 = 4'h5 == state ? _GEN_3460 : tag_1_6; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3743 = 4'h5 == state ? _GEN_3461 : tag_1_7; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3744 = 4'h5 == state ? _GEN_3462 : tag_1_8; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3745 = 4'h5 == state ? _GEN_3463 : tag_1_9; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3746 = 4'h5 == state ? _GEN_3464 : tag_1_10; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3747 = 4'h5 == state ? _GEN_3465 : tag_1_11; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3748 = 4'h5 == state ? _GEN_3466 : tag_1_12; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3749 = 4'h5 == state ? _GEN_3467 : tag_1_13; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3750 = 4'h5 == state ? _GEN_3468 : tag_1_14; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_3751 = 4'h5 == state ? _GEN_3469 : tag_1_15; // @[d_cache.scala 105:18 25:24]
  wire  _GEN_3752 = 4'h5 == state ? _GEN_3470 : valid_1_0; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3753 = 4'h5 == state ? _GEN_3471 : valid_1_1; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3754 = 4'h5 == state ? _GEN_3472 : valid_1_2; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3755 = 4'h5 == state ? _GEN_3473 : valid_1_3; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3756 = 4'h5 == state ? _GEN_3474 : valid_1_4; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3757 = 4'h5 == state ? _GEN_3475 : valid_1_5; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3758 = 4'h5 == state ? _GEN_3476 : valid_1_6; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3759 = 4'h5 == state ? _GEN_3477 : valid_1_7; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3760 = 4'h5 == state ? _GEN_3478 : valid_1_8; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3761 = 4'h5 == state ? _GEN_3479 : valid_1_9; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3762 = 4'h5 == state ? _GEN_3480 : valid_1_10; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3763 = 4'h5 == state ? _GEN_3481 : valid_1_11; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3764 = 4'h5 == state ? _GEN_3482 : valid_1_12; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3765 = 4'h5 == state ? _GEN_3483 : valid_1_13; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3766 = 4'h5 == state ? _GEN_3484 : valid_1_14; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_3767 = 4'h5 == state ? _GEN_3485 : valid_1_15; // @[d_cache.scala 105:18 30:26]
  wire [511:0] _GEN_3768 = 4'h5 == state ? _GEN_3486 : ram_2_0; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3769 = 4'h5 == state ? _GEN_3487 : ram_2_1; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3770 = 4'h5 == state ? _GEN_3488 : ram_2_2; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3771 = 4'h5 == state ? _GEN_3489 : ram_2_3; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3772 = 4'h5 == state ? _GEN_3490 : ram_2_4; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3773 = 4'h5 == state ? _GEN_3491 : ram_2_5; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3774 = 4'h5 == state ? _GEN_3492 : ram_2_6; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3775 = 4'h5 == state ? _GEN_3493 : ram_2_7; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3776 = 4'h5 == state ? _GEN_3494 : ram_2_8; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3777 = 4'h5 == state ? _GEN_3495 : ram_2_9; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3778 = 4'h5 == state ? _GEN_3496 : ram_2_10; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3779 = 4'h5 == state ? _GEN_3497 : ram_2_11; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3780 = 4'h5 == state ? _GEN_3498 : ram_2_12; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3781 = 4'h5 == state ? _GEN_3499 : ram_2_13; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3782 = 4'h5 == state ? _GEN_3500 : ram_2_14; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_3783 = 4'h5 == state ? _GEN_3501 : ram_2_15; // @[d_cache.scala 105:18 21:24]
  wire [31:0] _GEN_3784 = 4'h5 == state ? _GEN_3502 : tag_2_0; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3785 = 4'h5 == state ? _GEN_3503 : tag_2_1; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3786 = 4'h5 == state ? _GEN_3504 : tag_2_2; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3787 = 4'h5 == state ? _GEN_3505 : tag_2_3; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3788 = 4'h5 == state ? _GEN_3506 : tag_2_4; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3789 = 4'h5 == state ? _GEN_3507 : tag_2_5; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3790 = 4'h5 == state ? _GEN_3508 : tag_2_6; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3791 = 4'h5 == state ? _GEN_3509 : tag_2_7; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3792 = 4'h5 == state ? _GEN_3510 : tag_2_8; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3793 = 4'h5 == state ? _GEN_3511 : tag_2_9; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3794 = 4'h5 == state ? _GEN_3512 : tag_2_10; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3795 = 4'h5 == state ? _GEN_3513 : tag_2_11; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3796 = 4'h5 == state ? _GEN_3514 : tag_2_12; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3797 = 4'h5 == state ? _GEN_3515 : tag_2_13; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3798 = 4'h5 == state ? _GEN_3516 : tag_2_14; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_3799 = 4'h5 == state ? _GEN_3517 : tag_2_15; // @[d_cache.scala 105:18 26:24]
  wire  _GEN_3800 = 4'h5 == state ? _GEN_3518 : valid_2_0; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3801 = 4'h5 == state ? _GEN_3519 : valid_2_1; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3802 = 4'h5 == state ? _GEN_3520 : valid_2_2; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3803 = 4'h5 == state ? _GEN_3521 : valid_2_3; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3804 = 4'h5 == state ? _GEN_3522 : valid_2_4; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3805 = 4'h5 == state ? _GEN_3523 : valid_2_5; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3806 = 4'h5 == state ? _GEN_3524 : valid_2_6; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3807 = 4'h5 == state ? _GEN_3525 : valid_2_7; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3808 = 4'h5 == state ? _GEN_3526 : valid_2_8; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3809 = 4'h5 == state ? _GEN_3527 : valid_2_9; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3810 = 4'h5 == state ? _GEN_3528 : valid_2_10; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3811 = 4'h5 == state ? _GEN_3529 : valid_2_11; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3812 = 4'h5 == state ? _GEN_3530 : valid_2_12; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3813 = 4'h5 == state ? _GEN_3531 : valid_2_13; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3814 = 4'h5 == state ? _GEN_3532 : valid_2_14; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_3815 = 4'h5 == state ? _GEN_3533 : valid_2_15; // @[d_cache.scala 105:18 31:26]
  wire [511:0] _GEN_3816 = 4'h5 == state ? _GEN_3534 : ram_3_0; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3817 = 4'h5 == state ? _GEN_3535 : ram_3_1; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3818 = 4'h5 == state ? _GEN_3536 : ram_3_2; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3819 = 4'h5 == state ? _GEN_3537 : ram_3_3; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3820 = 4'h5 == state ? _GEN_3538 : ram_3_4; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3821 = 4'h5 == state ? _GEN_3539 : ram_3_5; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3822 = 4'h5 == state ? _GEN_3540 : ram_3_6; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3823 = 4'h5 == state ? _GEN_3541 : ram_3_7; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3824 = 4'h5 == state ? _GEN_3542 : ram_3_8; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3825 = 4'h5 == state ? _GEN_3543 : ram_3_9; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3826 = 4'h5 == state ? _GEN_3544 : ram_3_10; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3827 = 4'h5 == state ? _GEN_3545 : ram_3_11; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3828 = 4'h5 == state ? _GEN_3546 : ram_3_12; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3829 = 4'h5 == state ? _GEN_3547 : ram_3_13; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3830 = 4'h5 == state ? _GEN_3548 : ram_3_14; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_3831 = 4'h5 == state ? _GEN_3549 : ram_3_15; // @[d_cache.scala 105:18 22:24]
  wire [31:0] _GEN_3832 = 4'h5 == state ? _GEN_3550 : tag_3_0; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3833 = 4'h5 == state ? _GEN_3551 : tag_3_1; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3834 = 4'h5 == state ? _GEN_3552 : tag_3_2; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3835 = 4'h5 == state ? _GEN_3553 : tag_3_3; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3836 = 4'h5 == state ? _GEN_3554 : tag_3_4; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3837 = 4'h5 == state ? _GEN_3555 : tag_3_5; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3838 = 4'h5 == state ? _GEN_3556 : tag_3_6; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3839 = 4'h5 == state ? _GEN_3557 : tag_3_7; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3840 = 4'h5 == state ? _GEN_3558 : tag_3_8; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3841 = 4'h5 == state ? _GEN_3559 : tag_3_9; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3842 = 4'h5 == state ? _GEN_3560 : tag_3_10; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3843 = 4'h5 == state ? _GEN_3561 : tag_3_11; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3844 = 4'h5 == state ? _GEN_3562 : tag_3_12; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3845 = 4'h5 == state ? _GEN_3563 : tag_3_13; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3846 = 4'h5 == state ? _GEN_3564 : tag_3_14; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_3847 = 4'h5 == state ? _GEN_3565 : tag_3_15; // @[d_cache.scala 105:18 27:24]
  wire  _GEN_3848 = 4'h5 == state ? _GEN_3566 : valid_3_0; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3849 = 4'h5 == state ? _GEN_3567 : valid_3_1; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3850 = 4'h5 == state ? _GEN_3568 : valid_3_2; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3851 = 4'h5 == state ? _GEN_3569 : valid_3_3; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3852 = 4'h5 == state ? _GEN_3570 : valid_3_4; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3853 = 4'h5 == state ? _GEN_3571 : valid_3_5; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3854 = 4'h5 == state ? _GEN_3572 : valid_3_6; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3855 = 4'h5 == state ? _GEN_3573 : valid_3_7; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3856 = 4'h5 == state ? _GEN_3574 : valid_3_8; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3857 = 4'h5 == state ? _GEN_3575 : valid_3_9; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3858 = 4'h5 == state ? _GEN_3576 : valid_3_10; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3859 = 4'h5 == state ? _GEN_3577 : valid_3_11; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3860 = 4'h5 == state ? _GEN_3578 : valid_3_12; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3861 = 4'h5 == state ? _GEN_3579 : valid_3_13; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3862 = 4'h5 == state ? _GEN_3580 : valid_3_14; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_3863 = 4'h5 == state ? _GEN_3581 : valid_3_15; // @[d_cache.scala 105:18 32:26]
  wire [511:0] _GEN_3864 = 4'h5 == state ? _GEN_3582 : _GEN_3653; // @[d_cache.scala 105:18]
  wire [41:0] _GEN_3865 = 4'h5 == state ? _GEN_3583 : {{10'd0}, write_back_addr}; // @[d_cache.scala 105:18 45:34]
  wire  _GEN_3866 = 4'h5 == state ? _GEN_3584 : dirty_0_0; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3867 = 4'h5 == state ? _GEN_3585 : dirty_0_1; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3868 = 4'h5 == state ? _GEN_3586 : dirty_0_2; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3869 = 4'h5 == state ? _GEN_3587 : dirty_0_3; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3870 = 4'h5 == state ? _GEN_3588 : dirty_0_4; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3871 = 4'h5 == state ? _GEN_3589 : dirty_0_5; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3872 = 4'h5 == state ? _GEN_3590 : dirty_0_6; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3873 = 4'h5 == state ? _GEN_3591 : dirty_0_7; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3874 = 4'h5 == state ? _GEN_3592 : dirty_0_8; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3875 = 4'h5 == state ? _GEN_3593 : dirty_0_9; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3876 = 4'h5 == state ? _GEN_3594 : dirty_0_10; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3877 = 4'h5 == state ? _GEN_3595 : dirty_0_11; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3878 = 4'h5 == state ? _GEN_3596 : dirty_0_12; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3879 = 4'h5 == state ? _GEN_3597 : dirty_0_13; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3880 = 4'h5 == state ? _GEN_3598 : dirty_0_14; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3881 = 4'h5 == state ? _GEN_3599 : dirty_0_15; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_3882 = 4'h5 == state ? _GEN_3600 : dirty_1_0; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3883 = 4'h5 == state ? _GEN_3601 : dirty_1_1; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3884 = 4'h5 == state ? _GEN_3602 : dirty_1_2; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3885 = 4'h5 == state ? _GEN_3603 : dirty_1_3; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3886 = 4'h5 == state ? _GEN_3604 : dirty_1_4; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3887 = 4'h5 == state ? _GEN_3605 : dirty_1_5; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3888 = 4'h5 == state ? _GEN_3606 : dirty_1_6; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3889 = 4'h5 == state ? _GEN_3607 : dirty_1_7; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3890 = 4'h5 == state ? _GEN_3608 : dirty_1_8; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3891 = 4'h5 == state ? _GEN_3609 : dirty_1_9; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3892 = 4'h5 == state ? _GEN_3610 : dirty_1_10; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3893 = 4'h5 == state ? _GEN_3611 : dirty_1_11; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3894 = 4'h5 == state ? _GEN_3612 : dirty_1_12; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3895 = 4'h5 == state ? _GEN_3613 : dirty_1_13; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3896 = 4'h5 == state ? _GEN_3614 : dirty_1_14; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3897 = 4'h5 == state ? _GEN_3615 : dirty_1_15; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_3898 = 4'h5 == state ? _GEN_3616 : dirty_2_0; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3899 = 4'h5 == state ? _GEN_3617 : dirty_2_1; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3900 = 4'h5 == state ? _GEN_3618 : dirty_2_2; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3901 = 4'h5 == state ? _GEN_3619 : dirty_2_3; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3902 = 4'h5 == state ? _GEN_3620 : dirty_2_4; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3903 = 4'h5 == state ? _GEN_3621 : dirty_2_5; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3904 = 4'h5 == state ? _GEN_3622 : dirty_2_6; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3905 = 4'h5 == state ? _GEN_3623 : dirty_2_7; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3906 = 4'h5 == state ? _GEN_3624 : dirty_2_8; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3907 = 4'h5 == state ? _GEN_3625 : dirty_2_9; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3908 = 4'h5 == state ? _GEN_3626 : dirty_2_10; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3909 = 4'h5 == state ? _GEN_3627 : dirty_2_11; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3910 = 4'h5 == state ? _GEN_3628 : dirty_2_12; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3911 = 4'h5 == state ? _GEN_3629 : dirty_2_13; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3912 = 4'h5 == state ? _GEN_3630 : dirty_2_14; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3913 = 4'h5 == state ? _GEN_3631 : dirty_2_15; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_3914 = 4'h5 == state ? _GEN_3632 : dirty_3_0; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3915 = 4'h5 == state ? _GEN_3633 : dirty_3_1; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3916 = 4'h5 == state ? _GEN_3634 : dirty_3_2; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3917 = 4'h5 == state ? _GEN_3635 : dirty_3_3; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3918 = 4'h5 == state ? _GEN_3636 : dirty_3_4; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3919 = 4'h5 == state ? _GEN_3637 : dirty_3_5; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3920 = 4'h5 == state ? _GEN_3638 : dirty_3_6; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3921 = 4'h5 == state ? _GEN_3639 : dirty_3_7; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3922 = 4'h5 == state ? _GEN_3640 : dirty_3_8; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3923 = 4'h5 == state ? _GEN_3641 : dirty_3_9; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3924 = 4'h5 == state ? _GEN_3642 : dirty_3_10; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3925 = 4'h5 == state ? _GEN_3643 : dirty_3_11; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3926 = 4'h5 == state ? _GEN_3644 : dirty_3_12; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3927 = 4'h5 == state ? _GEN_3645 : dirty_3_13; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3928 = 4'h5 == state ? _GEN_3646 : dirty_3_14; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_3929 = 4'h5 == state ? _GEN_3647 : dirty_3_15; // @[d_cache.scala 105:18 37:26]
  wire [3:0] _GEN_3930 = 4'h4 == state ? _GEN_670 : _GEN_3655; // @[d_cache.scala 105:18]
  wire [511:0] _GEN_3931 = 4'h4 == state ? ram_0_0 : _GEN_3656; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3932 = 4'h4 == state ? ram_0_1 : _GEN_3657; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3933 = 4'h4 == state ? ram_0_2 : _GEN_3658; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3934 = 4'h4 == state ? ram_0_3 : _GEN_3659; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3935 = 4'h4 == state ? ram_0_4 : _GEN_3660; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3936 = 4'h4 == state ? ram_0_5 : _GEN_3661; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3937 = 4'h4 == state ? ram_0_6 : _GEN_3662; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3938 = 4'h4 == state ? ram_0_7 : _GEN_3663; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3939 = 4'h4 == state ? ram_0_8 : _GEN_3664; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3940 = 4'h4 == state ? ram_0_9 : _GEN_3665; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3941 = 4'h4 == state ? ram_0_10 : _GEN_3666; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3942 = 4'h4 == state ? ram_0_11 : _GEN_3667; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3943 = 4'h4 == state ? ram_0_12 : _GEN_3668; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3944 = 4'h4 == state ? ram_0_13 : _GEN_3669; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3945 = 4'h4 == state ? ram_0_14 : _GEN_3670; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_3946 = 4'h4 == state ? ram_0_15 : _GEN_3671; // @[d_cache.scala 105:18 19:24]
  wire [31:0] _GEN_3947 = 4'h4 == state ? tag_0_0 : _GEN_3672; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3948 = 4'h4 == state ? tag_0_1 : _GEN_3673; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3949 = 4'h4 == state ? tag_0_2 : _GEN_3674; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3950 = 4'h4 == state ? tag_0_3 : _GEN_3675; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3951 = 4'h4 == state ? tag_0_4 : _GEN_3676; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3952 = 4'h4 == state ? tag_0_5 : _GEN_3677; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3953 = 4'h4 == state ? tag_0_6 : _GEN_3678; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3954 = 4'h4 == state ? tag_0_7 : _GEN_3679; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3955 = 4'h4 == state ? tag_0_8 : _GEN_3680; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3956 = 4'h4 == state ? tag_0_9 : _GEN_3681; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3957 = 4'h4 == state ? tag_0_10 : _GEN_3682; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3958 = 4'h4 == state ? tag_0_11 : _GEN_3683; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3959 = 4'h4 == state ? tag_0_12 : _GEN_3684; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3960 = 4'h4 == state ? tag_0_13 : _GEN_3685; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3961 = 4'h4 == state ? tag_0_14 : _GEN_3686; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_3962 = 4'h4 == state ? tag_0_15 : _GEN_3687; // @[d_cache.scala 105:18 24:24]
  wire  _GEN_3963 = 4'h4 == state ? valid_0_0 : _GEN_3688; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3964 = 4'h4 == state ? valid_0_1 : _GEN_3689; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3965 = 4'h4 == state ? valid_0_2 : _GEN_3690; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3966 = 4'h4 == state ? valid_0_3 : _GEN_3691; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3967 = 4'h4 == state ? valid_0_4 : _GEN_3692; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3968 = 4'h4 == state ? valid_0_5 : _GEN_3693; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3969 = 4'h4 == state ? valid_0_6 : _GEN_3694; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3970 = 4'h4 == state ? valid_0_7 : _GEN_3695; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3971 = 4'h4 == state ? valid_0_8 : _GEN_3696; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3972 = 4'h4 == state ? valid_0_9 : _GEN_3697; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3973 = 4'h4 == state ? valid_0_10 : _GEN_3698; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3974 = 4'h4 == state ? valid_0_11 : _GEN_3699; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3975 = 4'h4 == state ? valid_0_12 : _GEN_3700; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3976 = 4'h4 == state ? valid_0_13 : _GEN_3701; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3977 = 4'h4 == state ? valid_0_14 : _GEN_3702; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_3978 = 4'h4 == state ? valid_0_15 : _GEN_3703; // @[d_cache.scala 105:18 29:26]
  wire [7:0] _GEN_3979 = 4'h4 == state ? quene_0 : _GEN_3704; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3980 = 4'h4 == state ? quene_1 : _GEN_3705; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3981 = 4'h4 == state ? quene_2 : _GEN_3706; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3982 = 4'h4 == state ? quene_3 : _GEN_3707; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3983 = 4'h4 == state ? quene_4 : _GEN_3708; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3984 = 4'h4 == state ? quene_5 : _GEN_3709; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3985 = 4'h4 == state ? quene_6 : _GEN_3710; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3986 = 4'h4 == state ? quene_7 : _GEN_3711; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3987 = 4'h4 == state ? quene_8 : _GEN_3712; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3988 = 4'h4 == state ? quene_9 : _GEN_3713; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3989 = 4'h4 == state ? quene_10 : _GEN_3714; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3990 = 4'h4 == state ? quene_11 : _GEN_3715; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3991 = 4'h4 == state ? quene_12 : _GEN_3716; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3992 = 4'h4 == state ? quene_13 : _GEN_3717; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3993 = 4'h4 == state ? quene_14 : _GEN_3718; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_3994 = 4'h4 == state ? quene_15 : _GEN_3719; // @[d_cache.scala 105:18 52:24]
  wire [511:0] _GEN_3995 = 4'h4 == state ? ram_1_0 : _GEN_3720; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3996 = 4'h4 == state ? ram_1_1 : _GEN_3721; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3997 = 4'h4 == state ? ram_1_2 : _GEN_3722; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3998 = 4'h4 == state ? ram_1_3 : _GEN_3723; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_3999 = 4'h4 == state ? ram_1_4 : _GEN_3724; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4000 = 4'h4 == state ? ram_1_5 : _GEN_3725; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4001 = 4'h4 == state ? ram_1_6 : _GEN_3726; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4002 = 4'h4 == state ? ram_1_7 : _GEN_3727; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4003 = 4'h4 == state ? ram_1_8 : _GEN_3728; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4004 = 4'h4 == state ? ram_1_9 : _GEN_3729; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4005 = 4'h4 == state ? ram_1_10 : _GEN_3730; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4006 = 4'h4 == state ? ram_1_11 : _GEN_3731; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4007 = 4'h4 == state ? ram_1_12 : _GEN_3732; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4008 = 4'h4 == state ? ram_1_13 : _GEN_3733; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4009 = 4'h4 == state ? ram_1_14 : _GEN_3734; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4010 = 4'h4 == state ? ram_1_15 : _GEN_3735; // @[d_cache.scala 105:18 20:24]
  wire [31:0] _GEN_4011 = 4'h4 == state ? tag_1_0 : _GEN_3736; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4012 = 4'h4 == state ? tag_1_1 : _GEN_3737; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4013 = 4'h4 == state ? tag_1_2 : _GEN_3738; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4014 = 4'h4 == state ? tag_1_3 : _GEN_3739; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4015 = 4'h4 == state ? tag_1_4 : _GEN_3740; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4016 = 4'h4 == state ? tag_1_5 : _GEN_3741; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4017 = 4'h4 == state ? tag_1_6 : _GEN_3742; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4018 = 4'h4 == state ? tag_1_7 : _GEN_3743; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4019 = 4'h4 == state ? tag_1_8 : _GEN_3744; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4020 = 4'h4 == state ? tag_1_9 : _GEN_3745; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4021 = 4'h4 == state ? tag_1_10 : _GEN_3746; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4022 = 4'h4 == state ? tag_1_11 : _GEN_3747; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4023 = 4'h4 == state ? tag_1_12 : _GEN_3748; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4024 = 4'h4 == state ? tag_1_13 : _GEN_3749; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4025 = 4'h4 == state ? tag_1_14 : _GEN_3750; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4026 = 4'h4 == state ? tag_1_15 : _GEN_3751; // @[d_cache.scala 105:18 25:24]
  wire  _GEN_4027 = 4'h4 == state ? valid_1_0 : _GEN_3752; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4028 = 4'h4 == state ? valid_1_1 : _GEN_3753; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4029 = 4'h4 == state ? valid_1_2 : _GEN_3754; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4030 = 4'h4 == state ? valid_1_3 : _GEN_3755; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4031 = 4'h4 == state ? valid_1_4 : _GEN_3756; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4032 = 4'h4 == state ? valid_1_5 : _GEN_3757; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4033 = 4'h4 == state ? valid_1_6 : _GEN_3758; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4034 = 4'h4 == state ? valid_1_7 : _GEN_3759; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4035 = 4'h4 == state ? valid_1_8 : _GEN_3760; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4036 = 4'h4 == state ? valid_1_9 : _GEN_3761; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4037 = 4'h4 == state ? valid_1_10 : _GEN_3762; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4038 = 4'h4 == state ? valid_1_11 : _GEN_3763; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4039 = 4'h4 == state ? valid_1_12 : _GEN_3764; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4040 = 4'h4 == state ? valid_1_13 : _GEN_3765; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4041 = 4'h4 == state ? valid_1_14 : _GEN_3766; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4042 = 4'h4 == state ? valid_1_15 : _GEN_3767; // @[d_cache.scala 105:18 30:26]
  wire [511:0] _GEN_4043 = 4'h4 == state ? ram_2_0 : _GEN_3768; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4044 = 4'h4 == state ? ram_2_1 : _GEN_3769; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4045 = 4'h4 == state ? ram_2_2 : _GEN_3770; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4046 = 4'h4 == state ? ram_2_3 : _GEN_3771; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4047 = 4'h4 == state ? ram_2_4 : _GEN_3772; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4048 = 4'h4 == state ? ram_2_5 : _GEN_3773; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4049 = 4'h4 == state ? ram_2_6 : _GEN_3774; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4050 = 4'h4 == state ? ram_2_7 : _GEN_3775; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4051 = 4'h4 == state ? ram_2_8 : _GEN_3776; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4052 = 4'h4 == state ? ram_2_9 : _GEN_3777; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4053 = 4'h4 == state ? ram_2_10 : _GEN_3778; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4054 = 4'h4 == state ? ram_2_11 : _GEN_3779; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4055 = 4'h4 == state ? ram_2_12 : _GEN_3780; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4056 = 4'h4 == state ? ram_2_13 : _GEN_3781; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4057 = 4'h4 == state ? ram_2_14 : _GEN_3782; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4058 = 4'h4 == state ? ram_2_15 : _GEN_3783; // @[d_cache.scala 105:18 21:24]
  wire [31:0] _GEN_4059 = 4'h4 == state ? tag_2_0 : _GEN_3784; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4060 = 4'h4 == state ? tag_2_1 : _GEN_3785; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4061 = 4'h4 == state ? tag_2_2 : _GEN_3786; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4062 = 4'h4 == state ? tag_2_3 : _GEN_3787; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4063 = 4'h4 == state ? tag_2_4 : _GEN_3788; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4064 = 4'h4 == state ? tag_2_5 : _GEN_3789; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4065 = 4'h4 == state ? tag_2_6 : _GEN_3790; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4066 = 4'h4 == state ? tag_2_7 : _GEN_3791; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4067 = 4'h4 == state ? tag_2_8 : _GEN_3792; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4068 = 4'h4 == state ? tag_2_9 : _GEN_3793; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4069 = 4'h4 == state ? tag_2_10 : _GEN_3794; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4070 = 4'h4 == state ? tag_2_11 : _GEN_3795; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4071 = 4'h4 == state ? tag_2_12 : _GEN_3796; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4072 = 4'h4 == state ? tag_2_13 : _GEN_3797; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4073 = 4'h4 == state ? tag_2_14 : _GEN_3798; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4074 = 4'h4 == state ? tag_2_15 : _GEN_3799; // @[d_cache.scala 105:18 26:24]
  wire  _GEN_4075 = 4'h4 == state ? valid_2_0 : _GEN_3800; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4076 = 4'h4 == state ? valid_2_1 : _GEN_3801; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4077 = 4'h4 == state ? valid_2_2 : _GEN_3802; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4078 = 4'h4 == state ? valid_2_3 : _GEN_3803; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4079 = 4'h4 == state ? valid_2_4 : _GEN_3804; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4080 = 4'h4 == state ? valid_2_5 : _GEN_3805; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4081 = 4'h4 == state ? valid_2_6 : _GEN_3806; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4082 = 4'h4 == state ? valid_2_7 : _GEN_3807; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4083 = 4'h4 == state ? valid_2_8 : _GEN_3808; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4084 = 4'h4 == state ? valid_2_9 : _GEN_3809; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4085 = 4'h4 == state ? valid_2_10 : _GEN_3810; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4086 = 4'h4 == state ? valid_2_11 : _GEN_3811; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4087 = 4'h4 == state ? valid_2_12 : _GEN_3812; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4088 = 4'h4 == state ? valid_2_13 : _GEN_3813; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4089 = 4'h4 == state ? valid_2_14 : _GEN_3814; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4090 = 4'h4 == state ? valid_2_15 : _GEN_3815; // @[d_cache.scala 105:18 31:26]
  wire [511:0] _GEN_4091 = 4'h4 == state ? ram_3_0 : _GEN_3816; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4092 = 4'h4 == state ? ram_3_1 : _GEN_3817; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4093 = 4'h4 == state ? ram_3_2 : _GEN_3818; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4094 = 4'h4 == state ? ram_3_3 : _GEN_3819; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4095 = 4'h4 == state ? ram_3_4 : _GEN_3820; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4096 = 4'h4 == state ? ram_3_5 : _GEN_3821; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4097 = 4'h4 == state ? ram_3_6 : _GEN_3822; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4098 = 4'h4 == state ? ram_3_7 : _GEN_3823; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4099 = 4'h4 == state ? ram_3_8 : _GEN_3824; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4100 = 4'h4 == state ? ram_3_9 : _GEN_3825; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4101 = 4'h4 == state ? ram_3_10 : _GEN_3826; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4102 = 4'h4 == state ? ram_3_11 : _GEN_3827; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4103 = 4'h4 == state ? ram_3_12 : _GEN_3828; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4104 = 4'h4 == state ? ram_3_13 : _GEN_3829; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4105 = 4'h4 == state ? ram_3_14 : _GEN_3830; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4106 = 4'h4 == state ? ram_3_15 : _GEN_3831; // @[d_cache.scala 105:18 22:24]
  wire [31:0] _GEN_4107 = 4'h4 == state ? tag_3_0 : _GEN_3832; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4108 = 4'h4 == state ? tag_3_1 : _GEN_3833; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4109 = 4'h4 == state ? tag_3_2 : _GEN_3834; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4110 = 4'h4 == state ? tag_3_3 : _GEN_3835; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4111 = 4'h4 == state ? tag_3_4 : _GEN_3836; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4112 = 4'h4 == state ? tag_3_5 : _GEN_3837; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4113 = 4'h4 == state ? tag_3_6 : _GEN_3838; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4114 = 4'h4 == state ? tag_3_7 : _GEN_3839; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4115 = 4'h4 == state ? tag_3_8 : _GEN_3840; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4116 = 4'h4 == state ? tag_3_9 : _GEN_3841; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4117 = 4'h4 == state ? tag_3_10 : _GEN_3842; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4118 = 4'h4 == state ? tag_3_11 : _GEN_3843; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4119 = 4'h4 == state ? tag_3_12 : _GEN_3844; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4120 = 4'h4 == state ? tag_3_13 : _GEN_3845; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4121 = 4'h4 == state ? tag_3_14 : _GEN_3846; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4122 = 4'h4 == state ? tag_3_15 : _GEN_3847; // @[d_cache.scala 105:18 27:24]
  wire  _GEN_4123 = 4'h4 == state ? valid_3_0 : _GEN_3848; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4124 = 4'h4 == state ? valid_3_1 : _GEN_3849; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4125 = 4'h4 == state ? valid_3_2 : _GEN_3850; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4126 = 4'h4 == state ? valid_3_3 : _GEN_3851; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4127 = 4'h4 == state ? valid_3_4 : _GEN_3852; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4128 = 4'h4 == state ? valid_3_5 : _GEN_3853; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4129 = 4'h4 == state ? valid_3_6 : _GEN_3854; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4130 = 4'h4 == state ? valid_3_7 : _GEN_3855; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4131 = 4'h4 == state ? valid_3_8 : _GEN_3856; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4132 = 4'h4 == state ? valid_3_9 : _GEN_3857; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4133 = 4'h4 == state ? valid_3_10 : _GEN_3858; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4134 = 4'h4 == state ? valid_3_11 : _GEN_3859; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4135 = 4'h4 == state ? valid_3_12 : _GEN_3860; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4136 = 4'h4 == state ? valid_3_13 : _GEN_3861; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4137 = 4'h4 == state ? valid_3_14 : _GEN_3862; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4138 = 4'h4 == state ? valid_3_15 : _GEN_3863; // @[d_cache.scala 105:18 32:26]
  wire [511:0] _GEN_4139 = 4'h4 == state ? write_back_data : _GEN_3864; // @[d_cache.scala 105:18 44:34]
  wire [41:0] _GEN_4140 = 4'h4 == state ? {{10'd0}, write_back_addr} : _GEN_3865; // @[d_cache.scala 105:18 45:34]
  wire  _GEN_4141 = 4'h4 == state ? dirty_0_0 : _GEN_3866; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4142 = 4'h4 == state ? dirty_0_1 : _GEN_3867; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4143 = 4'h4 == state ? dirty_0_2 : _GEN_3868; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4144 = 4'h4 == state ? dirty_0_3 : _GEN_3869; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4145 = 4'h4 == state ? dirty_0_4 : _GEN_3870; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4146 = 4'h4 == state ? dirty_0_5 : _GEN_3871; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4147 = 4'h4 == state ? dirty_0_6 : _GEN_3872; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4148 = 4'h4 == state ? dirty_0_7 : _GEN_3873; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4149 = 4'h4 == state ? dirty_0_8 : _GEN_3874; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4150 = 4'h4 == state ? dirty_0_9 : _GEN_3875; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4151 = 4'h4 == state ? dirty_0_10 : _GEN_3876; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4152 = 4'h4 == state ? dirty_0_11 : _GEN_3877; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4153 = 4'h4 == state ? dirty_0_12 : _GEN_3878; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4154 = 4'h4 == state ? dirty_0_13 : _GEN_3879; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4155 = 4'h4 == state ? dirty_0_14 : _GEN_3880; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4156 = 4'h4 == state ? dirty_0_15 : _GEN_3881; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4157 = 4'h4 == state ? dirty_1_0 : _GEN_3882; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4158 = 4'h4 == state ? dirty_1_1 : _GEN_3883; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4159 = 4'h4 == state ? dirty_1_2 : _GEN_3884; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4160 = 4'h4 == state ? dirty_1_3 : _GEN_3885; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4161 = 4'h4 == state ? dirty_1_4 : _GEN_3886; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4162 = 4'h4 == state ? dirty_1_5 : _GEN_3887; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4163 = 4'h4 == state ? dirty_1_6 : _GEN_3888; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4164 = 4'h4 == state ? dirty_1_7 : _GEN_3889; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4165 = 4'h4 == state ? dirty_1_8 : _GEN_3890; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4166 = 4'h4 == state ? dirty_1_9 : _GEN_3891; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4167 = 4'h4 == state ? dirty_1_10 : _GEN_3892; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4168 = 4'h4 == state ? dirty_1_11 : _GEN_3893; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4169 = 4'h4 == state ? dirty_1_12 : _GEN_3894; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4170 = 4'h4 == state ? dirty_1_13 : _GEN_3895; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4171 = 4'h4 == state ? dirty_1_14 : _GEN_3896; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4172 = 4'h4 == state ? dirty_1_15 : _GEN_3897; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4173 = 4'h4 == state ? dirty_2_0 : _GEN_3898; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4174 = 4'h4 == state ? dirty_2_1 : _GEN_3899; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4175 = 4'h4 == state ? dirty_2_2 : _GEN_3900; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4176 = 4'h4 == state ? dirty_2_3 : _GEN_3901; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4177 = 4'h4 == state ? dirty_2_4 : _GEN_3902; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4178 = 4'h4 == state ? dirty_2_5 : _GEN_3903; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4179 = 4'h4 == state ? dirty_2_6 : _GEN_3904; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4180 = 4'h4 == state ? dirty_2_7 : _GEN_3905; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4181 = 4'h4 == state ? dirty_2_8 : _GEN_3906; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4182 = 4'h4 == state ? dirty_2_9 : _GEN_3907; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4183 = 4'h4 == state ? dirty_2_10 : _GEN_3908; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4184 = 4'h4 == state ? dirty_2_11 : _GEN_3909; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4185 = 4'h4 == state ? dirty_2_12 : _GEN_3910; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4186 = 4'h4 == state ? dirty_2_13 : _GEN_3911; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4187 = 4'h4 == state ? dirty_2_14 : _GEN_3912; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4188 = 4'h4 == state ? dirty_2_15 : _GEN_3913; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4189 = 4'h4 == state ? dirty_3_0 : _GEN_3914; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4190 = 4'h4 == state ? dirty_3_1 : _GEN_3915; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4191 = 4'h4 == state ? dirty_3_2 : _GEN_3916; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4192 = 4'h4 == state ? dirty_3_3 : _GEN_3917; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4193 = 4'h4 == state ? dirty_3_4 : _GEN_3918; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4194 = 4'h4 == state ? dirty_3_5 : _GEN_3919; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4195 = 4'h4 == state ? dirty_3_6 : _GEN_3920; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4196 = 4'h4 == state ? dirty_3_7 : _GEN_3921; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4197 = 4'h4 == state ? dirty_3_8 : _GEN_3922; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4198 = 4'h4 == state ? dirty_3_9 : _GEN_3923; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4199 = 4'h4 == state ? dirty_3_10 : _GEN_3924; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4200 = 4'h4 == state ? dirty_3_11 : _GEN_3925; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4201 = 4'h4 == state ? dirty_3_12 : _GEN_3926; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4202 = 4'h4 == state ? dirty_3_13 : _GEN_3927; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4203 = 4'h4 == state ? dirty_3_14 : _GEN_3928; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4204 = 4'h4 == state ? dirty_3_15 : _GEN_3929; // @[d_cache.scala 105:18 37:26]
  wire [63:0] _GEN_4205 = 4'h3 == state ? _GEN_660 : receive_data_0; // @[d_cache.scala 105:18 50:31]
  wire [63:0] _GEN_4206 = 4'h3 == state ? _GEN_661 : receive_data_1; // @[d_cache.scala 105:18 50:31]
  wire [63:0] _GEN_4207 = 4'h3 == state ? _GEN_662 : receive_data_2; // @[d_cache.scala 105:18 50:31]
  wire [63:0] _GEN_4208 = 4'h3 == state ? _GEN_663 : receive_data_3; // @[d_cache.scala 105:18 50:31]
  wire [63:0] _GEN_4209 = 4'h3 == state ? _GEN_664 : receive_data_4; // @[d_cache.scala 105:18 50:31]
  wire [63:0] _GEN_4210 = 4'h3 == state ? _GEN_665 : receive_data_5; // @[d_cache.scala 105:18 50:31]
  wire [63:0] _GEN_4211 = 4'h3 == state ? _GEN_666 : receive_data_6; // @[d_cache.scala 105:18 50:31]
  wire [63:0] _GEN_4212 = 4'h3 == state ? _GEN_667 : receive_data_7; // @[d_cache.scala 105:18 50:31]
  wire [2:0] _GEN_4213 = 4'h3 == state ? _GEN_668 : receive_num; // @[d_cache.scala 105:18 51:30]
  wire [3:0] _GEN_4214 = 4'h3 == state ? _GEN_669 : _GEN_3930; // @[d_cache.scala 105:18]
  wire [511:0] _GEN_4215 = 4'h3 == state ? ram_0_0 : _GEN_3931; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4216 = 4'h3 == state ? ram_0_1 : _GEN_3932; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4217 = 4'h3 == state ? ram_0_2 : _GEN_3933; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4218 = 4'h3 == state ? ram_0_3 : _GEN_3934; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4219 = 4'h3 == state ? ram_0_4 : _GEN_3935; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4220 = 4'h3 == state ? ram_0_5 : _GEN_3936; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4221 = 4'h3 == state ? ram_0_6 : _GEN_3937; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4222 = 4'h3 == state ? ram_0_7 : _GEN_3938; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4223 = 4'h3 == state ? ram_0_8 : _GEN_3939; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4224 = 4'h3 == state ? ram_0_9 : _GEN_3940; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4225 = 4'h3 == state ? ram_0_10 : _GEN_3941; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4226 = 4'h3 == state ? ram_0_11 : _GEN_3942; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4227 = 4'h3 == state ? ram_0_12 : _GEN_3943; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4228 = 4'h3 == state ? ram_0_13 : _GEN_3944; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4229 = 4'h3 == state ? ram_0_14 : _GEN_3945; // @[d_cache.scala 105:18 19:24]
  wire [511:0] _GEN_4230 = 4'h3 == state ? ram_0_15 : _GEN_3946; // @[d_cache.scala 105:18 19:24]
  wire [31:0] _GEN_4231 = 4'h3 == state ? tag_0_0 : _GEN_3947; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4232 = 4'h3 == state ? tag_0_1 : _GEN_3948; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4233 = 4'h3 == state ? tag_0_2 : _GEN_3949; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4234 = 4'h3 == state ? tag_0_3 : _GEN_3950; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4235 = 4'h3 == state ? tag_0_4 : _GEN_3951; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4236 = 4'h3 == state ? tag_0_5 : _GEN_3952; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4237 = 4'h3 == state ? tag_0_6 : _GEN_3953; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4238 = 4'h3 == state ? tag_0_7 : _GEN_3954; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4239 = 4'h3 == state ? tag_0_8 : _GEN_3955; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4240 = 4'h3 == state ? tag_0_9 : _GEN_3956; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4241 = 4'h3 == state ? tag_0_10 : _GEN_3957; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4242 = 4'h3 == state ? tag_0_11 : _GEN_3958; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4243 = 4'h3 == state ? tag_0_12 : _GEN_3959; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4244 = 4'h3 == state ? tag_0_13 : _GEN_3960; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4245 = 4'h3 == state ? tag_0_14 : _GEN_3961; // @[d_cache.scala 105:18 24:24]
  wire [31:0] _GEN_4246 = 4'h3 == state ? tag_0_15 : _GEN_3962; // @[d_cache.scala 105:18 24:24]
  wire  _GEN_4247 = 4'h3 == state ? valid_0_0 : _GEN_3963; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4248 = 4'h3 == state ? valid_0_1 : _GEN_3964; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4249 = 4'h3 == state ? valid_0_2 : _GEN_3965; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4250 = 4'h3 == state ? valid_0_3 : _GEN_3966; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4251 = 4'h3 == state ? valid_0_4 : _GEN_3967; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4252 = 4'h3 == state ? valid_0_5 : _GEN_3968; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4253 = 4'h3 == state ? valid_0_6 : _GEN_3969; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4254 = 4'h3 == state ? valid_0_7 : _GEN_3970; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4255 = 4'h3 == state ? valid_0_8 : _GEN_3971; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4256 = 4'h3 == state ? valid_0_9 : _GEN_3972; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4257 = 4'h3 == state ? valid_0_10 : _GEN_3973; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4258 = 4'h3 == state ? valid_0_11 : _GEN_3974; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4259 = 4'h3 == state ? valid_0_12 : _GEN_3975; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4260 = 4'h3 == state ? valid_0_13 : _GEN_3976; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4261 = 4'h3 == state ? valid_0_14 : _GEN_3977; // @[d_cache.scala 105:18 29:26]
  wire  _GEN_4262 = 4'h3 == state ? valid_0_15 : _GEN_3978; // @[d_cache.scala 105:18 29:26]
  wire [7:0] _GEN_4263 = 4'h3 == state ? quene_0 : _GEN_3979; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4264 = 4'h3 == state ? quene_1 : _GEN_3980; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4265 = 4'h3 == state ? quene_2 : _GEN_3981; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4266 = 4'h3 == state ? quene_3 : _GEN_3982; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4267 = 4'h3 == state ? quene_4 : _GEN_3983; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4268 = 4'h3 == state ? quene_5 : _GEN_3984; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4269 = 4'h3 == state ? quene_6 : _GEN_3985; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4270 = 4'h3 == state ? quene_7 : _GEN_3986; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4271 = 4'h3 == state ? quene_8 : _GEN_3987; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4272 = 4'h3 == state ? quene_9 : _GEN_3988; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4273 = 4'h3 == state ? quene_10 : _GEN_3989; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4274 = 4'h3 == state ? quene_11 : _GEN_3990; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4275 = 4'h3 == state ? quene_12 : _GEN_3991; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4276 = 4'h3 == state ? quene_13 : _GEN_3992; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4277 = 4'h3 == state ? quene_14 : _GEN_3993; // @[d_cache.scala 105:18 52:24]
  wire [7:0] _GEN_4278 = 4'h3 == state ? quene_15 : _GEN_3994; // @[d_cache.scala 105:18 52:24]
  wire [511:0] _GEN_4279 = 4'h3 == state ? ram_1_0 : _GEN_3995; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4280 = 4'h3 == state ? ram_1_1 : _GEN_3996; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4281 = 4'h3 == state ? ram_1_2 : _GEN_3997; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4282 = 4'h3 == state ? ram_1_3 : _GEN_3998; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4283 = 4'h3 == state ? ram_1_4 : _GEN_3999; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4284 = 4'h3 == state ? ram_1_5 : _GEN_4000; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4285 = 4'h3 == state ? ram_1_6 : _GEN_4001; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4286 = 4'h3 == state ? ram_1_7 : _GEN_4002; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4287 = 4'h3 == state ? ram_1_8 : _GEN_4003; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4288 = 4'h3 == state ? ram_1_9 : _GEN_4004; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4289 = 4'h3 == state ? ram_1_10 : _GEN_4005; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4290 = 4'h3 == state ? ram_1_11 : _GEN_4006; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4291 = 4'h3 == state ? ram_1_12 : _GEN_4007; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4292 = 4'h3 == state ? ram_1_13 : _GEN_4008; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4293 = 4'h3 == state ? ram_1_14 : _GEN_4009; // @[d_cache.scala 105:18 20:24]
  wire [511:0] _GEN_4294 = 4'h3 == state ? ram_1_15 : _GEN_4010; // @[d_cache.scala 105:18 20:24]
  wire [31:0] _GEN_4295 = 4'h3 == state ? tag_1_0 : _GEN_4011; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4296 = 4'h3 == state ? tag_1_1 : _GEN_4012; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4297 = 4'h3 == state ? tag_1_2 : _GEN_4013; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4298 = 4'h3 == state ? tag_1_3 : _GEN_4014; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4299 = 4'h3 == state ? tag_1_4 : _GEN_4015; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4300 = 4'h3 == state ? tag_1_5 : _GEN_4016; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4301 = 4'h3 == state ? tag_1_6 : _GEN_4017; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4302 = 4'h3 == state ? tag_1_7 : _GEN_4018; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4303 = 4'h3 == state ? tag_1_8 : _GEN_4019; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4304 = 4'h3 == state ? tag_1_9 : _GEN_4020; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4305 = 4'h3 == state ? tag_1_10 : _GEN_4021; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4306 = 4'h3 == state ? tag_1_11 : _GEN_4022; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4307 = 4'h3 == state ? tag_1_12 : _GEN_4023; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4308 = 4'h3 == state ? tag_1_13 : _GEN_4024; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4309 = 4'h3 == state ? tag_1_14 : _GEN_4025; // @[d_cache.scala 105:18 25:24]
  wire [31:0] _GEN_4310 = 4'h3 == state ? tag_1_15 : _GEN_4026; // @[d_cache.scala 105:18 25:24]
  wire  _GEN_4311 = 4'h3 == state ? valid_1_0 : _GEN_4027; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4312 = 4'h3 == state ? valid_1_1 : _GEN_4028; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4313 = 4'h3 == state ? valid_1_2 : _GEN_4029; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4314 = 4'h3 == state ? valid_1_3 : _GEN_4030; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4315 = 4'h3 == state ? valid_1_4 : _GEN_4031; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4316 = 4'h3 == state ? valid_1_5 : _GEN_4032; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4317 = 4'h3 == state ? valid_1_6 : _GEN_4033; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4318 = 4'h3 == state ? valid_1_7 : _GEN_4034; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4319 = 4'h3 == state ? valid_1_8 : _GEN_4035; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4320 = 4'h3 == state ? valid_1_9 : _GEN_4036; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4321 = 4'h3 == state ? valid_1_10 : _GEN_4037; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4322 = 4'h3 == state ? valid_1_11 : _GEN_4038; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4323 = 4'h3 == state ? valid_1_12 : _GEN_4039; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4324 = 4'h3 == state ? valid_1_13 : _GEN_4040; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4325 = 4'h3 == state ? valid_1_14 : _GEN_4041; // @[d_cache.scala 105:18 30:26]
  wire  _GEN_4326 = 4'h3 == state ? valid_1_15 : _GEN_4042; // @[d_cache.scala 105:18 30:26]
  wire [511:0] _GEN_4327 = 4'h3 == state ? ram_2_0 : _GEN_4043; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4328 = 4'h3 == state ? ram_2_1 : _GEN_4044; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4329 = 4'h3 == state ? ram_2_2 : _GEN_4045; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4330 = 4'h3 == state ? ram_2_3 : _GEN_4046; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4331 = 4'h3 == state ? ram_2_4 : _GEN_4047; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4332 = 4'h3 == state ? ram_2_5 : _GEN_4048; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4333 = 4'h3 == state ? ram_2_6 : _GEN_4049; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4334 = 4'h3 == state ? ram_2_7 : _GEN_4050; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4335 = 4'h3 == state ? ram_2_8 : _GEN_4051; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4336 = 4'h3 == state ? ram_2_9 : _GEN_4052; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4337 = 4'h3 == state ? ram_2_10 : _GEN_4053; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4338 = 4'h3 == state ? ram_2_11 : _GEN_4054; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4339 = 4'h3 == state ? ram_2_12 : _GEN_4055; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4340 = 4'h3 == state ? ram_2_13 : _GEN_4056; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4341 = 4'h3 == state ? ram_2_14 : _GEN_4057; // @[d_cache.scala 105:18 21:24]
  wire [511:0] _GEN_4342 = 4'h3 == state ? ram_2_15 : _GEN_4058; // @[d_cache.scala 105:18 21:24]
  wire [31:0] _GEN_4343 = 4'h3 == state ? tag_2_0 : _GEN_4059; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4344 = 4'h3 == state ? tag_2_1 : _GEN_4060; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4345 = 4'h3 == state ? tag_2_2 : _GEN_4061; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4346 = 4'h3 == state ? tag_2_3 : _GEN_4062; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4347 = 4'h3 == state ? tag_2_4 : _GEN_4063; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4348 = 4'h3 == state ? tag_2_5 : _GEN_4064; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4349 = 4'h3 == state ? tag_2_6 : _GEN_4065; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4350 = 4'h3 == state ? tag_2_7 : _GEN_4066; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4351 = 4'h3 == state ? tag_2_8 : _GEN_4067; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4352 = 4'h3 == state ? tag_2_9 : _GEN_4068; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4353 = 4'h3 == state ? tag_2_10 : _GEN_4069; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4354 = 4'h3 == state ? tag_2_11 : _GEN_4070; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4355 = 4'h3 == state ? tag_2_12 : _GEN_4071; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4356 = 4'h3 == state ? tag_2_13 : _GEN_4072; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4357 = 4'h3 == state ? tag_2_14 : _GEN_4073; // @[d_cache.scala 105:18 26:24]
  wire [31:0] _GEN_4358 = 4'h3 == state ? tag_2_15 : _GEN_4074; // @[d_cache.scala 105:18 26:24]
  wire  _GEN_4359 = 4'h3 == state ? valid_2_0 : _GEN_4075; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4360 = 4'h3 == state ? valid_2_1 : _GEN_4076; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4361 = 4'h3 == state ? valid_2_2 : _GEN_4077; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4362 = 4'h3 == state ? valid_2_3 : _GEN_4078; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4363 = 4'h3 == state ? valid_2_4 : _GEN_4079; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4364 = 4'h3 == state ? valid_2_5 : _GEN_4080; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4365 = 4'h3 == state ? valid_2_6 : _GEN_4081; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4366 = 4'h3 == state ? valid_2_7 : _GEN_4082; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4367 = 4'h3 == state ? valid_2_8 : _GEN_4083; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4368 = 4'h3 == state ? valid_2_9 : _GEN_4084; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4369 = 4'h3 == state ? valid_2_10 : _GEN_4085; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4370 = 4'h3 == state ? valid_2_11 : _GEN_4086; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4371 = 4'h3 == state ? valid_2_12 : _GEN_4087; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4372 = 4'h3 == state ? valid_2_13 : _GEN_4088; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4373 = 4'h3 == state ? valid_2_14 : _GEN_4089; // @[d_cache.scala 105:18 31:26]
  wire  _GEN_4374 = 4'h3 == state ? valid_2_15 : _GEN_4090; // @[d_cache.scala 105:18 31:26]
  wire [511:0] _GEN_4375 = 4'h3 == state ? ram_3_0 : _GEN_4091; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4376 = 4'h3 == state ? ram_3_1 : _GEN_4092; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4377 = 4'h3 == state ? ram_3_2 : _GEN_4093; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4378 = 4'h3 == state ? ram_3_3 : _GEN_4094; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4379 = 4'h3 == state ? ram_3_4 : _GEN_4095; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4380 = 4'h3 == state ? ram_3_5 : _GEN_4096; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4381 = 4'h3 == state ? ram_3_6 : _GEN_4097; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4382 = 4'h3 == state ? ram_3_7 : _GEN_4098; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4383 = 4'h3 == state ? ram_3_8 : _GEN_4099; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4384 = 4'h3 == state ? ram_3_9 : _GEN_4100; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4385 = 4'h3 == state ? ram_3_10 : _GEN_4101; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4386 = 4'h3 == state ? ram_3_11 : _GEN_4102; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4387 = 4'h3 == state ? ram_3_12 : _GEN_4103; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4388 = 4'h3 == state ? ram_3_13 : _GEN_4104; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4389 = 4'h3 == state ? ram_3_14 : _GEN_4105; // @[d_cache.scala 105:18 22:24]
  wire [511:0] _GEN_4390 = 4'h3 == state ? ram_3_15 : _GEN_4106; // @[d_cache.scala 105:18 22:24]
  wire [31:0] _GEN_4391 = 4'h3 == state ? tag_3_0 : _GEN_4107; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4392 = 4'h3 == state ? tag_3_1 : _GEN_4108; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4393 = 4'h3 == state ? tag_3_2 : _GEN_4109; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4394 = 4'h3 == state ? tag_3_3 : _GEN_4110; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4395 = 4'h3 == state ? tag_3_4 : _GEN_4111; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4396 = 4'h3 == state ? tag_3_5 : _GEN_4112; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4397 = 4'h3 == state ? tag_3_6 : _GEN_4113; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4398 = 4'h3 == state ? tag_3_7 : _GEN_4114; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4399 = 4'h3 == state ? tag_3_8 : _GEN_4115; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4400 = 4'h3 == state ? tag_3_9 : _GEN_4116; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4401 = 4'h3 == state ? tag_3_10 : _GEN_4117; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4402 = 4'h3 == state ? tag_3_11 : _GEN_4118; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4403 = 4'h3 == state ? tag_3_12 : _GEN_4119; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4404 = 4'h3 == state ? tag_3_13 : _GEN_4120; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4405 = 4'h3 == state ? tag_3_14 : _GEN_4121; // @[d_cache.scala 105:18 27:24]
  wire [31:0] _GEN_4406 = 4'h3 == state ? tag_3_15 : _GEN_4122; // @[d_cache.scala 105:18 27:24]
  wire  _GEN_4407 = 4'h3 == state ? valid_3_0 : _GEN_4123; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4408 = 4'h3 == state ? valid_3_1 : _GEN_4124; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4409 = 4'h3 == state ? valid_3_2 : _GEN_4125; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4410 = 4'h3 == state ? valid_3_3 : _GEN_4126; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4411 = 4'h3 == state ? valid_3_4 : _GEN_4127; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4412 = 4'h3 == state ? valid_3_5 : _GEN_4128; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4413 = 4'h3 == state ? valid_3_6 : _GEN_4129; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4414 = 4'h3 == state ? valid_3_7 : _GEN_4130; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4415 = 4'h3 == state ? valid_3_8 : _GEN_4131; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4416 = 4'h3 == state ? valid_3_9 : _GEN_4132; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4417 = 4'h3 == state ? valid_3_10 : _GEN_4133; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4418 = 4'h3 == state ? valid_3_11 : _GEN_4134; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4419 = 4'h3 == state ? valid_3_12 : _GEN_4135; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4420 = 4'h3 == state ? valid_3_13 : _GEN_4136; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4421 = 4'h3 == state ? valid_3_14 : _GEN_4137; // @[d_cache.scala 105:18 32:26]
  wire  _GEN_4422 = 4'h3 == state ? valid_3_15 : _GEN_4138; // @[d_cache.scala 105:18 32:26]
  wire [511:0] _GEN_4423 = 4'h3 == state ? write_back_data : _GEN_4139; // @[d_cache.scala 105:18 44:34]
  wire [41:0] _GEN_4424 = 4'h3 == state ? {{10'd0}, write_back_addr} : _GEN_4140; // @[d_cache.scala 105:18 45:34]
  wire  _GEN_4425 = 4'h3 == state ? dirty_0_0 : _GEN_4141; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4426 = 4'h3 == state ? dirty_0_1 : _GEN_4142; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4427 = 4'h3 == state ? dirty_0_2 : _GEN_4143; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4428 = 4'h3 == state ? dirty_0_3 : _GEN_4144; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4429 = 4'h3 == state ? dirty_0_4 : _GEN_4145; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4430 = 4'h3 == state ? dirty_0_5 : _GEN_4146; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4431 = 4'h3 == state ? dirty_0_6 : _GEN_4147; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4432 = 4'h3 == state ? dirty_0_7 : _GEN_4148; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4433 = 4'h3 == state ? dirty_0_8 : _GEN_4149; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4434 = 4'h3 == state ? dirty_0_9 : _GEN_4150; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4435 = 4'h3 == state ? dirty_0_10 : _GEN_4151; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4436 = 4'h3 == state ? dirty_0_11 : _GEN_4152; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4437 = 4'h3 == state ? dirty_0_12 : _GEN_4153; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4438 = 4'h3 == state ? dirty_0_13 : _GEN_4154; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4439 = 4'h3 == state ? dirty_0_14 : _GEN_4155; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4440 = 4'h3 == state ? dirty_0_15 : _GEN_4156; // @[d_cache.scala 105:18 34:26]
  wire  _GEN_4441 = 4'h3 == state ? dirty_1_0 : _GEN_4157; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4442 = 4'h3 == state ? dirty_1_1 : _GEN_4158; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4443 = 4'h3 == state ? dirty_1_2 : _GEN_4159; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4444 = 4'h3 == state ? dirty_1_3 : _GEN_4160; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4445 = 4'h3 == state ? dirty_1_4 : _GEN_4161; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4446 = 4'h3 == state ? dirty_1_5 : _GEN_4162; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4447 = 4'h3 == state ? dirty_1_6 : _GEN_4163; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4448 = 4'h3 == state ? dirty_1_7 : _GEN_4164; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4449 = 4'h3 == state ? dirty_1_8 : _GEN_4165; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4450 = 4'h3 == state ? dirty_1_9 : _GEN_4166; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4451 = 4'h3 == state ? dirty_1_10 : _GEN_4167; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4452 = 4'h3 == state ? dirty_1_11 : _GEN_4168; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4453 = 4'h3 == state ? dirty_1_12 : _GEN_4169; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4454 = 4'h3 == state ? dirty_1_13 : _GEN_4170; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4455 = 4'h3 == state ? dirty_1_14 : _GEN_4171; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4456 = 4'h3 == state ? dirty_1_15 : _GEN_4172; // @[d_cache.scala 105:18 35:26]
  wire  _GEN_4457 = 4'h3 == state ? dirty_2_0 : _GEN_4173; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4458 = 4'h3 == state ? dirty_2_1 : _GEN_4174; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4459 = 4'h3 == state ? dirty_2_2 : _GEN_4175; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4460 = 4'h3 == state ? dirty_2_3 : _GEN_4176; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4461 = 4'h3 == state ? dirty_2_4 : _GEN_4177; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4462 = 4'h3 == state ? dirty_2_5 : _GEN_4178; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4463 = 4'h3 == state ? dirty_2_6 : _GEN_4179; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4464 = 4'h3 == state ? dirty_2_7 : _GEN_4180; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4465 = 4'h3 == state ? dirty_2_8 : _GEN_4181; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4466 = 4'h3 == state ? dirty_2_9 : _GEN_4182; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4467 = 4'h3 == state ? dirty_2_10 : _GEN_4183; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4468 = 4'h3 == state ? dirty_2_11 : _GEN_4184; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4469 = 4'h3 == state ? dirty_2_12 : _GEN_4185; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4470 = 4'h3 == state ? dirty_2_13 : _GEN_4186; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4471 = 4'h3 == state ? dirty_2_14 : _GEN_4187; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4472 = 4'h3 == state ? dirty_2_15 : _GEN_4188; // @[d_cache.scala 105:18 36:26]
  wire  _GEN_4473 = 4'h3 == state ? dirty_3_0 : _GEN_4189; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4474 = 4'h3 == state ? dirty_3_1 : _GEN_4190; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4475 = 4'h3 == state ? dirty_3_2 : _GEN_4191; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4476 = 4'h3 == state ? dirty_3_3 : _GEN_4192; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4477 = 4'h3 == state ? dirty_3_4 : _GEN_4193; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4478 = 4'h3 == state ? dirty_3_5 : _GEN_4194; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4479 = 4'h3 == state ? dirty_3_6 : _GEN_4195; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4480 = 4'h3 == state ? dirty_3_7 : _GEN_4196; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4481 = 4'h3 == state ? dirty_3_8 : _GEN_4197; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4482 = 4'h3 == state ? dirty_3_9 : _GEN_4198; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4483 = 4'h3 == state ? dirty_3_10 : _GEN_4199; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4484 = 4'h3 == state ? dirty_3_11 : _GEN_4200; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4485 = 4'h3 == state ? dirty_3_12 : _GEN_4201; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4486 = 4'h3 == state ? dirty_3_13 : _GEN_4202; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4487 = 4'h3 == state ? dirty_3_14 : _GEN_4203; // @[d_cache.scala 105:18 37:26]
  wire  _GEN_4488 = 4'h3 == state ? dirty_3_15 : _GEN_4204; // @[d_cache.scala 105:18 37:26]
  wire [41:0] _GEN_4772 = 4'h2 == state ? {{10'd0}, write_back_addr} : _GEN_4424; // @[d_cache.scala 105:18 45:34]
  wire [41:0] _GEN_5056 = 4'h1 == state ? {{10'd0}, write_back_addr} : _GEN_4772; // @[d_cache.scala 105:18 45:34]
  wire [41:0] _GEN_5340 = 4'h0 == state ? {{10'd0}, write_back_addr} : _GEN_5056; // @[d_cache.scala 105:18 45:34]
  wire [511:0] _io_to_lsu_rdata_T = _GEN_150 >> shift_bit; // @[d_cache.scala 316:56]
  wire [511:0] _io_to_lsu_rdata_T_1 = _GEN_198 >> shift_bit; // @[d_cache.scala 316:98]
  wire [511:0] _io_to_lsu_rdata_T_2 = _GEN_246 >> shift_bit; // @[d_cache.scala 316:140]
  wire [511:0] _io_to_lsu_rdata_T_3 = _GEN_294 >> shift_bit; // @[d_cache.scala 316:169]
  wire [511:0] _io_to_lsu_rdata_T_4 = way2_hit ? _io_to_lsu_rdata_T_2 : _io_to_lsu_rdata_T_3; // @[d_cache.scala 316:116]
  wire [511:0] _io_to_lsu_rdata_T_5 = way1_hit ? _io_to_lsu_rdata_T_1 : _io_to_lsu_rdata_T_4; // @[d_cache.scala 316:74]
  wire [511:0] _io_to_lsu_rdata_T_6 = way0_hit ? _io_to_lsu_rdata_T : _io_to_lsu_rdata_T_5; // @[d_cache.scala 316:32]
  wire [63:0] _GEN_5702 = {{32'd0}, io_from_lsu_araddr}; // @[d_cache.scala 358:49]
  wire [63:0] _io_to_axi_araddr_T = _GEN_5702 & 64'hffffffffffffffc0; // @[d_cache.scala 358:49]
  wire  _T_35 = state == 4'h7; // @[d_cache.scala 438:21]
  wire [63:0] _GEN_5342 = state == 4'h7 ? io_from_axi_rdata : 64'h0; // @[d_cache.scala 438:30 439:19 442:25]
  wire  _GEN_5344 = state == 4'h7 & io_from_axi_rvalid; // @[d_cache.scala 438:30 439:19 444:26]
  wire  _GEN_5346 = state == 4'h7 & io_from_axi_wready; // @[d_cache.scala 438:30 439:19 446:26]
  wire  _GEN_5352 = state == 4'h7 & io_from_lsu_arvalid; // @[d_cache.scala 438:30 440:19 449:27]
  wire [31:0] _GEN_5354 = state == 4'h7 ? io_from_lsu_awaddr : 32'h0; // @[d_cache.scala 438:30 440:19 455:26]
  wire  _GEN_5358 = state == 4'h7 & io_from_lsu_awvalid; // @[d_cache.scala 438:30 440:19 456:27]
  wire [63:0] _GEN_5359 = state == 4'h7 ? io_from_lsu_wdata : 64'h0; // @[d_cache.scala 438:30 440:19 460:25]
  wire [7:0] _GEN_5360 = state == 4'h7 ? io_from_lsu_wstrb : 8'h0; // @[d_cache.scala 438:30 440:19 461:25]
  wire  _GEN_5362 = state == 4'h7 & io_from_lsu_wvalid; // @[d_cache.scala 438:30 440:19 463:26]
  wire [63:0] _GEN_5364 = state == 4'h6 ? 64'h0 : _GEN_5342; // @[d_cache.scala 414:35 415:25]
  wire  _GEN_5366 = state == 4'h6 ? 1'h0 : _GEN_5344; // @[d_cache.scala 414:35 417:26]
  wire  _GEN_5368 = state == 4'h6 ? 1'h0 : _GEN_5346; // @[d_cache.scala 414:35 419:26]
  wire  _GEN_5371 = state == 4'h6 ? 1'h0 : _GEN_5352; // @[d_cache.scala 414:35 422:27]
  wire [31:0] _GEN_5372 = state == 4'h6 ? 32'h0 : io_from_lsu_araddr; // @[d_cache.scala 414:35 423:26]
  wire [7:0] _GEN_5373 = state == 4'h6 ? 8'h7 : 8'h0; // @[d_cache.scala 414:35 424:25]
  wire  _GEN_5376 = state == 4'h6 ? 1'h0 : 1'h1; // @[d_cache.scala 414:35 427:26]
  wire [31:0] _GEN_5377 = state == 4'h6 ? write_back_addr : _GEN_5354; // @[d_cache.scala 414:35 428:26]
  wire  _GEN_5378 = state == 4'h6 | _GEN_5358; // @[d_cache.scala 414:35 429:27]
  wire [63:0] _GEN_5382 = state == 4'h6 ? write_back_data[63:0] : _GEN_5359; // @[d_cache.scala 414:35 433:25]
  wire [7:0] _GEN_5383 = state == 4'h6 ? 8'hff : _GEN_5360; // @[d_cache.scala 414:35 434:25]
  wire  _GEN_5385 = state == 4'h6 | _GEN_5362; // @[d_cache.scala 414:35 436:26]
  wire  _GEN_5386 = state == 4'h6 | _T_35; // @[d_cache.scala 414:35 437:26]
  wire [63:0] _GEN_5387 = state == 4'h4 | state == 4'h8 ? 64'h0 : _GEN_5364; // @[d_cache.scala 373:50 374:25]
  wire  _GEN_5389 = state == 4'h4 | state == 4'h8 ? 1'h0 : _GEN_5366; // @[d_cache.scala 373:50 376:26]
  wire  _GEN_5391 = state == 4'h4 | state == 4'h8 ? io_from_axi_wready : _GEN_5368; // @[d_cache.scala 373:50 378:26]
  wire  _GEN_5394 = state == 4'h4 | state == 4'h8 ? 1'h0 : _GEN_5371; // @[d_cache.scala 373:50 381:27]
  wire [31:0] _GEN_5395 = state == 4'h4 | state == 4'h8 ? 32'h0 : _GEN_5372; // @[d_cache.scala 373:50 382:26]
  wire [7:0] _GEN_5396 = state == 4'h4 | state == 4'h8 ? 8'h0 : _GEN_5373; // @[d_cache.scala 373:50 383:25]
  wire  _GEN_5399 = state == 4'h4 | state == 4'h8 | _GEN_5376; // @[d_cache.scala 373:50 386:26]
  wire [31:0] _GEN_5400 = state == 4'h4 | state == 4'h8 ? io_from_lsu_awaddr : _GEN_5377; // @[d_cache.scala 373:50 387:26]
  wire  _GEN_5401 = state == 4'h4 | state == 4'h8 ? io_from_lsu_awvalid : _GEN_5378; // @[d_cache.scala 373:50 388:27]
  wire [63:0] _GEN_5405 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wdata : _GEN_5382; // @[d_cache.scala 373:50 392:25]
  wire [7:0] _GEN_5406 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wstrb : _GEN_5383; // @[d_cache.scala 373:50 393:25]
  wire  _GEN_5408 = state == 4'h4 | state == 4'h8 ? io_from_lsu_wvalid : _GEN_5385; // @[d_cache.scala 373:50 395:26]
  wire  _GEN_5409 = state == 4'h4 | state == 4'h8 | _GEN_5386; // @[d_cache.scala 373:50 396:26]
  wire [63:0] _GEN_5410 = state == 4'h3 ? 64'h0 : _GEN_5387; // @[d_cache.scala 349:31 350:25]
  wire  _GEN_5412 = state == 4'h3 ? 1'h0 : _GEN_5389; // @[d_cache.scala 349:31 352:26]
  wire  _GEN_5414 = state == 4'h3 ? 1'h0 : _GEN_5391; // @[d_cache.scala 349:31 354:26]
  wire  _GEN_5417 = state == 4'h3 | _GEN_5394; // @[d_cache.scala 349:31 357:27]
  wire [63:0] _GEN_5418 = state == 4'h3 ? _io_to_axi_araddr_T : {{32'd0}, _GEN_5395}; // @[d_cache.scala 349:31 358:26]
  wire [7:0] _GEN_5419 = state == 4'h3 ? 8'h7 : _GEN_5396; // @[d_cache.scala 349:31 359:25]
  wire  _GEN_5422 = state == 4'h3 | _GEN_5399; // @[d_cache.scala 349:31 362:26]
  wire [31:0] _GEN_5423 = state == 4'h3 ? 32'h0 : _GEN_5400; // @[d_cache.scala 349:31 363:26]
  wire  _GEN_5424 = state == 4'h3 ? 1'h0 : _GEN_5401; // @[d_cache.scala 349:31 364:27]
  wire [7:0] _GEN_5425 = state == 4'h3 ? 8'h0 : _GEN_5396; // @[d_cache.scala 349:31 365:25]
  wire [63:0] _GEN_5428 = state == 4'h3 ? 64'h0 : _GEN_5405; // @[d_cache.scala 349:31 368:25]
  wire [7:0] _GEN_5429 = state == 4'h3 ? 8'h0 : _GEN_5406; // @[d_cache.scala 349:31 369:25]
  wire  _GEN_5431 = state == 4'h3 ? 1'h0 : _GEN_5408; // @[d_cache.scala 349:31 371:26]
  wire  _GEN_5432 = state == 4'h3 ? 1'h0 : _GEN_5409; // @[d_cache.scala 349:31 372:26]
  wire  _GEN_5433 = state == 4'h2 ? 1'h0 : _GEN_5417; // @[d_cache.scala 323:33 324:27]
  wire [63:0] _GEN_5434 = state == 4'h2 ? {{32'd0}, io_from_lsu_araddr} : _GEN_5418; // @[d_cache.scala 323:33 325:26]
  wire [7:0] _GEN_5435 = state == 4'h2 ? 8'h0 : _GEN_5419; // @[d_cache.scala 323:33 326:25]
  wire  _GEN_5438 = state == 4'h2 ? 1'h0 : _GEN_5422; // @[d_cache.scala 323:33 329:26]
  wire [31:0] _GEN_5439 = state == 4'h2 ? 32'h0 : _GEN_5423; // @[d_cache.scala 323:33 330:26]
  wire  _GEN_5440 = state == 4'h2 ? 1'h0 : _GEN_5424; // @[d_cache.scala 323:33 331:27]
  wire [7:0] _GEN_5441 = state == 4'h2 ? 8'h0 : _GEN_5425; // @[d_cache.scala 323:33 332:25]
  wire [63:0] _GEN_5444 = state == 4'h2 ? 64'h0 : _GEN_5428; // @[d_cache.scala 323:33 335:25]
  wire [7:0] _GEN_5445 = state == 4'h2 ? 8'h0 : _GEN_5429; // @[d_cache.scala 323:33 336:25]
  wire  _GEN_5447 = state == 4'h2 ? 1'h0 : _GEN_5431; // @[d_cache.scala 323:33 338:26]
  wire  _GEN_5448 = state == 4'h2 ? 1'h0 : _GEN_5432; // @[d_cache.scala 323:33 339:26]
  wire [63:0] _GEN_5449 = state == 4'h2 ? 64'h0 : _GEN_5410; // @[d_cache.scala 323:33 341:25]
  wire  _GEN_5451 = state == 4'h2 ? 1'h0 : _GEN_5412; // @[d_cache.scala 323:33 343:26]
  wire  _GEN_5453 = state == 4'h2 ? _T_6 : _GEN_5414; // @[d_cache.scala 323:33 345:26]
  wire [63:0] _GEN_5457 = state == 4'h1 ? {{32'd0}, io_from_lsu_araddr} : _GEN_5434; // @[d_cache.scala 299:27 301:26]
  wire [511:0] _GEN_5472 = state == 4'h1 ? _io_to_lsu_rdata_T_6 : {{448'd0}, _GEN_5449}; // @[d_cache.scala 299:27 316:25]
  wire [41:0] _GEN_5703 = reset ? 42'h0 : _GEN_5340; // @[d_cache.scala 45:{34,34}]
  assign io_to_lsu_rdata = _GEN_5472[63:0];
  assign io_to_lsu_rvalid = state == 4'h1 ? _T_6 : _GEN_5451; // @[d_cache.scala 299:27 318:26]
  assign io_to_lsu_wready = state == 4'h1 ? 1'h0 : _GEN_5453; // @[d_cache.scala 299:27 320:26]
  assign io_to_axi_araddr = _GEN_5457[31:0];
  assign io_to_axi_arlen = state == 4'h1 ? 8'h0 : _GEN_5435; // @[d_cache.scala 299:27 302:25]
  assign io_to_axi_arvalid = state == 4'h1 ? 1'h0 : _GEN_5433; // @[d_cache.scala 299:27 300:27]
  assign io_to_axi_rready = state == 4'h1 ? 1'h0 : _GEN_5438; // @[d_cache.scala 299:27 305:26]
  assign io_to_axi_awaddr = state == 4'h1 ? 32'h0 : _GEN_5439; // @[d_cache.scala 299:27 306:26]
  assign io_to_axi_awlen = state == 4'h1 ? 8'h0 : _GEN_5441; // @[d_cache.scala 299:27 308:25]
  assign io_to_axi_awvalid = state == 4'h1 ? 1'h0 : _GEN_5440; // @[d_cache.scala 299:27 307:27]
  assign io_to_axi_wdata = state == 4'h1 ? 64'h0 : _GEN_5444; // @[d_cache.scala 299:27 311:25]
  assign io_to_axi_wstrb = state == 4'h1 ? 8'h0 : _GEN_5445; // @[d_cache.scala 299:27 312:25]
  assign io_to_axi_wvalid = state == 4'h1 ? 1'h0 : _GEN_5447; // @[d_cache.scala 299:27 314:26]
  assign io_to_axi_bready = state == 4'h1 ? 1'h0 : _GEN_5448; // @[d_cache.scala 299:27 315:26]
  always @(posedge clock) begin
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_0 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_0 <= _GEN_523;
        end else begin
          ram_0_0 <= _GEN_4215;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_1 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_1 <= _GEN_524;
        end else begin
          ram_0_1 <= _GEN_4216;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_2 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_2 <= _GEN_525;
        end else begin
          ram_0_2 <= _GEN_4217;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_3 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_3 <= _GEN_526;
        end else begin
          ram_0_3 <= _GEN_4218;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_4 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_4 <= _GEN_527;
        end else begin
          ram_0_4 <= _GEN_4219;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_5 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_5 <= _GEN_528;
        end else begin
          ram_0_5 <= _GEN_4220;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_6 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_6 <= _GEN_529;
        end else begin
          ram_0_6 <= _GEN_4221;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_7 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_7 <= _GEN_530;
        end else begin
          ram_0_7 <= _GEN_4222;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_8 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_8 <= _GEN_531;
        end else begin
          ram_0_8 <= _GEN_4223;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_9 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_9 <= _GEN_532;
        end else begin
          ram_0_9 <= _GEN_4224;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_10 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_10 <= _GEN_533;
        end else begin
          ram_0_10 <= _GEN_4225;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_11 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_11 <= _GEN_534;
        end else begin
          ram_0_11 <= _GEN_4226;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_12 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_12 <= _GEN_535;
        end else begin
          ram_0_12 <= _GEN_4227;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_13 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_13 <= _GEN_536;
        end else begin
          ram_0_13 <= _GEN_4228;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_14 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_14 <= _GEN_537;
        end else begin
          ram_0_14 <= _GEN_4229;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 19:24]
      ram_0_15 <= 512'h0; // @[d_cache.scala 19:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_0_15 <= _GEN_538;
        end else begin
          ram_0_15 <= _GEN_4230;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_0 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_0 <= _GEN_555;
        end else begin
          ram_1_0 <= _GEN_4279;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_1 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_1 <= _GEN_556;
        end else begin
          ram_1_1 <= _GEN_4280;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_2 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_2 <= _GEN_557;
        end else begin
          ram_1_2 <= _GEN_4281;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_3 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_3 <= _GEN_558;
        end else begin
          ram_1_3 <= _GEN_4282;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_4 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_4 <= _GEN_559;
        end else begin
          ram_1_4 <= _GEN_4283;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_5 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_5 <= _GEN_560;
        end else begin
          ram_1_5 <= _GEN_4284;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_6 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_6 <= _GEN_561;
        end else begin
          ram_1_6 <= _GEN_4285;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_7 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_7 <= _GEN_562;
        end else begin
          ram_1_7 <= _GEN_4286;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_8 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_8 <= _GEN_563;
        end else begin
          ram_1_8 <= _GEN_4287;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_9 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_9 <= _GEN_564;
        end else begin
          ram_1_9 <= _GEN_4288;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_10 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_10 <= _GEN_565;
        end else begin
          ram_1_10 <= _GEN_4289;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_11 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_11 <= _GEN_566;
        end else begin
          ram_1_11 <= _GEN_4290;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_12 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_12 <= _GEN_567;
        end else begin
          ram_1_12 <= _GEN_4291;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_13 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_13 <= _GEN_568;
        end else begin
          ram_1_13 <= _GEN_4292;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_14 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_14 <= _GEN_569;
        end else begin
          ram_1_14 <= _GEN_4293;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 20:24]
      ram_1_15 <= 512'h0; // @[d_cache.scala 20:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_1_15 <= _GEN_570;
        end else begin
          ram_1_15 <= _GEN_4294;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_0 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_0 <= _GEN_587;
        end else begin
          ram_2_0 <= _GEN_4327;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_1 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_1 <= _GEN_588;
        end else begin
          ram_2_1 <= _GEN_4328;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_2 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_2 <= _GEN_589;
        end else begin
          ram_2_2 <= _GEN_4329;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_3 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_3 <= _GEN_590;
        end else begin
          ram_2_3 <= _GEN_4330;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_4 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_4 <= _GEN_591;
        end else begin
          ram_2_4 <= _GEN_4331;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_5 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_5 <= _GEN_592;
        end else begin
          ram_2_5 <= _GEN_4332;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_6 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_6 <= _GEN_593;
        end else begin
          ram_2_6 <= _GEN_4333;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_7 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_7 <= _GEN_594;
        end else begin
          ram_2_7 <= _GEN_4334;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_8 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_8 <= _GEN_595;
        end else begin
          ram_2_8 <= _GEN_4335;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_9 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_9 <= _GEN_596;
        end else begin
          ram_2_9 <= _GEN_4336;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_10 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_10 <= _GEN_597;
        end else begin
          ram_2_10 <= _GEN_4337;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_11 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_11 <= _GEN_598;
        end else begin
          ram_2_11 <= _GEN_4338;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_12 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_12 <= _GEN_599;
        end else begin
          ram_2_12 <= _GEN_4339;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_13 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_13 <= _GEN_600;
        end else begin
          ram_2_13 <= _GEN_4340;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_14 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_14 <= _GEN_601;
        end else begin
          ram_2_14 <= _GEN_4341;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 21:24]
      ram_2_15 <= 512'h0; // @[d_cache.scala 21:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_2_15 <= _GEN_602;
        end else begin
          ram_2_15 <= _GEN_4342;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_0 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_0 <= _GEN_619;
        end else begin
          ram_3_0 <= _GEN_4375;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_1 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_1 <= _GEN_620;
        end else begin
          ram_3_1 <= _GEN_4376;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_2 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_2 <= _GEN_621;
        end else begin
          ram_3_2 <= _GEN_4377;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_3 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_3 <= _GEN_622;
        end else begin
          ram_3_3 <= _GEN_4378;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_4 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_4 <= _GEN_623;
        end else begin
          ram_3_4 <= _GEN_4379;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_5 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_5 <= _GEN_624;
        end else begin
          ram_3_5 <= _GEN_4380;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_6 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_6 <= _GEN_625;
        end else begin
          ram_3_6 <= _GEN_4381;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_7 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_7 <= _GEN_626;
        end else begin
          ram_3_7 <= _GEN_4382;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_8 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_8 <= _GEN_627;
        end else begin
          ram_3_8 <= _GEN_4383;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_9 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_9 <= _GEN_628;
        end else begin
          ram_3_9 <= _GEN_4384;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_10 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_10 <= _GEN_629;
        end else begin
          ram_3_10 <= _GEN_4385;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_11 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_11 <= _GEN_630;
        end else begin
          ram_3_11 <= _GEN_4386;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_12 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_12 <= _GEN_631;
        end else begin
          ram_3_12 <= _GEN_4387;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_13 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_13 <= _GEN_632;
        end else begin
          ram_3_13 <= _GEN_4388;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_14 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_14 <= _GEN_633;
        end else begin
          ram_3_14 <= _GEN_4389;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 22:24]
      ram_3_15 <= 512'h0; // @[d_cache.scala 22:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          ram_3_15 <= _GEN_634;
        end else begin
          ram_3_15 <= _GEN_4390;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_0 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_0 <= _GEN_4231;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_1 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_1 <= _GEN_4232;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_2 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_2 <= _GEN_4233;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_3 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_3 <= _GEN_4234;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_4 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_4 <= _GEN_4235;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_5 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_5 <= _GEN_4236;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_6 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_6 <= _GEN_4237;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_7 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_7 <= _GEN_4238;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_8 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_8 <= _GEN_4239;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_9 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_9 <= _GEN_4240;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_10 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_10 <= _GEN_4241;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_11 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_11 <= _GEN_4242;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_12 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_12 <= _GEN_4243;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_13 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_13 <= _GEN_4244;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_14 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_14 <= _GEN_4245;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 24:24]
      tag_0_15 <= 32'h0; // @[d_cache.scala 24:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_0_15 <= _GEN_4246;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_0 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_0 <= _GEN_4295;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_1 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_1 <= _GEN_4296;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_2 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_2 <= _GEN_4297;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_3 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_3 <= _GEN_4298;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_4 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_4 <= _GEN_4299;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_5 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_5 <= _GEN_4300;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_6 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_6 <= _GEN_4301;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_7 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_7 <= _GEN_4302;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_8 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_8 <= _GEN_4303;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_9 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_9 <= _GEN_4304;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_10 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_10 <= _GEN_4305;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_11 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_11 <= _GEN_4306;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_12 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_12 <= _GEN_4307;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_13 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_13 <= _GEN_4308;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_14 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_14 <= _GEN_4309;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 25:24]
      tag_1_15 <= 32'h0; // @[d_cache.scala 25:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_1_15 <= _GEN_4310;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_0 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_0 <= _GEN_4343;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_1 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_1 <= _GEN_4344;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_2 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_2 <= _GEN_4345;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_3 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_3 <= _GEN_4346;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_4 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_4 <= _GEN_4347;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_5 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_5 <= _GEN_4348;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_6 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_6 <= _GEN_4349;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_7 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_7 <= _GEN_4350;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_8 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_8 <= _GEN_4351;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_9 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_9 <= _GEN_4352;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_10 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_10 <= _GEN_4353;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_11 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_11 <= _GEN_4354;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_12 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_12 <= _GEN_4355;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_13 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_13 <= _GEN_4356;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_14 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_14 <= _GEN_4357;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 26:24]
      tag_2_15 <= 32'h0; // @[d_cache.scala 26:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_2_15 <= _GEN_4358;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_0 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_0 <= _GEN_4391;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_1 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_1 <= _GEN_4392;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_2 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_2 <= _GEN_4393;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_3 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_3 <= _GEN_4394;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_4 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_4 <= _GEN_4395;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_5 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_5 <= _GEN_4396;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_6 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_6 <= _GEN_4397;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_7 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_7 <= _GEN_4398;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_8 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_8 <= _GEN_4399;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_9 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_9 <= _GEN_4400;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_10 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_10 <= _GEN_4401;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_11 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_11 <= _GEN_4402;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_12 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_12 <= _GEN_4403;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_13 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_13 <= _GEN_4404;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_14 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_14 <= _GEN_4405;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 27:24]
      tag_3_15 <= 32'h0; // @[d_cache.scala 27:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          tag_3_15 <= _GEN_4406;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_0 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_0 <= _GEN_4247;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_1 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_1 <= _GEN_4248;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_2 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_2 <= _GEN_4249;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_3 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_3 <= _GEN_4250;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_4 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_4 <= _GEN_4251;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_5 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_5 <= _GEN_4252;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_6 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_6 <= _GEN_4253;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_7 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_7 <= _GEN_4254;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_8 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_8 <= _GEN_4255;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_9 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_9 <= _GEN_4256;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_10 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_10 <= _GEN_4257;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_11 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_11 <= _GEN_4258;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_12 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_12 <= _GEN_4259;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_13 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_13 <= _GEN_4260;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_14 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_14 <= _GEN_4261;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 29:26]
      valid_0_15 <= 1'h0; // @[d_cache.scala 29:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_0_15 <= _GEN_4262;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_0 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_0 <= _GEN_4311;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_1 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_1 <= _GEN_4312;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_2 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_2 <= _GEN_4313;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_3 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_3 <= _GEN_4314;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_4 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_4 <= _GEN_4315;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_5 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_5 <= _GEN_4316;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_6 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_6 <= _GEN_4317;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_7 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_7 <= _GEN_4318;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_8 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_8 <= _GEN_4319;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_9 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_9 <= _GEN_4320;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_10 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_10 <= _GEN_4321;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_11 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_11 <= _GEN_4322;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_12 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_12 <= _GEN_4323;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_13 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_13 <= _GEN_4324;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_14 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_14 <= _GEN_4325;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 30:26]
      valid_1_15 <= 1'h0; // @[d_cache.scala 30:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_1_15 <= _GEN_4326;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_0 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_0 <= _GEN_4359;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_1 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_1 <= _GEN_4360;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_2 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_2 <= _GEN_4361;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_3 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_3 <= _GEN_4362;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_4 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_4 <= _GEN_4363;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_5 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_5 <= _GEN_4364;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_6 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_6 <= _GEN_4365;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_7 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_7 <= _GEN_4366;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_8 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_8 <= _GEN_4367;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_9 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_9 <= _GEN_4368;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_10 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_10 <= _GEN_4369;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_11 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_11 <= _GEN_4370;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_12 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_12 <= _GEN_4371;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_13 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_13 <= _GEN_4372;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_14 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_14 <= _GEN_4373;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 31:26]
      valid_2_15 <= 1'h0; // @[d_cache.scala 31:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_2_15 <= _GEN_4374;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_0 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_0 <= _GEN_4407;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_1 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_1 <= _GEN_4408;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_2 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_2 <= _GEN_4409;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_3 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_3 <= _GEN_4410;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_4 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_4 <= _GEN_4411;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_5 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_5 <= _GEN_4412;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_6 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_6 <= _GEN_4413;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_7 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_7 <= _GEN_4414;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_8 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_8 <= _GEN_4415;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_9 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_9 <= _GEN_4416;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_10 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_10 <= _GEN_4417;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_11 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_11 <= _GEN_4418;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_12 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_12 <= _GEN_4419;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_13 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_13 <= _GEN_4420;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_14 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_14 <= _GEN_4421;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 32:26]
      valid_3_15 <= 1'h0; // @[d_cache.scala 32:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          valid_3_15 <= _GEN_4422;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_0 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_0 <= _GEN_539;
        end else begin
          dirty_0_0 <= _GEN_4425;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_1 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_1 <= _GEN_540;
        end else begin
          dirty_0_1 <= _GEN_4426;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_2 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_2 <= _GEN_541;
        end else begin
          dirty_0_2 <= _GEN_4427;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_3 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_3 <= _GEN_542;
        end else begin
          dirty_0_3 <= _GEN_4428;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_4 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_4 <= _GEN_543;
        end else begin
          dirty_0_4 <= _GEN_4429;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_5 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_5 <= _GEN_544;
        end else begin
          dirty_0_5 <= _GEN_4430;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_6 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_6 <= _GEN_545;
        end else begin
          dirty_0_6 <= _GEN_4431;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_7 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_7 <= _GEN_546;
        end else begin
          dirty_0_7 <= _GEN_4432;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_8 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_8 <= _GEN_547;
        end else begin
          dirty_0_8 <= _GEN_4433;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_9 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_9 <= _GEN_548;
        end else begin
          dirty_0_9 <= _GEN_4434;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_10 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_10 <= _GEN_549;
        end else begin
          dirty_0_10 <= _GEN_4435;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_11 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_11 <= _GEN_550;
        end else begin
          dirty_0_11 <= _GEN_4436;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_12 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_12 <= _GEN_551;
        end else begin
          dirty_0_12 <= _GEN_4437;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_13 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_13 <= _GEN_552;
        end else begin
          dirty_0_13 <= _GEN_4438;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_14 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_14 <= _GEN_553;
        end else begin
          dirty_0_14 <= _GEN_4439;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 34:26]
      dirty_0_15 <= 1'h0; // @[d_cache.scala 34:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_0_15 <= _GEN_554;
        end else begin
          dirty_0_15 <= _GEN_4440;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_0 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_0 <= _GEN_571;
        end else begin
          dirty_1_0 <= _GEN_4441;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_1 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_1 <= _GEN_572;
        end else begin
          dirty_1_1 <= _GEN_4442;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_2 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_2 <= _GEN_573;
        end else begin
          dirty_1_2 <= _GEN_4443;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_3 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_3 <= _GEN_574;
        end else begin
          dirty_1_3 <= _GEN_4444;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_4 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_4 <= _GEN_575;
        end else begin
          dirty_1_4 <= _GEN_4445;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_5 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_5 <= _GEN_576;
        end else begin
          dirty_1_5 <= _GEN_4446;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_6 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_6 <= _GEN_577;
        end else begin
          dirty_1_6 <= _GEN_4447;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_7 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_7 <= _GEN_578;
        end else begin
          dirty_1_7 <= _GEN_4448;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_8 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_8 <= _GEN_579;
        end else begin
          dirty_1_8 <= _GEN_4449;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_9 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_9 <= _GEN_580;
        end else begin
          dirty_1_9 <= _GEN_4450;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_10 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_10 <= _GEN_581;
        end else begin
          dirty_1_10 <= _GEN_4451;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_11 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_11 <= _GEN_582;
        end else begin
          dirty_1_11 <= _GEN_4452;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_12 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_12 <= _GEN_583;
        end else begin
          dirty_1_12 <= _GEN_4453;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_13 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_13 <= _GEN_584;
        end else begin
          dirty_1_13 <= _GEN_4454;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_14 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_14 <= _GEN_585;
        end else begin
          dirty_1_14 <= _GEN_4455;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 35:26]
      dirty_1_15 <= 1'h0; // @[d_cache.scala 35:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_1_15 <= _GEN_586;
        end else begin
          dirty_1_15 <= _GEN_4456;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_0 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_0 <= _GEN_603;
        end else begin
          dirty_2_0 <= _GEN_4457;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_1 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_1 <= _GEN_604;
        end else begin
          dirty_2_1 <= _GEN_4458;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_2 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_2 <= _GEN_605;
        end else begin
          dirty_2_2 <= _GEN_4459;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_3 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_3 <= _GEN_606;
        end else begin
          dirty_2_3 <= _GEN_4460;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_4 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_4 <= _GEN_607;
        end else begin
          dirty_2_4 <= _GEN_4461;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_5 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_5 <= _GEN_608;
        end else begin
          dirty_2_5 <= _GEN_4462;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_6 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_6 <= _GEN_609;
        end else begin
          dirty_2_6 <= _GEN_4463;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_7 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_7 <= _GEN_610;
        end else begin
          dirty_2_7 <= _GEN_4464;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_8 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_8 <= _GEN_611;
        end else begin
          dirty_2_8 <= _GEN_4465;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_9 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_9 <= _GEN_612;
        end else begin
          dirty_2_9 <= _GEN_4466;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_10 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_10 <= _GEN_613;
        end else begin
          dirty_2_10 <= _GEN_4467;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_11 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_11 <= _GEN_614;
        end else begin
          dirty_2_11 <= _GEN_4468;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_12 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_12 <= _GEN_615;
        end else begin
          dirty_2_12 <= _GEN_4469;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_13 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_13 <= _GEN_616;
        end else begin
          dirty_2_13 <= _GEN_4470;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_14 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_14 <= _GEN_617;
        end else begin
          dirty_2_14 <= _GEN_4471;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 36:26]
      dirty_2_15 <= 1'h0; // @[d_cache.scala 36:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_2_15 <= _GEN_618;
        end else begin
          dirty_2_15 <= _GEN_4472;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_0 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_0 <= _GEN_635;
        end else begin
          dirty_3_0 <= _GEN_4473;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_1 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_1 <= _GEN_636;
        end else begin
          dirty_3_1 <= _GEN_4474;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_2 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_2 <= _GEN_637;
        end else begin
          dirty_3_2 <= _GEN_4475;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_3 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_3 <= _GEN_638;
        end else begin
          dirty_3_3 <= _GEN_4476;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_4 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_4 <= _GEN_639;
        end else begin
          dirty_3_4 <= _GEN_4477;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_5 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_5 <= _GEN_640;
        end else begin
          dirty_3_5 <= _GEN_4478;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_6 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_6 <= _GEN_641;
        end else begin
          dirty_3_6 <= _GEN_4479;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_7 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_7 <= _GEN_642;
        end else begin
          dirty_3_7 <= _GEN_4480;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_8 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_8 <= _GEN_643;
        end else begin
          dirty_3_8 <= _GEN_4481;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_9 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_9 <= _GEN_644;
        end else begin
          dirty_3_9 <= _GEN_4482;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_10 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_10 <= _GEN_645;
        end else begin
          dirty_3_10 <= _GEN_4483;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_11 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_11 <= _GEN_646;
        end else begin
          dirty_3_11 <= _GEN_4484;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_12 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_12 <= _GEN_647;
        end else begin
          dirty_3_12 <= _GEN_4485;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_13 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_13 <= _GEN_648;
        end else begin
          dirty_3_13 <= _GEN_4486;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_14 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_14 <= _GEN_649;
        end else begin
          dirty_3_14 <= _GEN_4487;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 37:26]
      dirty_3_15 <= 1'h0; // @[d_cache.scala 37:26]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (4'h2 == state) begin // @[d_cache.scala 105:18]
          dirty_3_15 <= _GEN_650;
        end else begin
          dirty_3_15 <= _GEN_4488;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 44:34]
      write_back_data <= 512'h0; // @[d_cache.scala 44:34]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          write_back_data <= _GEN_4423;
        end
      end
    end
    write_back_addr <= _GEN_5703[31:0]; // @[d_cache.scala 45:{34,34}]
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_0 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          receive_data_0 <= _GEN_4205;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_1 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          receive_data_1 <= _GEN_4206;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_2 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          receive_data_2 <= _GEN_4207;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_3 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          receive_data_3 <= _GEN_4208;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_4 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          receive_data_4 <= _GEN_4209;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_5 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          receive_data_5 <= _GEN_4210;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_6 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          receive_data_6 <= _GEN_4211;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 50:31]
      receive_data_7 <= 64'h0; // @[d_cache.scala 50:31]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          receive_data_7 <= _GEN_4212;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 51:30]
      receive_num <= 3'h0; // @[d_cache.scala 51:30]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (4'h1 == state) begin // @[d_cache.scala 105:18]
        if (!(way0_hit | way1_hit | way2_hit | way3_hit)) begin // @[d_cache.scala 123:57]
          receive_num <= 3'h0; // @[d_cache.scala 129:29]
        end
      end else if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
        receive_num <= _GEN_4213;
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_0 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_0 <= _GEN_4263;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_1 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_1 <= _GEN_4264;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_2 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_2 <= _GEN_4265;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_3 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_3 <= _GEN_4266;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_4 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_4 <= _GEN_4267;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_5 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_5 <= _GEN_4268;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_6 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_6 <= _GEN_4269;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_7 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_7 <= _GEN_4270;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_8 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_8 <= _GEN_4271;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_9 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_9 <= _GEN_4272;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_10 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_10 <= _GEN_4273;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_11 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_11 <= _GEN_4274;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_12 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_12 <= _GEN_4275;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_13 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_13 <= _GEN_4276;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_14 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_14 <= _GEN_4277;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 52:24]
      quene_15 <= 8'h0; // @[d_cache.scala 52:24]
    end else if (!(4'h0 == state)) begin // @[d_cache.scala 105:18]
      if (!(4'h1 == state)) begin // @[d_cache.scala 105:18]
        if (!(4'h2 == state)) begin // @[d_cache.scala 105:18]
          quene_15 <= _GEN_4278;
        end
      end
    end
    if (reset) begin // @[d_cache.scala 100:24]
      state <= 4'h0; // @[d_cache.scala 100:24]
    end else if (4'h0 == state) begin // @[d_cache.scala 105:18]
      if (io_from_lsu_arvalid) begin // @[d_cache.scala 107:38]
        if (io_from_lsu_araddr >= 32'ha0000000) begin // @[d_cache.scala 108:58]
          state <= 4'h7; // @[d_cache.scala 109:27]
        end else begin
          state <= 4'h1; // @[d_cache.scala 111:27]
        end
      end else if (io_from_lsu_awvalid) begin // @[d_cache.scala 113:44]
        state <= _GEN_129;
      end
    end else if (4'h1 == state) begin // @[d_cache.scala 105:18]
      if (way0_hit | way1_hit | way2_hit | way3_hit) begin // @[d_cache.scala 123:57]
        state <= 4'h0;
      end else begin
        state <= 4'h3; // @[d_cache.scala 128:23]
      end
    end else if (4'h2 == state) begin // @[d_cache.scala 105:18]
      state <= _GEN_522;
    end else begin
      state <= _GEN_4214;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  ram_0_0 = _RAND_0[511:0];
  _RAND_1 = {16{`RANDOM}};
  ram_0_1 = _RAND_1[511:0];
  _RAND_2 = {16{`RANDOM}};
  ram_0_2 = _RAND_2[511:0];
  _RAND_3 = {16{`RANDOM}};
  ram_0_3 = _RAND_3[511:0];
  _RAND_4 = {16{`RANDOM}};
  ram_0_4 = _RAND_4[511:0];
  _RAND_5 = {16{`RANDOM}};
  ram_0_5 = _RAND_5[511:0];
  _RAND_6 = {16{`RANDOM}};
  ram_0_6 = _RAND_6[511:0];
  _RAND_7 = {16{`RANDOM}};
  ram_0_7 = _RAND_7[511:0];
  _RAND_8 = {16{`RANDOM}};
  ram_0_8 = _RAND_8[511:0];
  _RAND_9 = {16{`RANDOM}};
  ram_0_9 = _RAND_9[511:0];
  _RAND_10 = {16{`RANDOM}};
  ram_0_10 = _RAND_10[511:0];
  _RAND_11 = {16{`RANDOM}};
  ram_0_11 = _RAND_11[511:0];
  _RAND_12 = {16{`RANDOM}};
  ram_0_12 = _RAND_12[511:0];
  _RAND_13 = {16{`RANDOM}};
  ram_0_13 = _RAND_13[511:0];
  _RAND_14 = {16{`RANDOM}};
  ram_0_14 = _RAND_14[511:0];
  _RAND_15 = {16{`RANDOM}};
  ram_0_15 = _RAND_15[511:0];
  _RAND_16 = {16{`RANDOM}};
  ram_1_0 = _RAND_16[511:0];
  _RAND_17 = {16{`RANDOM}};
  ram_1_1 = _RAND_17[511:0];
  _RAND_18 = {16{`RANDOM}};
  ram_1_2 = _RAND_18[511:0];
  _RAND_19 = {16{`RANDOM}};
  ram_1_3 = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  ram_1_4 = _RAND_20[511:0];
  _RAND_21 = {16{`RANDOM}};
  ram_1_5 = _RAND_21[511:0];
  _RAND_22 = {16{`RANDOM}};
  ram_1_6 = _RAND_22[511:0];
  _RAND_23 = {16{`RANDOM}};
  ram_1_7 = _RAND_23[511:0];
  _RAND_24 = {16{`RANDOM}};
  ram_1_8 = _RAND_24[511:0];
  _RAND_25 = {16{`RANDOM}};
  ram_1_9 = _RAND_25[511:0];
  _RAND_26 = {16{`RANDOM}};
  ram_1_10 = _RAND_26[511:0];
  _RAND_27 = {16{`RANDOM}};
  ram_1_11 = _RAND_27[511:0];
  _RAND_28 = {16{`RANDOM}};
  ram_1_12 = _RAND_28[511:0];
  _RAND_29 = {16{`RANDOM}};
  ram_1_13 = _RAND_29[511:0];
  _RAND_30 = {16{`RANDOM}};
  ram_1_14 = _RAND_30[511:0];
  _RAND_31 = {16{`RANDOM}};
  ram_1_15 = _RAND_31[511:0];
  _RAND_32 = {16{`RANDOM}};
  ram_2_0 = _RAND_32[511:0];
  _RAND_33 = {16{`RANDOM}};
  ram_2_1 = _RAND_33[511:0];
  _RAND_34 = {16{`RANDOM}};
  ram_2_2 = _RAND_34[511:0];
  _RAND_35 = {16{`RANDOM}};
  ram_2_3 = _RAND_35[511:0];
  _RAND_36 = {16{`RANDOM}};
  ram_2_4 = _RAND_36[511:0];
  _RAND_37 = {16{`RANDOM}};
  ram_2_5 = _RAND_37[511:0];
  _RAND_38 = {16{`RANDOM}};
  ram_2_6 = _RAND_38[511:0];
  _RAND_39 = {16{`RANDOM}};
  ram_2_7 = _RAND_39[511:0];
  _RAND_40 = {16{`RANDOM}};
  ram_2_8 = _RAND_40[511:0];
  _RAND_41 = {16{`RANDOM}};
  ram_2_9 = _RAND_41[511:0];
  _RAND_42 = {16{`RANDOM}};
  ram_2_10 = _RAND_42[511:0];
  _RAND_43 = {16{`RANDOM}};
  ram_2_11 = _RAND_43[511:0];
  _RAND_44 = {16{`RANDOM}};
  ram_2_12 = _RAND_44[511:0];
  _RAND_45 = {16{`RANDOM}};
  ram_2_13 = _RAND_45[511:0];
  _RAND_46 = {16{`RANDOM}};
  ram_2_14 = _RAND_46[511:0];
  _RAND_47 = {16{`RANDOM}};
  ram_2_15 = _RAND_47[511:0];
  _RAND_48 = {16{`RANDOM}};
  ram_3_0 = _RAND_48[511:0];
  _RAND_49 = {16{`RANDOM}};
  ram_3_1 = _RAND_49[511:0];
  _RAND_50 = {16{`RANDOM}};
  ram_3_2 = _RAND_50[511:0];
  _RAND_51 = {16{`RANDOM}};
  ram_3_3 = _RAND_51[511:0];
  _RAND_52 = {16{`RANDOM}};
  ram_3_4 = _RAND_52[511:0];
  _RAND_53 = {16{`RANDOM}};
  ram_3_5 = _RAND_53[511:0];
  _RAND_54 = {16{`RANDOM}};
  ram_3_6 = _RAND_54[511:0];
  _RAND_55 = {16{`RANDOM}};
  ram_3_7 = _RAND_55[511:0];
  _RAND_56 = {16{`RANDOM}};
  ram_3_8 = _RAND_56[511:0];
  _RAND_57 = {16{`RANDOM}};
  ram_3_9 = _RAND_57[511:0];
  _RAND_58 = {16{`RANDOM}};
  ram_3_10 = _RAND_58[511:0];
  _RAND_59 = {16{`RANDOM}};
  ram_3_11 = _RAND_59[511:0];
  _RAND_60 = {16{`RANDOM}};
  ram_3_12 = _RAND_60[511:0];
  _RAND_61 = {16{`RANDOM}};
  ram_3_13 = _RAND_61[511:0];
  _RAND_62 = {16{`RANDOM}};
  ram_3_14 = _RAND_62[511:0];
  _RAND_63 = {16{`RANDOM}};
  ram_3_15 = _RAND_63[511:0];
  _RAND_64 = {1{`RANDOM}};
  tag_0_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  tag_0_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  tag_0_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  tag_0_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  tag_0_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  tag_0_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  tag_0_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  tag_0_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  tag_0_8 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  tag_0_9 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  tag_0_10 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  tag_0_11 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  tag_0_12 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  tag_0_13 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  tag_0_14 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  tag_0_15 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  tag_1_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  tag_1_1 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  tag_1_2 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  tag_1_3 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  tag_1_4 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  tag_1_5 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  tag_1_6 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  tag_1_7 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  tag_1_8 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  tag_1_9 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  tag_1_10 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  tag_1_11 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  tag_1_12 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  tag_1_13 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  tag_1_14 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  tag_1_15 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  tag_2_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  tag_2_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  tag_2_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  tag_2_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  tag_2_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  tag_2_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  tag_2_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  tag_2_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  tag_2_8 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  tag_2_9 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  tag_2_10 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  tag_2_11 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  tag_2_12 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  tag_2_13 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  tag_2_14 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  tag_2_15 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  tag_3_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  tag_3_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  tag_3_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  tag_3_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  tag_3_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  tag_3_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  tag_3_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  tag_3_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  tag_3_8 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  tag_3_9 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  tag_3_10 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  tag_3_11 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  tag_3_12 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  tag_3_13 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  tag_3_14 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  tag_3_15 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_1_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_1_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_1_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_1_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_1_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_1_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_1_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_1_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_1_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_1_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_1_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_1_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_1_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_1_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_1_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_1_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_2_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_2_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_2_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_2_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_2_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_2_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_2_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_2_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_2_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_2_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_2_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_2_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_2_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_2_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_2_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_2_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_3_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_3_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_3_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_3_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_3_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_3_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_3_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_3_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_3_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_3_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_3_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_3_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_3_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_3_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_3_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_3_15 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  dirty_0_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  dirty_0_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dirty_0_2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  dirty_0_3 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  dirty_0_4 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  dirty_0_5 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  dirty_0_6 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  dirty_0_7 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dirty_0_8 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  dirty_0_9 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  dirty_0_10 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  dirty_0_11 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  dirty_0_12 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  dirty_0_13 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dirty_0_14 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  dirty_0_15 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  dirty_1_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  dirty_1_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  dirty_1_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  dirty_1_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dirty_1_4 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  dirty_1_5 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  dirty_1_6 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  dirty_1_7 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  dirty_1_8 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  dirty_1_9 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  dirty_1_10 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  dirty_1_11 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  dirty_1_12 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  dirty_1_13 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  dirty_1_14 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  dirty_1_15 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  dirty_2_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  dirty_2_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  dirty_2_2 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  dirty_2_3 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  dirty_2_4 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  dirty_2_5 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  dirty_2_6 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  dirty_2_7 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  dirty_2_8 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  dirty_2_9 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  dirty_2_10 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  dirty_2_11 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  dirty_2_12 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  dirty_2_13 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  dirty_2_14 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  dirty_2_15 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  dirty_3_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  dirty_3_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  dirty_3_2 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  dirty_3_3 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  dirty_3_4 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  dirty_3_5 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  dirty_3_6 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  dirty_3_7 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  dirty_3_8 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  dirty_3_9 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  dirty_3_10 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  dirty_3_11 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  dirty_3_12 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  dirty_3_13 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  dirty_3_14 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  dirty_3_15 = _RAND_255[0:0];
  _RAND_256 = {16{`RANDOM}};
  write_back_data = _RAND_256[511:0];
  _RAND_257 = {1{`RANDOM}};
  write_back_addr = _RAND_257[31:0];
  _RAND_258 = {2{`RANDOM}};
  receive_data_0 = _RAND_258[63:0];
  _RAND_259 = {2{`RANDOM}};
  receive_data_1 = _RAND_259[63:0];
  _RAND_260 = {2{`RANDOM}};
  receive_data_2 = _RAND_260[63:0];
  _RAND_261 = {2{`RANDOM}};
  receive_data_3 = _RAND_261[63:0];
  _RAND_262 = {2{`RANDOM}};
  receive_data_4 = _RAND_262[63:0];
  _RAND_263 = {2{`RANDOM}};
  receive_data_5 = _RAND_263[63:0];
  _RAND_264 = {2{`RANDOM}};
  receive_data_6 = _RAND_264[63:0];
  _RAND_265 = {2{`RANDOM}};
  receive_data_7 = _RAND_265[63:0];
  _RAND_266 = {1{`RANDOM}};
  receive_num = _RAND_266[2:0];
  _RAND_267 = {1{`RANDOM}};
  quene_0 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  quene_1 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  quene_2 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  quene_3 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  quene_4 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  quene_5 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  quene_6 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  quene_7 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  quene_8 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  quene_9 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  quene_10 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  quene_11 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  quene_12 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  quene_13 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  quene_14 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  quene_15 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  state = _RAND_283[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
